<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-476.906,-594.272,684.937,-1168.55</PageViewport></page 0>
<page 1>
<PageViewport>-410.29,-113.219,813.71,-718.219</PageViewport></page 1>
<page 2>
<PageViewport>-115.222,-806.511,175.239,-950.08</PageViewport>
<gate>
<ID>6151</ID>
<type>AE_DFF_LOW</type>
<position>99,-1631</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4504 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW</type>
<position>142,-3826</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6152</ID>
<type>AE_DFF_LOW</type>
<position>74,-1571</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4417 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>BA_TRI_STATE</type>
<position>175,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6153</ID>
<type>BA_TRI_STATE</type>
<position>109,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4504 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_TRI_STATE</type>
<position>152,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6154</ID>
<type>BA_TRI_STATE</type>
<position>84,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4417 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>188,-3886</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>132 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6155</ID>
<type>AE_DFF_LOW</type>
<position>122,-1631</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4505 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_DFF_LOW</type>
<position>165,-3826</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6156</ID>
<type>AE_DFF_LOW</type>
<position>99,-1571</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4418 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_TRI_STATE</type>
<position>198,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6157</ID>
<type>BA_TRI_STATE</type>
<position>132,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4505 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>BA_TRI_STATE</type>
<position>175,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6158</ID>
<type>BA_TRI_STATE</type>
<position>109,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4418 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_DFF_LOW</type>
<position>213,-3886</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>133 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6159</ID>
<type>AE_DFF_LOW</type>
<position>145,-1631</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4506 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_DFF_LOW</type>
<position>188,-3826</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6160</ID>
<type>AE_DFF_LOW</type>
<position>122,-1571</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4419 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_TRI_STATE</type>
<position>223,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6161</ID>
<type>BA_TRI_STATE</type>
<position>155,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4506 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>BA_TRI_STATE</type>
<position>198,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6162</ID>
<type>BA_TRI_STATE</type>
<position>132,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4419 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_DFF_LOW</type>
<position>236,-3886</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6163</ID>
<type>AE_DFF_LOW</type>
<position>168,-1631</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4507 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_DFF_LOW</type>
<position>213,-3826</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6164</ID>
<type>AE_DFF_LOW</type>
<position>145,-1571</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4420 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_TRI_STATE</type>
<position>246,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6165</ID>
<type>BA_TRI_STATE</type>
<position>178,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4507 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>BA_TRI_STATE</type>
<position>223,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6166</ID>
<type>BA_TRI_STATE</type>
<position>155,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4420 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>43.5,-3868.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6167</ID>
<type>AE_DFF_LOW</type>
<position>193,-1631</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4508 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_DFF_LOW</type>
<position>236,-3826</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6168</ID>
<type>AE_DFF_LOW</type>
<position>168,-1571</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4421 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>55,-3878</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6169</ID>
<type>BA_TRI_STATE</type>
<position>203,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4508 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>BA_TRI_STATE</type>
<position>246,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6170</ID>
<type>BA_TRI_STATE</type>
<position>178,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4421 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_DFF_LOW</type>
<position>71,-3867.5</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>137 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6171</ID>
<type>AE_DFF_LOW</type>
<position>216,-1631</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4509 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>43.5,-3808.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6172</ID>
<type>AE_DFF_LOW</type>
<position>193,-1571</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4422 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>22</ID>
<type>BA_TRI_STATE</type>
<position>81,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>137 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6173</ID>
<type>BA_TRI_STATE</type>
<position>226,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4509 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>54.5,-3818</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6174</ID>
<type>BA_TRI_STATE</type>
<position>203,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4422 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>94,-3867.5</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>138 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6175</ID>
<type>AA_AND2</type>
<position>23.5,-1766</position>
<input>
<ID>IN_0</ID>4575 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>71,-3807.5</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6176</ID>
<type>AE_DFF_LOW</type>
<position>216,-1571</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4423 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_TRI_STATE</type>
<position>104,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>138 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6177</ID>
<type>AA_AND2</type>
<position>34.5,-1775.5</position>
<input>
<ID>IN_0</ID>4575 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4521 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>BA_TRI_STATE</type>
<position>81,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6178</ID>
<type>BA_TRI_STATE</type>
<position>226,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4423 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_DFF_LOW</type>
<position>119,-3867.5</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>139 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6179</ID>
<type>AE_DFF_LOW</type>
<position>51,-1765</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4512 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>94,-3807.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6180</ID>
<type>AA_AND2</type>
<position>34.5,-1738</position>
<input>
<ID>IN_0</ID>4573 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4541 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>BA_TRI_STATE</type>
<position>129,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>139 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6181</ID>
<type>AA_AND2</type>
<position>23.5,-1553</position>
<input>
<ID>IN_0</ID>4467 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>BA_TRI_STATE</type>
<position>104,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6182</ID>
<type>BA_TRI_STATE</type>
<position>61,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4512 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_DFF_LOW</type>
<position>142,-3867.5</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>140 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6183</ID>
<type>AA_AND2</type>
<position>34.5,-1562.5</position>
<input>
<ID>IN_0</ID>4467 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>119,-3807.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6184</ID>
<type>AE_DFF_LOW</type>
<position>74,-1765</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4513 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>BA_TRI_STATE</type>
<position>152,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>140 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6185</ID>
<type>AE_DFF_LOW</type>
<position>51,-1727.5</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4532 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>BA_TRI_STATE</type>
<position>129,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6186</ID>
<type>AE_DFF_LOW</type>
<position>51,-1552</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4426 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_DFF_LOW</type>
<position>165,-3867.5</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>141 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6187</ID>
<type>BA_TRI_STATE</type>
<position>84,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4513 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_DFF_LOW</type>
<position>142,-3807.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6188</ID>
<type>BA_TRI_STATE</type>
<position>61,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4426 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>38</ID>
<type>BA_TRI_STATE</type>
<position>175,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>141 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6189</ID>
<type>AE_DFF_LOW</type>
<position>99,-1765</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4514 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>39</ID>
<type>BA_TRI_STATE</type>
<position>152,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6190</ID>
<type>BA_TRI_STATE</type>
<position>61,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4532 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_DFF_LOW</type>
<position>188,-3867.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>142 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6191</ID>
<type>AE_DFF_LOW</type>
<position>74,-1552</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4427 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_DFF_LOW</type>
<position>165,-3807.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>55 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6192</ID>
<type>BA_TRI_STATE</type>
<position>109,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4514 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>BA_TRI_STATE</type>
<position>198,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6193</ID>
<type>BA_TRI_STATE</type>
<position>84,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4427 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>43</ID>
<type>BA_TRI_STATE</type>
<position>175,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6194</ID>
<type>AE_DFF_LOW</type>
<position>122,-1765</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4515 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>44</ID>
<type>AE_DFF_LOW</type>
<position>213,-3867.5</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>143 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6195</ID>
<type>AE_DFF_LOW</type>
<position>74,-1727.5</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4533 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>188,-3807.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>56 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6196</ID>
<type>AE_DFF_LOW</type>
<position>99,-1552</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4428 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>BA_TRI_STATE</type>
<position>223,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>143 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6197</ID>
<type>BA_TRI_STATE</type>
<position>132,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4515 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>BA_TRI_STATE</type>
<position>198,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6198</ID>
<type>BA_TRI_STATE</type>
<position>109,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4428 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW</type>
<position>236,-3867.5</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>144 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6199</ID>
<type>AE_DFF_LOW</type>
<position>145,-1765</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4516 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_DFF_LOW</type>
<position>213,-3807.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>57 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6200</ID>
<type>BA_TRI_STATE</type>
<position>84,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4533 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>BA_TRI_STATE</type>
<position>246,-3878</position>
<input>
<ID>ENABLE_0</ID>146 </input>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6201</ID>
<type>AE_DFF_LOW</type>
<position>122,-1552</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4429 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>51</ID>
<type>BA_TRI_STATE</type>
<position>223,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6202</ID>
<type>BA_TRI_STATE</type>
<position>155,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4516 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>43.5,-4002.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6203</ID>
<type>BA_TRI_STATE</type>
<position>132,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4429 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_DFF_LOW</type>
<position>236,-3807.5</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6204</ID>
<type>AE_DFF_LOW</type>
<position>168,-1765</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4517 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>54.5,-4012</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6205</ID>
<type>AE_DFF_LOW</type>
<position>99,-1727.5</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4534 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>BA_TRI_STATE</type>
<position>246,-3818</position>
<input>
<ID>ENABLE_0</ID>60 </input>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6206</ID>
<type>AE_DFF_LOW</type>
<position>145,-1552</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4430 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_DFF_LOW</type>
<position>71,-4001.5</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>147 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6207</ID>
<type>BA_TRI_STATE</type>
<position>178,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4517 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND2</type>
<position>54.5,-3974.5</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6208</ID>
<type>BA_TRI_STATE</type>
<position>155,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4430 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>43.5,-3789.5</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6209</ID>
<type>BA_TRI_STATE</type>
<position>109,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4534 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_TRI_STATE</type>
<position>81,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>147 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6210</ID>
<type>AE_DFF_LOW</type>
<position>168,-1552</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4431 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND2</type>
<position>54.5,-3799</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6211</ID>
<type>BA_TRI_STATE</type>
<position>178,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4431 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_DFF_LOW</type>
<position>94,-4001.5</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>148 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6212</ID>
<type>AE_DFF_LOW</type>
<position>122,-1727.5</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4535 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_DFF_LOW</type>
<position>71,-3964</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>167 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6213</ID>
<type>AE_DFF_LOW</type>
<position>193,-1552</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4432 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_DFF_LOW</type>
<position>71,-3788.5</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>61 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6214</ID>
<type>BA_TRI_STATE</type>
<position>203,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4432 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>BA_TRI_STATE</type>
<position>104,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6215</ID>
<type>AE_DFF_LOW</type>
<position>216,-1552</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4433 </output>
<input>
<ID>clock</ID>4434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_TRI_STATE</type>
<position>81,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6216</ID>
<type>BA_TRI_STATE</type>
<position>226,-1562.5</position>
<input>
<ID>ENABLE_0</ID>4435 </input>
<input>
<ID>IN_0</ID>4433 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_DFF_LOW</type>
<position>119,-4001.5</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>149 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6217</ID>
<type>AA_AND2</type>
<position>23.5,-1534.5</position>
<input>
<ID>IN_0</ID>4466 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4444 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>BA_TRI_STATE</type>
<position>81,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6218</ID>
<type>AA_AND2</type>
<position>34.5,-1544</position>
<input>
<ID>IN_0</ID>4466 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_DFF_LOW</type>
<position>94,-3788.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>62 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6219</ID>
<type>AE_DFF_LOW</type>
<position>51,-1533.5</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4436 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>BA_TRI_STATE</type>
<position>129,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>149 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6220</ID>
<type>BA_TRI_STATE</type>
<position>61,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4436 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>BA_TRI_STATE</type>
<position>104,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6221</ID>
<type>AE_DFF_LOW</type>
<position>74,-1533.5</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4437 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_DFF_LOW</type>
<position>142,-4001.5</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>150 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6222</ID>
<type>BA_TRI_STATE</type>
<position>84,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4437 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_DFF_LOW</type>
<position>94,-3964</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>168 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6223</ID>
<type>AE_DFF_LOW</type>
<position>99,-1533.5</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4438 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_DFF_LOW</type>
<position>119,-3788.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>63 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6224</ID>
<type>BA_TRI_STATE</type>
<position>109,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4438 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_TRI_STATE</type>
<position>152,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6225</ID>
<type>AE_DFF_LOW</type>
<position>122,-1533.5</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4439 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>BA_TRI_STATE</type>
<position>129,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6226</ID>
<type>BA_TRI_STATE</type>
<position>132,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4439 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_DFF_LOW</type>
<position>165,-4001.5</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>151 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6227</ID>
<type>AE_DFF_LOW</type>
<position>145,-1533.5</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4440 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>77</ID>
<type>BA_TRI_STATE</type>
<position>104,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6228</ID>
<type>BA_TRI_STATE</type>
<position>155,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4440 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>142,-3788.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6229</ID>
<type>AE_DFF_LOW</type>
<position>168,-1533.5</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4441 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>79</ID>
<type>BA_TRI_STATE</type>
<position>175,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>151 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6230</ID>
<type>BA_TRI_STATE</type>
<position>178,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4441 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>80</ID>
<type>BA_TRI_STATE</type>
<position>152,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6231</ID>
<type>AE_DFF_LOW</type>
<position>193,-1533.5</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4442 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_DFF_LOW</type>
<position>188,-4001.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>152 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6232</ID>
<type>BA_TRI_STATE</type>
<position>203,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4442 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_DFF_LOW</type>
<position>119,-3964</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>169 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6233</ID>
<type>AE_DFF_LOW</type>
<position>216,-1533.5</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4443 </output>
<input>
<ID>clock</ID>4444 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_DFF_LOW</type>
<position>165,-3788.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6234</ID>
<type>BA_TRI_STATE</type>
<position>226,-1544</position>
<input>
<ID>ENABLE_0</ID>4445 </input>
<input>
<ID>IN_0</ID>4443 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>BA_TRI_STATE</type>
<position>198,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6235</ID>
<type>HA_JUNC_2</type>
<position>42.5,-1447</position>
<input>
<ID>N_in0</ID>4446 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>85</ID>
<type>BA_TRI_STATE</type>
<position>175,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6236</ID>
<type>HA_JUNC_2</type>
<position>65.5,-1446.5</position>
<input>
<ID>N_in0</ID>4447 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>86</ID>
<type>BA_TRI_STATE</type>
<position>129,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6237</ID>
<type>HA_JUNC_2</type>
<position>68.5,-1447</position>
<input>
<ID>N_in0</ID>4448 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>87</ID>
<type>AE_DFF_LOW</type>
<position>188,-3788.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6238</ID>
<type>HA_JUNC_2</type>
<position>88,-1446.5</position>
<input>
<ID>N_in0</ID>4449 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>88</ID>
<type>BA_TRI_STATE</type>
<position>198,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6239</ID>
<type>HA_JUNC_2</type>
<position>91.5,-1446.5</position>
<input>
<ID>N_in0</ID>4450 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>89</ID>
<type>AE_DFF_LOW</type>
<position>142,-3964</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>170 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6240</ID>
<type>HA_JUNC_2</type>
<position>112.5,-1447</position>
<input>
<ID>N_in0</ID>4451 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>90</ID>
<type>AE_DFF_LOW</type>
<position>213,-3788.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6241</ID>
<type>HA_JUNC_2</type>
<position>116.5,-1446.5</position>
<input>
<ID>N_in0</ID>4452 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>91</ID>
<type>BA_TRI_STATE</type>
<position>223,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6242</ID>
<type>HA_JUNC_2</type>
<position>135,-1446.5</position>
<input>
<ID>N_in0</ID>4453 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>92</ID>
<type>AE_DFF_LOW</type>
<position>236,-3788.5</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6243</ID>
<type>HA_JUNC_2</type>
<position>139,-1446.5</position>
<input>
<ID>N_in0</ID>4454 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>93</ID>
<type>BA_TRI_STATE</type>
<position>246,-3799</position>
<input>
<ID>ENABLE_0</ID>70 </input>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6244</ID>
<type>HA_JUNC_2</type>
<position>158,-1446.5</position>
<input>
<ID>N_in0</ID>4455 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND2</type>
<position>43.5,-3771</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6245</ID>
<type>HA_JUNC_2</type>
<position>163,-1446.5</position>
<input>
<ID>N_in0</ID>4456 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND2</type>
<position>54.5,-3780.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6246</ID>
<type>HA_JUNC_2</type>
<position>185.5,-1446.5</position>
<input>
<ID>N_in0</ID>4458 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>96</ID>
<type>AE_DFF_LOW</type>
<position>71,-3770</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>71 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6247</ID>
<type>HA_JUNC_2</type>
<position>181,-1446.5</position>
<input>
<ID>N_in0</ID>4457 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>97</ID>
<type>BA_TRI_STATE</type>
<position>81,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6248</ID>
<type>HA_JUNC_2</type>
<position>206.5,-1447</position>
<input>
<ID>N_in0</ID>4459 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>98</ID>
<type>AE_DFF_LOW</type>
<position>94,-3770</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>72 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6249</ID>
<type>HA_JUNC_2</type>
<position>231,-1448</position>
<input>
<ID>N_in0</ID>4461 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>99</ID>
<type>BA_TRI_STATE</type>
<position>104,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6250</ID>
<type>HA_JUNC_2</type>
<position>42.5,-1614</position>
<input>
<ID>N_in0</ID>4580 </input>
<input>
<ID>N_in1</ID>4446 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>100</ID>
<type>AE_DFF_LOW</type>
<position>119,-3770</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6251</ID>
<type>HA_JUNC_2</type>
<position>65.5,-1613.5</position>
<input>
<ID>N_in0</ID>4581 </input>
<input>
<ID>N_in1</ID>4447 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>101</ID>
<type>BA_TRI_STATE</type>
<position>129,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6252</ID>
<type>HA_JUNC_2</type>
<position>68.5,-1613.5</position>
<input>
<ID>N_in0</ID>4582 </input>
<input>
<ID>N_in1</ID>4448 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>102</ID>
<type>AE_DFF_LOW</type>
<position>142,-3770</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6253</ID>
<type>HA_JUNC_2</type>
<position>88,-1613.5</position>
<input>
<ID>N_in0</ID>4583 </input>
<input>
<ID>N_in1</ID>4449 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>103</ID>
<type>BA_TRI_STATE</type>
<position>152,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>74 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6254</ID>
<type>HA_JUNC_2</type>
<position>91.5,-1613.5</position>
<input>
<ID>N_in0</ID>4584 </input>
<input>
<ID>N_in1</ID>4450 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>104</ID>
<type>AE_DFF_LOW</type>
<position>165,-3770</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>75 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6255</ID>
<type>HA_JUNC_2</type>
<position>112.5,-1613.5</position>
<input>
<ID>N_in0</ID>4585 </input>
<input>
<ID>N_in1</ID>4451 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>105</ID>
<type>BA_TRI_STATE</type>
<position>175,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6256</ID>
<type>HA_JUNC_2</type>
<position>116.5,-1613.5</position>
<input>
<ID>N_in0</ID>4586 </input>
<input>
<ID>N_in1</ID>4452 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>106</ID>
<type>AE_DFF_LOW</type>
<position>188,-3770</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6257</ID>
<type>HA_JUNC_2</type>
<position>135,-1613.5</position>
<input>
<ID>N_in0</ID>4587 </input>
<input>
<ID>N_in1</ID>4453 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>107</ID>
<type>BA_TRI_STATE</type>
<position>198,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6258</ID>
<type>HA_JUNC_2</type>
<position>139,-1613.5</position>
<input>
<ID>N_in0</ID>4588 </input>
<input>
<ID>N_in1</ID>4454 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>108</ID>
<type>AE_DFF_LOW</type>
<position>213,-3770</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>77 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6259</ID>
<type>HA_JUNC_2</type>
<position>158,-1613</position>
<input>
<ID>N_in0</ID>4589 </input>
<input>
<ID>N_in1</ID>4455 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>109</ID>
<type>BA_TRI_STATE</type>
<position>223,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6260</ID>
<type>HA_JUNC_2</type>
<position>163,-1613</position>
<input>
<ID>N_in0</ID>4590 </input>
<input>
<ID>N_in1</ID>4456 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>110</ID>
<type>AE_DFF_LOW</type>
<position>236,-3770</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>78 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6261</ID>
<type>HA_JUNC_2</type>
<position>181,-1612.5</position>
<input>
<ID>N_in0</ID>4591 </input>
<input>
<ID>N_in1</ID>4457 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>111</ID>
<type>BA_TRI_STATE</type>
<position>246,-3780.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6262</ID>
<type>HA_JUNC_2</type>
<position>185.5,-1612.5</position>
<input>
<ID>N_in0</ID>4592 </input>
<input>
<ID>N_in1</ID>4458 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>112</ID>
<type>HA_JUNC_2</type>
<position>62.5,-3683.5</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6263</ID>
<type>HA_JUNC_2</type>
<position>206.5,-1612</position>
<input>
<ID>N_in0</ID>4593 </input>
<input>
<ID>N_in1</ID>4459 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>113</ID>
<type>HA_JUNC_2</type>
<position>85.5,-3683</position>
<input>
<ID>N_in0</ID>82 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6264</ID>
<type>HA_JUNC_2</type>
<position>210,-1612</position>
<input>
<ID>N_in0</ID>4594 </input>
<input>
<ID>N_in1</ID>4460 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>114</ID>
<type>HA_JUNC_2</type>
<position>88.5,-3683.5</position>
<input>
<ID>N_in0</ID>83 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6265</ID>
<type>HA_JUNC_2</type>
<position>210,-1447</position>
<input>
<ID>N_in0</ID>4460 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>115</ID>
<type>HA_JUNC_2</type>
<position>108,-3683</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6266</ID>
<type>HA_JUNC_2</type>
<position>231,-1612</position>
<input>
<ID>N_in0</ID>4595 </input>
<input>
<ID>N_in1</ID>4461 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>116</ID>
<type>HA_JUNC_2</type>
<position>111.5,-3683</position>
<input>
<ID>N_in0</ID>85 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6267</ID>
<type>HA_JUNC_2</type>
<position>29.5,-1447</position>
<input>
<ID>N_in0</ID>4471 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>117</ID>
<type>HA_JUNC_2</type>
<position>132.5,-3683.5</position>
<input>
<ID>N_in0</ID>86 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6268</ID>
<type>HA_JUNC_2</type>
<position>19.5,-1447</position>
<input>
<ID>N_in0</ID>4470 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>118</ID>
<type>HA_JUNC_2</type>
<position>136.5,-3683</position>
<input>
<ID>N_in0</ID>87 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6269</ID>
<type>HA_JUNC_2</type>
<position>29.5,-1614</position>
<input>
<ID>N_in0</ID>4579 </input>
<input>
<ID>N_in1</ID>4471 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>119</ID>
<type>HA_JUNC_2</type>
<position>155,-3683</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6270</ID>
<type>HA_JUNC_2</type>
<position>19.5,-1614</position>
<input>
<ID>N_in0</ID>4578 </input>
<input>
<ID>N_in1</ID>4470 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>120</ID>
<type>HA_JUNC_2</type>
<position>159,-3683</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6271</ID>
<type>AA_LABEL</type>
<position>10.5,-1447.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>HA_JUNC_2</type>
<position>178,-3683</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6272</ID>
<type>BI_DECODER_4x16</type>
<position>-129,-1614.5</position>
<output>
<ID>OUT_0</ID>4575 </output>
<output>
<ID>OUT_1</ID>4574 </output>
<output>
<ID>OUT_10</ID>4467 </output>
<output>
<ID>OUT_11</ID>4466 </output>
<output>
<ID>OUT_12</ID>4465 </output>
<output>
<ID>OUT_13</ID>4464 </output>
<output>
<ID>OUT_14</ID>4463 </output>
<output>
<ID>OUT_15</ID>4462 </output>
<output>
<ID>OUT_2</ID>4573 </output>
<output>
<ID>OUT_3</ID>4572 </output>
<output>
<ID>OUT_4</ID>4571 </output>
<output>
<ID>OUT_5</ID>4570 </output>
<output>
<ID>OUT_6</ID>4569 </output>
<output>
<ID>OUT_7</ID>4568 </output>
<output>
<ID>OUT_8</ID>4469 </output>
<output>
<ID>OUT_9</ID>4468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>122</ID>
<type>HA_JUNC_2</type>
<position>183,-3683</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6273</ID>
<type>AE_DFF_LOW</type>
<position>193,-1765</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4518 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>HA_JUNC_2</type>
<position>205.5,-3683</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6274</ID>
<type>BA_TRI_STATE</type>
<position>203,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4518 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>124</ID>
<type>HA_JUNC_2</type>
<position>201,-3683</position>
<input>
<ID>N_in0</ID>92 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6275</ID>
<type>AE_DFF_LOW</type>
<position>216,-1765</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4519 </output>
<input>
<ID>clock</ID>4520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>125</ID>
<type>HA_JUNC_2</type>
<position>226.5,-3683.5</position>
<input>
<ID>N_in0</ID>94 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6276</ID>
<type>BA_TRI_STATE</type>
<position>226,-1775.5</position>
<input>
<ID>ENABLE_0</ID>4521 </input>
<input>
<ID>IN_0</ID>4519 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>126</ID>
<type>HA_JUNC_2</type>
<position>251,-3684.5</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6277</ID>
<type>AA_AND2</type>
<position>23.5,-1747.5</position>
<input>
<ID>IN_0</ID>4574 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4530 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>HA_JUNC_2</type>
<position>62.5,-3850.5</position>
<input>
<ID>N_in0</ID>215 </input>
<input>
<ID>N_in1</ID>81 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6278</ID>
<type>AA_AND2</type>
<position>34.5,-1757</position>
<input>
<ID>IN_0</ID>4574 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4531 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>HA_JUNC_2</type>
<position>85.5,-3850</position>
<input>
<ID>N_in0</ID>216 </input>
<input>
<ID>N_in1</ID>82 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6279</ID>
<type>AE_DFF_LOW</type>
<position>51,-1746.5</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4522 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>129</ID>
<type>HA_JUNC_2</type>
<position>88.5,-3850</position>
<input>
<ID>N_in0</ID>217 </input>
<input>
<ID>N_in1</ID>83 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6280</ID>
<type>BA_TRI_STATE</type>
<position>61,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4522 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>HA_JUNC_2</type>
<position>108,-3850</position>
<input>
<ID>N_in0</ID>218 </input>
<input>
<ID>N_in1</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6281</ID>
<type>AE_DFF_LOW</type>
<position>74,-1746.5</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4523 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>131</ID>
<type>HA_JUNC_2</type>
<position>111.5,-3850</position>
<input>
<ID>N_in0</ID>219 </input>
<input>
<ID>N_in1</ID>85 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6282</ID>
<type>BA_TRI_STATE</type>
<position>84,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4523 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>HA_JUNC_2</type>
<position>132.5,-3850</position>
<input>
<ID>N_in0</ID>220 </input>
<input>
<ID>N_in1</ID>86 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6283</ID>
<type>AE_DFF_LOW</type>
<position>99,-1746.5</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4524 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>133</ID>
<type>HA_JUNC_2</type>
<position>136.5,-3850</position>
<input>
<ID>N_in0</ID>221 </input>
<input>
<ID>N_in1</ID>87 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6284</ID>
<type>BA_TRI_STATE</type>
<position>109,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4524 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>HA_JUNC_2</type>
<position>155,-3850</position>
<input>
<ID>N_in0</ID>222 </input>
<input>
<ID>N_in1</ID>88 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6285</ID>
<type>AE_DFF_LOW</type>
<position>122,-1746.5</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4525 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>135</ID>
<type>HA_JUNC_2</type>
<position>159,-3850</position>
<input>
<ID>N_in0</ID>223 </input>
<input>
<ID>N_in1</ID>89 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6286</ID>
<type>BA_TRI_STATE</type>
<position>132,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4525 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>HA_JUNC_2</type>
<position>178,-3849.5</position>
<input>
<ID>N_in0</ID>224 </input>
<input>
<ID>N_in1</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6287</ID>
<type>AE_DFF_LOW</type>
<position>145,-1746.5</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4526 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>137</ID>
<type>HA_JUNC_2</type>
<position>183,-3849.5</position>
<input>
<ID>N_in0</ID>225 </input>
<input>
<ID>N_in1</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6288</ID>
<type>BA_TRI_STATE</type>
<position>155,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4526 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>HA_JUNC_2</type>
<position>201,-3849</position>
<input>
<ID>N_in0</ID>226 </input>
<input>
<ID>N_in1</ID>92 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6289</ID>
<type>AE_DFF_LOW</type>
<position>168,-1746.5</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4527 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>139</ID>
<type>HA_JUNC_2</type>
<position>205.5,-3849</position>
<input>
<ID>N_in0</ID>227 </input>
<input>
<ID>N_in1</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6290</ID>
<type>BA_TRI_STATE</type>
<position>178,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4527 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>HA_JUNC_2</type>
<position>226.5,-3848.5</position>
<input>
<ID>N_in0</ID>228 </input>
<input>
<ID>N_in1</ID>94 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6291</ID>
<type>AE_DFF_LOW</type>
<position>193,-1746.5</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4528 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>141</ID>
<type>HA_JUNC_2</type>
<position>230,-3848.5</position>
<input>
<ID>N_in0</ID>229 </input>
<input>
<ID>N_in1</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6292</ID>
<type>BA_TRI_STATE</type>
<position>203,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4528 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>142</ID>
<type>HA_JUNC_2</type>
<position>230,-3683.5</position>
<input>
<ID>N_in0</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6293</ID>
<type>AE_DFF_LOW</type>
<position>216,-1746.5</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4529 </output>
<input>
<ID>clock</ID>4530 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>143</ID>
<type>HA_JUNC_2</type>
<position>251,-3848.5</position>
<input>
<ID>N_in0</ID>230 </input>
<input>
<ID>N_in1</ID>96 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6294</ID>
<type>BA_TRI_STATE</type>
<position>226,-1757</position>
<input>
<ID>ENABLE_0</ID>4531 </input>
<input>
<ID>IN_0</ID>4529 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>144</ID>
<type>HA_JUNC_2</type>
<position>49.5,-3683.5</position>
<input>
<ID>N_in0</ID>106 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6295</ID>
<type>AA_AND2</type>
<position>23.5,-1728.5</position>
<input>
<ID>IN_0</ID>4573 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4540 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>HA_JUNC_2</type>
<position>39.5,-3683.5</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6296</ID>
<type>BA_TRI_STATE</type>
<position>132,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4535 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>146</ID>
<type>HA_JUNC_2</type>
<position>49.5,-3850.5</position>
<input>
<ID>N_in0</ID>214 </input>
<input>
<ID>N_in1</ID>106 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6297</ID>
<type>AE_DFF_LOW</type>
<position>145,-1727.5</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4536 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>147</ID>
<type>HA_JUNC_2</type>
<position>39.5,-3850.5</position>
<input>
<ID>N_in0</ID>213 </input>
<input>
<ID>N_in1</ID>105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6298</ID>
<type>BA_TRI_STATE</type>
<position>155,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4536 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_LABEL</type>
<position>30.5,-3684</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6299</ID>
<type>AE_DFF_LOW</type>
<position>168,-1727.5</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4537 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>149</ID>
<type>BI_DECODER_4x16</type>
<position>-109,-3851</position>
<output>
<ID>OUT_0</ID>210 </output>
<output>
<ID>OUT_1</ID>209 </output>
<output>
<ID>OUT_10</ID>102 </output>
<output>
<ID>OUT_11</ID>101 </output>
<output>
<ID>OUT_12</ID>100 </output>
<output>
<ID>OUT_13</ID>99 </output>
<output>
<ID>OUT_14</ID>98 </output>
<output>
<ID>OUT_15</ID>97 </output>
<output>
<ID>OUT_2</ID>208 </output>
<output>
<ID>OUT_3</ID>207 </output>
<output>
<ID>OUT_4</ID>206 </output>
<output>
<ID>OUT_5</ID>205 </output>
<output>
<ID>OUT_6</ID>204 </output>
<output>
<ID>OUT_7</ID>203 </output>
<output>
<ID>OUT_8</ID>104 </output>
<output>
<ID>OUT_9</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6300</ID>
<type>BA_TRI_STATE</type>
<position>178,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4537 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_DFF_LOW</type>
<position>213,-4001.5</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>153 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6301</ID>
<type>AE_DFF_LOW</type>
<position>193,-1727.5</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4538 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>151</ID>
<type>BA_TRI_STATE</type>
<position>223,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6302</ID>
<type>BA_TRI_STATE</type>
<position>203,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4538 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_DFF_LOW</type>
<position>236,-4001.5</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>154 </output>
<input>
<ID>clock</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6303</ID>
<type>AA_AND2</type>
<position>23.5,-1512.5</position>
<input>
<ID>IN_0</ID>4465 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>BA_TRI_STATE</type>
<position>246,-4012</position>
<input>
<ID>ENABLE_0</ID>156 </input>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6304</ID>
<type>AE_DFF_LOW</type>
<position>216,-1727.5</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4539 </output>
<input>
<ID>clock</ID>4540 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND2</type>
<position>43.5,-3984</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6305</ID>
<type>BA_TRI_STATE</type>
<position>226,-1738</position>
<input>
<ID>ENABLE_0</ID>4541 </input>
<input>
<ID>IN_0</ID>4539 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>54.5,-3993.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6306</ID>
<type>AA_AND2</type>
<position>23.5,-1710</position>
<input>
<ID>IN_0</ID>4572 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4550 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>AE_DFF_LOW</type>
<position>71,-3983</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>157 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6307</ID>
<type>AA_AND2</type>
<position>34.5,-1719.5</position>
<input>
<ID>IN_0</ID>4572 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4551 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>BA_TRI_STATE</type>
<position>81,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6308</ID>
<type>AA_AND2</type>
<position>35,-1522</position>
<input>
<ID>IN_0</ID>4465 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4375 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>AE_DFF_LOW</type>
<position>94,-3983</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>158 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6309</ID>
<type>AE_DFF_LOW</type>
<position>51,-1709</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4542 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>159</ID>
<type>BA_TRI_STATE</type>
<position>104,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6310</ID>
<type>BA_TRI_STATE</type>
<position>61,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4542 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_DFF_LOW</type>
<position>119,-3983</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>159 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6311</ID>
<type>AE_DFF_LOW</type>
<position>74,-1709</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4543 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>BA_TRI_STATE</type>
<position>129,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6312</ID>
<type>BA_TRI_STATE</type>
<position>84,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4543 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_DFF_LOW</type>
<position>142,-3983</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>160 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6313</ID>
<type>AE_DFF_LOW</type>
<position>51,-1511.5</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4366 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>163</ID>
<type>BA_TRI_STATE</type>
<position>152,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6314</ID>
<type>AE_DFF_LOW</type>
<position>99,-1709</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4544 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_DFF_LOW</type>
<position>165,-3983</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>161 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6315</ID>
<type>BA_TRI_STATE</type>
<position>109,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4544 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>BA_TRI_STATE</type>
<position>175,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6316</ID>
<type>AE_DFF_LOW</type>
<position>122,-1709</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4545 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_DFF_LOW</type>
<position>188,-3983</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>162 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6317</ID>
<type>BA_TRI_STATE</type>
<position>132,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4545 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>BA_TRI_STATE</type>
<position>198,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>162 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6318</ID>
<type>AE_DFF_LOW</type>
<position>145,-1709</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4546 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_DFF_LOW</type>
<position>213,-3983</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>163 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6319</ID>
<type>BA_TRI_STATE</type>
<position>61,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4366 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>BA_TRI_STATE</type>
<position>223,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6320</ID>
<type>BA_TRI_STATE</type>
<position>155,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4546 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>170</ID>
<type>AE_DFF_LOW</type>
<position>236,-3983</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>164 </output>
<input>
<ID>clock</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6321</ID>
<type>AE_DFF_LOW</type>
<position>168,-1709</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4547 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>BA_TRI_STATE</type>
<position>246,-3993.5</position>
<input>
<ID>ENABLE_0</ID>166 </input>
<input>
<ID>IN_0</ID>164 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6322</ID>
<type>BA_TRI_STATE</type>
<position>178,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4547 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND2</type>
<position>43.5,-3965</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6323</ID>
<type>AE_DFF_LOW</type>
<position>193,-1709</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4548 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>173</ID>
<type>BA_TRI_STATE</type>
<position>152,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6324</ID>
<type>BA_TRI_STATE</type>
<position>203,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4548 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>174</ID>
<type>AE_DFF_LOW</type>
<position>165,-3964</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>171 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6325</ID>
<type>AE_DFF_LOW</type>
<position>216,-1709</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4549 </output>
<input>
<ID>clock</ID>4550 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>175</ID>
<type>BA_TRI_STATE</type>
<position>175,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>171 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6326</ID>
<type>BA_TRI_STATE</type>
<position>226,-1719.5</position>
<input>
<ID>ENABLE_0</ID>4551 </input>
<input>
<ID>IN_0</ID>4549 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_DFF_LOW</type>
<position>188,-3964</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>172 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6327</ID>
<type>HA_JUNC_2</type>
<position>42.5,-1622.5</position>
<input>
<ID>N_in0</ID>4552 </input>
<input>
<ID>N_in1</ID>4580 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>177</ID>
<type>BA_TRI_STATE</type>
<position>198,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6328</ID>
<type>HA_JUNC_2</type>
<position>65.5,-1622</position>
<input>
<ID>N_in0</ID>4553 </input>
<input>
<ID>N_in1</ID>4581 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>178</ID>
<type>AE_DFF_LOW</type>
<position>213,-3964</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>173 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6329</ID>
<type>HA_JUNC_2</type>
<position>68.5,-1622.5</position>
<input>
<ID>N_in0</ID>4554 </input>
<input>
<ID>N_in1</ID>4582 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>179</ID>
<type>BA_TRI_STATE</type>
<position>223,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>173 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6330</ID>
<type>HA_JUNC_2</type>
<position>88,-1622</position>
<input>
<ID>N_in0</ID>4555 </input>
<input>
<ID>N_in1</ID>4583 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_AND2</type>
<position>43.5,-3749</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6331</ID>
<type>HA_JUNC_2</type>
<position>91.5,-1622</position>
<input>
<ID>N_in0</ID>4556 </input>
<input>
<ID>N_in1</ID>4584 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>181</ID>
<type>AE_DFF_LOW</type>
<position>236,-3964</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>174 </output>
<input>
<ID>clock</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6332</ID>
<type>HA_JUNC_2</type>
<position>112.5,-1622.5</position>
<input>
<ID>N_in0</ID>4557 </input>
<input>
<ID>N_in1</ID>4585 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>182</ID>
<type>BA_TRI_STATE</type>
<position>246,-3974.5</position>
<input>
<ID>ENABLE_0</ID>176 </input>
<input>
<ID>IN_0</ID>174 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6333</ID>
<type>HA_JUNC_2</type>
<position>116.5,-1622</position>
<input>
<ID>N_in0</ID>4558 </input>
<input>
<ID>N_in1</ID>4586 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND2</type>
<position>43.5,-3946.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6334</ID>
<type>HA_JUNC_2</type>
<position>135,-1622</position>
<input>
<ID>N_in0</ID>4559 </input>
<input>
<ID>N_in1</ID>4587 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_AND2</type>
<position>54.5,-3956</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6335</ID>
<type>AE_DFF_LOW</type>
<position>74,-1511.5</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4367 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>55,-3758.5</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6336</ID>
<type>HA_JUNC_2</type>
<position>139,-1622</position>
<input>
<ID>N_in0</ID>4560 </input>
<input>
<ID>N_in1</ID>4588 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>186</ID>
<type>AE_DFF_LOW</type>
<position>71,-3945.5</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>177 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6337</ID>
<type>BA_TRI_STATE</type>
<position>84,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4367 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>BA_TRI_STATE</type>
<position>81,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6338</ID>
<type>HA_JUNC_2</type>
<position>158,-1622</position>
<input>
<ID>N_in0</ID>4561 </input>
<input>
<ID>N_in1</ID>4589 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>188</ID>
<type>AE_DFF_LOW</type>
<position>94,-3945.5</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>178 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6339</ID>
<type>AE_DFF_LOW</type>
<position>99,-1511.5</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4368 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>189</ID>
<type>BA_TRI_STATE</type>
<position>104,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>178 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6340</ID>
<type>HA_JUNC_2</type>
<position>163,-1622</position>
<input>
<ID>N_in0</ID>4562 </input>
<input>
<ID>N_in1</ID>4590 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>190</ID>
<type>AE_DFF_LOW</type>
<position>71,-3748</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>1 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6341</ID>
<type>BA_TRI_STATE</type>
<position>109,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4368 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_DFF_LOW</type>
<position>119,-3945.5</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>179 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6342</ID>
<type>HA_JUNC_2</type>
<position>185.5,-1622</position>
<input>
<ID>N_in0</ID>4564 </input>
<input>
<ID>N_in1</ID>4592 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>192</ID>
<type>BA_TRI_STATE</type>
<position>129,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6343</ID>
<type>AE_DFF_LOW</type>
<position>122,-1511.5</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4369 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>193</ID>
<type>AE_DFF_LOW</type>
<position>142,-3945.5</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>180 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6344</ID>
<type>HA_JUNC_2</type>
<position>181,-1622</position>
<input>
<ID>N_in0</ID>4563 </input>
<input>
<ID>N_in1</ID>4591 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>194</ID>
<type>BA_TRI_STATE</type>
<position>152,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6345</ID>
<type>BA_TRI_STATE</type>
<position>132,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4369 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_DFF_LOW</type>
<position>165,-3945.5</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>181 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6346</ID>
<type>HA_JUNC_2</type>
<position>206.5,-1622.5</position>
<input>
<ID>N_in0</ID>4565 </input>
<input>
<ID>N_in1</ID>4593 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>196</ID>
<type>BA_TRI_STATE</type>
<position>81,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6347</ID>
<type>AE_DFF_LOW</type>
<position>145,-1511.5</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4370 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_TRI_STATE</type>
<position>175,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>181 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6348</ID>
<type>HA_JUNC_2</type>
<position>231,-1623.5</position>
<input>
<ID>N_in0</ID>4567 </input>
<input>
<ID>N_in1</ID>4595 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>198</ID>
<type>AE_DFF_LOW</type>
<position>188,-3945.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>182 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6349</ID>
<type>BA_TRI_STATE</type>
<position>155,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4370 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>199</ID>
<type>BA_TRI_STATE</type>
<position>198,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6350</ID>
<type>AA_AND2</type>
<position>23.5,-1688</position>
<input>
<ID>IN_0</ID>4571 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4480 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_DFF_LOW</type>
<position>213,-3945.5</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>183 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6351</ID>
<type>AE_DFF_LOW</type>
<position>168,-1511.5</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4371 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>201</ID>
<type>BA_TRI_STATE</type>
<position>223,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>183 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6352</ID>
<type>AA_AND2</type>
<position>35,-1697.5</position>
<input>
<ID>IN_0</ID>4571 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_DFF_LOW</type>
<position>236,-3945.5</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>184 </output>
<input>
<ID>clock</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6353</ID>
<type>BA_TRI_STATE</type>
<position>178,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4371 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>BA_TRI_STATE</type>
<position>246,-3956</position>
<input>
<ID>ENABLE_0</ID>186 </input>
<input>
<ID>IN_0</ID>184 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6354</ID>
<type>HA_JUNC_2</type>
<position>42.5,-1789.5</position>
<input>
<ID>N_in1</ID>4552 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>204</ID>
<type>HA_JUNC_2</type>
<position>62.5,-3859</position>
<input>
<ID>N_in0</ID>187 </input>
<input>
<ID>N_in1</ID>215 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6355</ID>
<type>AE_DFF_LOW</type>
<position>193,-1511.5</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4372 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>205</ID>
<type>HA_JUNC_2</type>
<position>85.5,-3858.5</position>
<input>
<ID>N_in0</ID>188 </input>
<input>
<ID>N_in1</ID>216 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6356</ID>
<type>AE_DFF_LOW</type>
<position>51,-1687</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4472 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>206</ID>
<type>HA_JUNC_2</type>
<position>88.5,-3859</position>
<input>
<ID>N_in0</ID>189 </input>
<input>
<ID>N_in1</ID>217 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6357</ID>
<type>BA_TRI_STATE</type>
<position>203,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4372 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>HA_JUNC_2</type>
<position>108,-3858.5</position>
<input>
<ID>N_in0</ID>190 </input>
<input>
<ID>N_in1</ID>218 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6358</ID>
<type>HA_JUNC_2</type>
<position>65.5,-1789</position>
<input>
<ID>N_in1</ID>4553 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>208</ID>
<type>HA_JUNC_2</type>
<position>111.5,-3858.5</position>
<input>
<ID>N_in0</ID>191 </input>
<input>
<ID>N_in1</ID>219 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6359</ID>
<type>AE_DFF_LOW</type>
<position>216,-1511.5</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4373 </output>
<input>
<ID>clock</ID>4374 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>209</ID>
<type>HA_JUNC_2</type>
<position>132.5,-3859</position>
<input>
<ID>N_in0</ID>192 </input>
<input>
<ID>N_in1</ID>220 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6360</ID>
<type>HA_JUNC_2</type>
<position>68.5,-1789</position>
<input>
<ID>N_in1</ID>4554 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>210</ID>
<type>HA_JUNC_2</type>
<position>136.5,-3858.5</position>
<input>
<ID>N_in0</ID>193 </input>
<input>
<ID>N_in1</ID>221 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6361</ID>
<type>BA_TRI_STATE</type>
<position>226,-1522</position>
<input>
<ID>ENABLE_0</ID>4375 </input>
<input>
<ID>IN_0</ID>4373 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>211</ID>
<type>HA_JUNC_2</type>
<position>155,-3858.5</position>
<input>
<ID>N_in0</ID>194 </input>
<input>
<ID>N_in1</ID>222 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6362</ID>
<type>HA_JUNC_2</type>
<position>88,-1789</position>
<input>
<ID>N_in1</ID>4555 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>212</ID>
<type>AE_DFF_LOW</type>
<position>94,-3748</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>2 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6363</ID>
<type>AA_AND2</type>
<position>23.5,-1494</position>
<input>
<ID>IN_0</ID>4464 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4384 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>HA_JUNC_2</type>
<position>159,-3858.5</position>
<input>
<ID>N_in0</ID>195 </input>
<input>
<ID>N_in1</ID>223 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6364</ID>
<type>HA_JUNC_2</type>
<position>91.5,-1789</position>
<input>
<ID>N_in1</ID>4556 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>214</ID>
<type>BA_TRI_STATE</type>
<position>104,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6365</ID>
<type>AA_AND2</type>
<position>35,-1503.5</position>
<input>
<ID>IN_0</ID>4464 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4385 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>HA_JUNC_2</type>
<position>178,-3858.5</position>
<input>
<ID>N_in0</ID>196 </input>
<input>
<ID>N_in1</ID>224 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6366</ID>
<type>HA_JUNC_2</type>
<position>112.5,-1789</position>
<input>
<ID>N_in1</ID>4557 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>216</ID>
<type>AE_DFF_LOW</type>
<position>119,-3748</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6367</ID>
<type>AE_DFF_LOW</type>
<position>51,-1493</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4376 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>217</ID>
<type>HA_JUNC_2</type>
<position>183,-3858.5</position>
<input>
<ID>N_in0</ID>197 </input>
<input>
<ID>N_in1</ID>225 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6368</ID>
<type>BA_TRI_STATE</type>
<position>61,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4472 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>BA_TRI_STATE</type>
<position>129,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6369</ID>
<type>BA_TRI_STATE</type>
<position>61,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4376 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>219</ID>
<type>HA_JUNC_2</type>
<position>205.5,-3858.5</position>
<input>
<ID>N_in0</ID>199 </input>
<input>
<ID>N_in1</ID>227 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6370</ID>
<type>HA_JUNC_2</type>
<position>116.5,-1789</position>
<input>
<ID>N_in1</ID>4558 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>220</ID>
<type>AE_DFF_LOW</type>
<position>142,-3748</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>4 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6371</ID>
<type>AE_DFF_LOW</type>
<position>74,-1493</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4377 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>221</ID>
<type>HA_JUNC_2</type>
<position>201,-3858.5</position>
<input>
<ID>N_in0</ID>198 </input>
<input>
<ID>N_in1</ID>226 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6372</ID>
<type>HA_JUNC_2</type>
<position>135,-1789</position>
<input>
<ID>N_in1</ID>4559 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>222</ID>
<type>BA_TRI_STATE</type>
<position>152,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6373</ID>
<type>BA_TRI_STATE</type>
<position>84,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4377 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>223</ID>
<type>HA_JUNC_2</type>
<position>226.5,-3859</position>
<input>
<ID>N_in0</ID>200 </input>
<input>
<ID>N_in1</ID>228 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6374</ID>
<type>HA_JUNC_2</type>
<position>139,-1789</position>
<input>
<ID>N_in1</ID>4560 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>224</ID>
<type>AE_DFF_LOW</type>
<position>165,-3748</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6375</ID>
<type>AE_DFF_LOW</type>
<position>99,-1493</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4378 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>225</ID>
<type>HA_JUNC_2</type>
<position>251,-3860</position>
<input>
<ID>N_in0</ID>202 </input>
<input>
<ID>N_in1</ID>230 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6376</ID>
<type>HA_JUNC_2</type>
<position>158,-1788.5</position>
<input>
<ID>N_in1</ID>4561 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>226</ID>
<type>BA_TRI_STATE</type>
<position>175,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6377</ID>
<type>BA_TRI_STATE</type>
<position>109,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4378 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>43.5,-3924.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6378</ID>
<type>HA_JUNC_2</type>
<position>163,-1788.5</position>
<input>
<ID>N_in1</ID>4562 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>228</ID>
<type>AE_DFF_LOW</type>
<position>188,-3748</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6379</ID>
<type>AE_DFF_LOW</type>
<position>122,-1493</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4379 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND2</type>
<position>55,-3934</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6380</ID>
<type>HA_JUNC_2</type>
<position>181,-1788</position>
<input>
<ID>N_in1</ID>4563 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>230</ID>
<type>BA_TRI_STATE</type>
<position>198,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6381</ID>
<type>BA_TRI_STATE</type>
<position>132,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4379 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>HA_JUNC_2</type>
<position>62.5,-4026</position>
<input>
<ID>N_in1</ID>187 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6382</ID>
<type>HA_JUNC_2</type>
<position>185.5,-1788</position>
<input>
<ID>N_in1</ID>4564 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>232</ID>
<type>AE_DFF_LOW</type>
<position>213,-3748</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6383</ID>
<type>AE_DFF_LOW</type>
<position>145,-1493</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4380 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>233</ID>
<type>AE_DFF_LOW</type>
<position>71,-3923.5</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>107 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6384</ID>
<type>HA_JUNC_2</type>
<position>206.5,-1787.5</position>
<input>
<ID>N_in1</ID>4565 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>234</ID>
<type>BA_TRI_STATE</type>
<position>223,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6385</ID>
<type>BA_TRI_STATE</type>
<position>155,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4380 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>235</ID>
<type>HA_JUNC_2</type>
<position>85.5,-4025.5</position>
<input>
<ID>N_in1</ID>188 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6386</ID>
<type>HA_JUNC_2</type>
<position>210,-1787.5</position>
<input>
<ID>N_in1</ID>4566 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>236</ID>
<type>AE_DFF_LOW</type>
<position>236,-3748</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>8 </output>
<input>
<ID>clock</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6387</ID>
<type>AE_DFF_LOW</type>
<position>168,-1493</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4381 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>237</ID>
<type>HA_JUNC_2</type>
<position>88.5,-4025.5</position>
<input>
<ID>N_in1</ID>189 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6388</ID>
<type>HA_JUNC_2</type>
<position>210,-1622.5</position>
<input>
<ID>N_in0</ID>4566 </input>
<input>
<ID>N_in1</ID>4594 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>238</ID>
<type>BA_TRI_STATE</type>
<position>246,-3758.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6389</ID>
<type>BA_TRI_STATE</type>
<position>178,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4381 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>239</ID>
<type>HA_JUNC_2</type>
<position>108,-4025.5</position>
<input>
<ID>N_in1</ID>190 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6390</ID>
<type>HA_JUNC_2</type>
<position>231,-1787.5</position>
<input>
<ID>N_in1</ID>4567 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>43.5,-3730.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6391</ID>
<type>AE_DFF_LOW</type>
<position>193,-1493</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4382 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>241</ID>
<type>HA_JUNC_2</type>
<position>111.5,-4025.5</position>
<input>
<ID>N_in1</ID>191 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6392</ID>
<type>AE_DFF_LOW</type>
<position>74,-1687</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4473 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_AND2</type>
<position>55,-3740</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6393</ID>
<type>BA_TRI_STATE</type>
<position>203,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4382 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>243</ID>
<type>HA_JUNC_2</type>
<position>132.5,-4025.5</position>
<input>
<ID>N_in1</ID>192 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6394</ID>
<type>BA_TRI_STATE</type>
<position>84,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4473 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_DFF_LOW</type>
<position>71,-3729.5</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>11 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6395</ID>
<type>AE_DFF_LOW</type>
<position>216,-1493</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4383 </output>
<input>
<ID>clock</ID>4384 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>245</ID>
<type>BA_TRI_STATE</type>
<position>81,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>107 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6396</ID>
<type>HA_JUNC_2</type>
<position>29.5,-1622.5</position>
<input>
<ID>N_in0</ID>4577 </input>
<input>
<ID>N_in1</ID>4579 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>246</ID>
<type>BA_TRI_STATE</type>
<position>81,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6397</ID>
<type>BA_TRI_STATE</type>
<position>226,-1503.5</position>
<input>
<ID>ENABLE_0</ID>4385 </input>
<input>
<ID>IN_0</ID>4383 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>247</ID>
<type>HA_JUNC_2</type>
<position>136.5,-4025.5</position>
<input>
<ID>N_in1</ID>193 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6398</ID>
<type>AE_DFF_LOW</type>
<position>99,-1687</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4474 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>248</ID>
<type>AE_DFF_LOW</type>
<position>94,-3729.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6399</ID>
<type>AA_AND2</type>
<position>23.5,-1475</position>
<input>
<ID>IN_0</ID>4463 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>HA_JUNC_2</type>
<position>155,-4025.5</position>
<input>
<ID>N_in1</ID>194 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6400</ID>
<type>HA_JUNC_2</type>
<position>19.5,-1622.5</position>
<input>
<ID>N_in0</ID>4576 </input>
<input>
<ID>N_in1</ID>4578 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>250</ID>
<type>BA_TRI_STATE</type>
<position>104,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6401</ID>
<type>AA_AND2</type>
<position>35,-1484.5</position>
<input>
<ID>IN_0</ID>4463 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4395 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>HA_JUNC_2</type>
<position>159,-4025.5</position>
<input>
<ID>N_in1</ID>195 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6402</ID>
<type>BA_TRI_STATE</type>
<position>109,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4474 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AE_DFF_LOW</type>
<position>119,-3729.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6403</ID>
<type>AE_DFF_LOW</type>
<position>51,-1474</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4386 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>253</ID>
<type>HA_JUNC_2</type>
<position>178,-4025</position>
<input>
<ID>N_in1</ID>196 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6404</ID>
<type>HA_JUNC_2</type>
<position>29.5,-1789.5</position>
<input>
<ID>N_in1</ID>4577 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>254</ID>
<type>BA_TRI_STATE</type>
<position>129,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6405</ID>
<type>BA_TRI_STATE</type>
<position>61,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4386 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>255</ID>
<type>HA_JUNC_2</type>
<position>183,-4025</position>
<input>
<ID>N_in1</ID>197 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6406</ID>
<type>AE_DFF_LOW</type>
<position>122,-1687</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4475 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>256</ID>
<type>AE_DFF_LOW</type>
<position>142,-3729.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6407</ID>
<type>AE_DFF_LOW</type>
<position>74,-1474</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4387 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>257</ID>
<type>HA_JUNC_2</type>
<position>201,-4024.5</position>
<input>
<ID>N_in1</ID>198 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6408</ID>
<type>HA_JUNC_2</type>
<position>19.5,-1789.5</position>
<input>
<ID>N_in1</ID>4576 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>258</ID>
<type>BA_TRI_STATE</type>
<position>152,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6409</ID>
<type>BA_TRI_STATE</type>
<position>84,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4387 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>259</ID>
<type>HA_JUNC_2</type>
<position>205.5,-4024.5</position>
<input>
<ID>N_in1</ID>199 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6410</ID>
<type>BA_TRI_STATE</type>
<position>132,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4475 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_DFF_LOW</type>
<position>165,-3729.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6411</ID>
<type>AE_DFF_LOW</type>
<position>99,-1474</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4388 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>261</ID>
<type>HA_JUNC_2</type>
<position>226.5,-4024</position>
<input>
<ID>N_in1</ID>200 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6412</ID>
<type>AE_DFF_LOW</type>
<position>145,-1687</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4476 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>262</ID>
<type>BA_TRI_STATE</type>
<position>175,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6413</ID>
<type>BA_TRI_STATE</type>
<position>109,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4388 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>263</ID>
<type>HA_JUNC_2</type>
<position>230,-4024</position>
<input>
<ID>N_in1</ID>201 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6414</ID>
<type>AA_LABEL</type>
<position>10.5,-1623</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AE_DFF_LOW</type>
<position>188,-3729.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6415</ID>
<type>AE_DFF_LOW</type>
<position>122,-1474</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4389 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>265</ID>
<type>HA_JUNC_2</type>
<position>230,-3859</position>
<input>
<ID>N_in0</ID>201 </input>
<input>
<ID>N_in1</ID>229 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6416</ID>
<type>BA_TRI_STATE</type>
<position>155,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4476 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>266</ID>
<type>BA_TRI_STATE</type>
<position>198,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6417</ID>
<type>BA_TRI_STATE</type>
<position>132,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4389 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>267</ID>
<type>HA_JUNC_2</type>
<position>251,-4024</position>
<input>
<ID>N_in1</ID>202 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6418</ID>
<type>AE_DFF_LOW</type>
<position>168,-1687</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4477 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>268</ID>
<type>AE_DFF_LOW</type>
<position>213,-3729.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6419</ID>
<type>AE_DFF_LOW</type>
<position>145,-1474</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4390 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_DFF_LOW</type>
<position>94,-3923.5</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>108 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6420</ID>
<type>BA_TRI_STATE</type>
<position>178,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4477 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>BA_TRI_STATE</type>
<position>223,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6421</ID>
<type>BA_TRI_STATE</type>
<position>155,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4390 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>271</ID>
<type>BA_TRI_STATE</type>
<position>104,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6422</ID>
<type>AE_DFF_LOW</type>
<position>193,-1687</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4478 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>272</ID>
<type>AE_DFF_LOW</type>
<position>236,-3729.5</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>18 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6423</ID>
<type>AE_DFF_LOW</type>
<position>168,-1474</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4391 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>273</ID>
<type>HA_JUNC_2</type>
<position>49.5,-3859</position>
<input>
<ID>N_in0</ID>212 </input>
<input>
<ID>N_in1</ID>214 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6424</ID>
<type>BA_TRI_STATE</type>
<position>203,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4478 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>274</ID>
<type>BA_TRI_STATE</type>
<position>246,-3740</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6425</ID>
<type>BA_TRI_STATE</type>
<position>178,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4391 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>275</ID>
<type>AE_DFF_LOW</type>
<position>119,-3923.5</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>109 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6426</ID>
<type>AE_DFF_LOW</type>
<position>216,-1687</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4479 </output>
<input>
<ID>clock</ID>4480 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>43.5,-3711.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6427</ID>
<type>AE_DFF_LOW</type>
<position>193,-1474</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4392 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>277</ID>
<type>HA_JUNC_2</type>
<position>39.5,-3859</position>
<input>
<ID>N_in0</ID>211 </input>
<input>
<ID>N_in1</ID>213 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6428</ID>
<type>BA_TRI_STATE</type>
<position>226,-1697.5</position>
<input>
<ID>ENABLE_0</ID>4481 </input>
<input>
<ID>IN_0</ID>4479 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>55,-3721</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6429</ID>
<type>BA_TRI_STATE</type>
<position>203,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4392 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>279</ID>
<type>BA_TRI_STATE</type>
<position>129,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>109 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6430</ID>
<type>AA_AND2</type>
<position>23.5,-1669.5</position>
<input>
<ID>IN_0</ID>4570 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4490 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AE_DFF_LOW</type>
<position>71,-3710.5</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>21 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6431</ID>
<type>AE_DFF_LOW</type>
<position>216,-1474</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4393 </output>
<input>
<ID>clock</ID>4394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>281</ID>
<type>HA_JUNC_2</type>
<position>49.5,-4026</position>
<input>
<ID>N_in1</ID>212 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6432</ID>
<type>AA_AND2</type>
<position>35,-1679</position>
<input>
<ID>IN_0</ID>4570 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4491 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>BA_TRI_STATE</type>
<position>81,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6433</ID>
<type>BA_TRI_STATE</type>
<position>226,-1484.5</position>
<input>
<ID>ENABLE_0</ID>4395 </input>
<input>
<ID>IN_0</ID>4393 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>283</ID>
<type>AE_DFF_LOW</type>
<position>142,-3923.5</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>110 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6434</ID>
<type>AE_DFF_LOW</type>
<position>51,-1668.5</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4482 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>284</ID>
<type>AE_DFF_LOW</type>
<position>94,-3710.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6435</ID>
<type>AA_AND2</type>
<position>23.5,-1456.5</position>
<input>
<ID>IN_0</ID>4462 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4404 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>HA_JUNC_2</type>
<position>39.5,-4026</position>
<input>
<ID>N_in1</ID>211 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6436</ID>
<type>BA_TRI_STATE</type>
<position>61,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4482 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>286</ID>
<type>BA_TRI_STATE</type>
<position>104,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6437</ID>
<type>AA_AND2</type>
<position>35,-1466</position>
<input>
<ID>IN_0</ID>4462 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4405 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>BA_TRI_STATE</type>
<position>152,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>110 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6438</ID>
<type>AE_DFF_LOW</type>
<position>74,-1668.5</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4483 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_DFF_LOW</type>
<position>119,-3710.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6439</ID>
<type>AE_DFF_LOW</type>
<position>51,-1455.5</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4396 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_DFF_LOW</type>
<position>165,-3923.5</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>111 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6440</ID>
<type>BA_TRI_STATE</type>
<position>84,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4483 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>290</ID>
<type>BA_TRI_STATE</type>
<position>129,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6441</ID>
<type>BA_TRI_STATE</type>
<position>61,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4396 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>30.5,-3859.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6442</ID>
<type>AE_DFF_LOW</type>
<position>99,-1668.5</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4484 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_DFF_LOW</type>
<position>142,-3710.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6443</ID>
<type>AE_DFF_LOW</type>
<position>74,-1455.5</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4397 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>293</ID>
<type>BA_TRI_STATE</type>
<position>175,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>111 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6444</ID>
<type>BA_TRI_STATE</type>
<position>109,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4484 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>294</ID>
<type>BA_TRI_STATE</type>
<position>152,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6445</ID>
<type>BA_TRI_STATE</type>
<position>84,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4397 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>295</ID>
<type>AE_DFF_LOW</type>
<position>188,-3923.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>112 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6446</ID>
<type>AE_DFF_LOW</type>
<position>122,-1668.5</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4485 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>296</ID>
<type>AE_DFF_LOW</type>
<position>165,-3710.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>25 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6447</ID>
<type>AE_DFF_LOW</type>
<position>99,-1455.5</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4398 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>297</ID>
<type>BA_TRI_STATE</type>
<position>198,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6448</ID>
<type>BA_TRI_STATE</type>
<position>132,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4485 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>298</ID>
<type>BA_TRI_STATE</type>
<position>175,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6449</ID>
<type>BA_TRI_STATE</type>
<position>109,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4398 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>299</ID>
<type>AE_DFF_LOW</type>
<position>213,-3923.5</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>113 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6450</ID>
<type>AE_DFF_LOW</type>
<position>145,-1668.5</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4486 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_DFF_LOW</type>
<position>188,-3710.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6451</ID>
<type>AE_DFF_LOW</type>
<position>122,-1455.5</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4399 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>301</ID>
<type>BA_TRI_STATE</type>
<position>223,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6452</ID>
<type>BA_TRI_STATE</type>
<position>155,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4486 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>302</ID>
<type>BA_TRI_STATE</type>
<position>198,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6453</ID>
<type>BA_TRI_STATE</type>
<position>132,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4399 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_DFF_LOW</type>
<position>236,-3923.5</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>114 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6454</ID>
<type>AE_DFF_LOW</type>
<position>168,-1668.5</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4487 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_DFF_LOW</type>
<position>213,-3710.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>27 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6455</ID>
<type>AE_DFF_LOW</type>
<position>145,-1455.5</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4400 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>305</ID>
<type>BA_TRI_STATE</type>
<position>246,-3934</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6456</ID>
<type>BA_TRI_STATE</type>
<position>178,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4487 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>306</ID>
<type>BA_TRI_STATE</type>
<position>223,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6457</ID>
<type>BA_TRI_STATE</type>
<position>155,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4400 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_AND2</type>
<position>43.5,-3906</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6458</ID>
<type>AE_DFF_LOW</type>
<position>193,-1668.5</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4488 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_DFF_LOW</type>
<position>236,-3710.5</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clock</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6459</ID>
<type>AE_DFF_LOW</type>
<position>168,-1455.5</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4401 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_AND2</type>
<position>55,-3915.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6460</ID>
<type>BA_TRI_STATE</type>
<position>203,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4488 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>310</ID>
<type>BA_TRI_STATE</type>
<position>246,-3721</position>
<input>
<ID>ENABLE_0</ID>30 </input>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6461</ID>
<type>BA_TRI_STATE</type>
<position>178,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4401 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>311</ID>
<type>AE_DFF_LOW</type>
<position>71,-3905</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>117 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6462</ID>
<type>AE_DFF_LOW</type>
<position>216,-1668.5</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4489 </output>
<input>
<ID>clock</ID>4490 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_AND2</type>
<position>43.5,-3693</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6463</ID>
<type>AE_DFF_LOW</type>
<position>193,-1455.5</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4402 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>313</ID>
<type>BA_TRI_STATE</type>
<position>81,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6464</ID>
<type>BA_TRI_STATE</type>
<position>226,-1679</position>
<input>
<ID>ENABLE_0</ID>4491 </input>
<input>
<ID>IN_0</ID>4489 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>55,-3702.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6465</ID>
<type>BA_TRI_STATE</type>
<position>203,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4402 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>315</ID>
<type>AE_DFF_LOW</type>
<position>94,-3905</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>118 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6466</ID>
<type>AA_AND2</type>
<position>23.5,-1650.5</position>
<input>
<ID>IN_0</ID>4569 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4500 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AE_DFF_LOW</type>
<position>71,-3692</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>31 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6467</ID>
<type>AE_DFF_LOW</type>
<position>216,-1455.5</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4403 </output>
<input>
<ID>clock</ID>4404 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>317</ID>
<type>BA_TRI_STATE</type>
<position>104,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>118 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6468</ID>
<type>AA_AND2</type>
<position>35,-1660</position>
<input>
<ID>IN_0</ID>4569 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4501 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>BA_TRI_STATE</type>
<position>81,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6469</ID>
<type>BA_TRI_STATE</type>
<position>226,-1466</position>
<input>
<ID>ENABLE_0</ID>4405 </input>
<input>
<ID>IN_0</ID>4403 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_DFF_LOW</type>
<position>119,-3905</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>119 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6470</ID>
<type>AE_DFF_LOW</type>
<position>51,-1649.5</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4492 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_DFF_LOW</type>
<position>94,-3692</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6471</ID>
<type>AA_AND2</type>
<position>23.5,-1590.5</position>
<input>
<ID>IN_0</ID>4469 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>BA_TRI_STATE</type>
<position>129,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6472</ID>
<type>BA_TRI_STATE</type>
<position>61,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4492 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>322</ID>
<type>BA_TRI_STATE</type>
<position>104,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6473</ID>
<type>AA_AND2</type>
<position>34.5,-1600</position>
<input>
<ID>IN_0</ID>4469 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_DFF_LOW</type>
<position>142,-3905</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>120 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6474</ID>
<type>AE_DFF_LOW</type>
<position>74,-1649.5</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4493 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_DFF_LOW</type>
<position>119,-3692</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>33 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6475</ID>
<type>AE_DFF_LOW</type>
<position>51,-1589.5</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4406 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>325</ID>
<type>BA_TRI_STATE</type>
<position>152,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>120 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6476</ID>
<type>BA_TRI_STATE</type>
<position>84,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4493 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>326</ID>
<type>BA_TRI_STATE</type>
<position>129,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6477</ID>
<type>BA_TRI_STATE</type>
<position>61,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4406 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>327</ID>
<type>AE_DFF_LOW</type>
<position>165,-3905</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>121 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6478</ID>
<type>AE_DFF_LOW</type>
<position>99,-1649.5</position>
<input>
<ID>IN_0</ID>4556 </input>
<output>
<ID>OUT_0</ID>4494 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>328</ID>
<type>AE_DFF_LOW</type>
<position>142,-3692</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6479</ID>
<type>AE_DFF_LOW</type>
<position>74,-1589.5</position>
<input>
<ID>IN_0</ID>4448 </input>
<output>
<ID>OUT_0</ID>4407 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>329</ID>
<type>BA_TRI_STATE</type>
<position>175,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6480</ID>
<type>BA_TRI_STATE</type>
<position>109,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4494 </input>
<output>
<ID>OUT_0</ID>4557 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>330</ID>
<type>BA_TRI_STATE</type>
<position>152,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6481</ID>
<type>BA_TRI_STATE</type>
<position>84,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4407 </input>
<output>
<ID>OUT_0</ID>4449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>331</ID>
<type>AE_DFF_LOW</type>
<position>188,-3905</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>122 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6482</ID>
<type>AE_DFF_LOW</type>
<position>122,-1649.5</position>
<input>
<ID>IN_0</ID>4558 </input>
<output>
<ID>OUT_0</ID>4495 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_DFF_LOW</type>
<position>165,-3692</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6483</ID>
<type>AE_DFF_LOW</type>
<position>99,-1589.5</position>
<input>
<ID>IN_0</ID>4450 </input>
<output>
<ID>OUT_0</ID>4408 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>333</ID>
<type>BA_TRI_STATE</type>
<position>198,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>122 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6484</ID>
<type>BA_TRI_STATE</type>
<position>132,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4495 </input>
<output>
<ID>OUT_0</ID>4559 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>334</ID>
<type>BA_TRI_STATE</type>
<position>175,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6485</ID>
<type>BA_TRI_STATE</type>
<position>109,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4408 </input>
<output>
<ID>OUT_0</ID>4451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_DFF_LOW</type>
<position>213,-3905</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>123 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6486</ID>
<type>AE_DFF_LOW</type>
<position>145,-1649.5</position>
<input>
<ID>IN_0</ID>4560 </input>
<output>
<ID>OUT_0</ID>4496 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_DFF_LOW</type>
<position>188,-3692</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>36 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>337</ID>
<type>BA_TRI_STATE</type>
<position>223,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6488</ID>
<type>AA_LABEL</type>
<position>267,-1617.5</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>BA_TRI_STATE</type>
<position>198,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6489</ID>
<type>AE_DFF_LOW</type>
<position>120,-1962.5</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4639 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>339</ID>
<type>AE_DFF_LOW</type>
<position>236,-3905</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>124 </output>
<input>
<ID>clock</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6490</ID>
<type>BA_TRI_STATE</type>
<position>153,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4726 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>340</ID>
<type>AE_DFF_LOW</type>
<position>213,-3692</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6491</ID>
<type>BA_TRI_STATE</type>
<position>130,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4639 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>341</ID>
<type>BA_TRI_STATE</type>
<position>246,-3915.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6492</ID>
<type>AE_DFF_LOW</type>
<position>166,-2022.5</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4727 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>342</ID>
<type>BA_TRI_STATE</type>
<position>223,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6493</ID>
<type>AE_DFF_LOW</type>
<position>143,-1962.5</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4640 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_AND2</type>
<position>43.5,-3887</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6494</ID>
<type>BA_TRI_STATE</type>
<position>176,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4727 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_DFF_LOW</type>
<position>236,-3692</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6495</ID>
<type>BA_TRI_STATE</type>
<position>153,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4640 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_AND2</type>
<position>55,-3896.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6496</ID>
<type>AE_DFF_LOW</type>
<position>191,-2022.5</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4728 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>346</ID>
<type>BA_TRI_STATE</type>
<position>246,-3702.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6497</ID>
<type>AE_DFF_LOW</type>
<position>166,-1962.5</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4641 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>347</ID>
<type>AE_DFF_LOW</type>
<position>71,-3886</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>127 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6498</ID>
<type>BA_TRI_STATE</type>
<position>201,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4728 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_AND2</type>
<position>43.5,-3827</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6499</ID>
<type>BA_TRI_STATE</type>
<position>176,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4641 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>349</ID>
<type>BA_TRI_STATE</type>
<position>81,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6500</ID>
<type>AE_DFF_LOW</type>
<position>214,-2022.5</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4729 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_AND2</type>
<position>54.5,-3836.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6501</ID>
<type>AE_DFF_LOW</type>
<position>191,-1962.5</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4642 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>351</ID>
<type>AE_DFF_LOW</type>
<position>94,-3886</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>128 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6502</ID>
<type>BA_TRI_STATE</type>
<position>224,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4729 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>352</ID>
<type>AE_DFF_LOW</type>
<position>71,-3826</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6503</ID>
<type>BA_TRI_STATE</type>
<position>201,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4642 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>353</ID>
<type>BA_TRI_STATE</type>
<position>104,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>128 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6504</ID>
<type>AA_AND2</type>
<position>21.5,-2005</position>
<input>
<ID>IN_0</ID>4798 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4740 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>BA_TRI_STATE</type>
<position>81,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6505</ID>
<type>AE_DFF_LOW</type>
<position>214,-1962.5</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4643 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>355</ID>
<type>AE_DFF_LOW</type>
<position>119,-3886</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>129 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6506</ID>
<type>AA_AND2</type>
<position>33,-2014.5</position>
<input>
<ID>IN_0</ID>4798 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4741 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AE_DFF_LOW</type>
<position>94,-3826</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>42 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6507</ID>
<type>BA_TRI_STATE</type>
<position>224,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4643 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>357</ID>
<type>BA_TRI_STATE</type>
<position>129,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6508</ID>
<type>AE_DFF_LOW</type>
<position>49,-2004</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4732 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>358</ID>
<type>BA_TRI_STATE</type>
<position>104,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6509</ID>
<type>AA_AND2</type>
<position>21.5,-1945</position>
<input>
<ID>IN_0</ID>4698 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AE_DFF_LOW</type>
<position>142,-3886</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>130 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6510</ID>
<type>BA_TRI_STATE</type>
<position>59,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4732 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>360</ID>
<type>AE_DFF_LOW</type>
<position>119,-3826</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6511</ID>
<type>AA_AND2</type>
<position>32.5,-1954.5</position>
<input>
<ID>IN_0</ID>4698 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4655 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>BA_TRI_STATE</type>
<position>152,-3896.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6512</ID>
<type>AE_DFF_LOW</type>
<position>72,-2004</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4733 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>362</ID>
<type>BA_TRI_STATE</type>
<position>129,-3836.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6513</ID>
<type>AE_DFF_LOW</type>
<position>49,-1944</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4646 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>363</ID>
<type>AE_DFF_LOW</type>
<position>165,-3886</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>131 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6514</ID>
<type>BA_TRI_STATE</type>
<position>82,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4733 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6515</ID>
<type>BA_TRI_STATE</type>
<position>59,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4646 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6516</ID>
<type>AE_DFF_LOW</type>
<position>97,-2004</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4734 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6517</ID>
<type>AE_DFF_LOW</type>
<position>72,-1944</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4647 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6518</ID>
<type>BA_TRI_STATE</type>
<position>107,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4734 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6519</ID>
<type>BA_TRI_STATE</type>
<position>82,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4647 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6520</ID>
<type>AE_DFF_LOW</type>
<position>120,-2004</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4735 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6521</ID>
<type>AE_DFF_LOW</type>
<position>97,-1944</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4648 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6522</ID>
<type>BA_TRI_STATE</type>
<position>130,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4735 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6523</ID>
<type>BA_TRI_STATE</type>
<position>107,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4648 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6524</ID>
<type>AE_DFF_LOW</type>
<position>143,-2004</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4736 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6525</ID>
<type>AE_DFF_LOW</type>
<position>120,-1944</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4649 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6526</ID>
<type>BA_TRI_STATE</type>
<position>153,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4736 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6527</ID>
<type>BA_TRI_STATE</type>
<position>130,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4649 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6528</ID>
<type>AE_DFF_LOW</type>
<position>166,-2004</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4737 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6529</ID>
<type>AE_DFF_LOW</type>
<position>143,-1944</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4650 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6530</ID>
<type>BA_TRI_STATE</type>
<position>176,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4737 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6531</ID>
<type>BA_TRI_STATE</type>
<position>153,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4650 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6532</ID>
<type>AE_DFF_LOW</type>
<position>191,-2004</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4738 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6533</ID>
<type>AE_DFF_LOW</type>
<position>166,-1944</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4651 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6534</ID>
<type>BA_TRI_STATE</type>
<position>201,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4738 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6535</ID>
<type>BA_TRI_STATE</type>
<position>176,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4651 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6536</ID>
<type>AE_DFF_LOW</type>
<position>214,-2004</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4739 </output>
<input>
<ID>clock</ID>4740 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6537</ID>
<type>AE_DFF_LOW</type>
<position>191,-1944</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4652 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6538</ID>
<type>BA_TRI_STATE</type>
<position>224,-2014.5</position>
<input>
<ID>ENABLE_0</ID>4741 </input>
<input>
<ID>IN_0</ID>4739 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6539</ID>
<type>BA_TRI_STATE</type>
<position>201,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4652 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6540</ID>
<type>AA_AND2</type>
<position>21.5,-2139</position>
<input>
<ID>IN_0</ID>4805 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4750 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6541</ID>
<type>AE_DFF_LOW</type>
<position>214,-1944</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4653 </output>
<input>
<ID>clock</ID>4654 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6542</ID>
<type>AA_AND2</type>
<position>32.5,-2148.5</position>
<input>
<ID>IN_0</ID>4805 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4751 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6543</ID>
<type>BA_TRI_STATE</type>
<position>224,-1954.5</position>
<input>
<ID>ENABLE_0</ID>4655 </input>
<input>
<ID>IN_0</ID>4653 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6544</ID>
<type>AE_DFF_LOW</type>
<position>49,-2138</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4742 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6545</ID>
<type>AA_AND2</type>
<position>32.5,-2111</position>
<input>
<ID>IN_0</ID>4803 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6546</ID>
<type>AA_AND2</type>
<position>21.5,-1926</position>
<input>
<ID>IN_0</ID>4697 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4664 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6547</ID>
<type>BA_TRI_STATE</type>
<position>59,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4742 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6548</ID>
<type>AA_AND2</type>
<position>32.5,-1935.5</position>
<input>
<ID>IN_0</ID>4697 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4665 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6549</ID>
<type>AE_DFF_LOW</type>
<position>72,-2138</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4743 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6550</ID>
<type>AE_DFF_LOW</type>
<position>49,-2100.5</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4762 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6551</ID>
<type>AE_DFF_LOW</type>
<position>49,-1925</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4656 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6552</ID>
<type>BA_TRI_STATE</type>
<position>82,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4743 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6553</ID>
<type>BA_TRI_STATE</type>
<position>59,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4656 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6554</ID>
<type>AE_DFF_LOW</type>
<position>97,-2138</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4744 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6555</ID>
<type>BA_TRI_STATE</type>
<position>59,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4762 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6556</ID>
<type>AE_DFF_LOW</type>
<position>72,-1925</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4657 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6557</ID>
<type>BA_TRI_STATE</type>
<position>107,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4744 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6558</ID>
<type>BA_TRI_STATE</type>
<position>82,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4657 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6559</ID>
<type>AE_DFF_LOW</type>
<position>120,-2138</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4745 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6560</ID>
<type>AE_DFF_LOW</type>
<position>72,-2100.5</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4763 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6561</ID>
<type>AE_DFF_LOW</type>
<position>97,-1925</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4658 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6562</ID>
<type>BA_TRI_STATE</type>
<position>130,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4745 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6563</ID>
<type>BA_TRI_STATE</type>
<position>107,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4658 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6564</ID>
<type>AE_DFF_LOW</type>
<position>143,-2138</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4746 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6565</ID>
<type>BA_TRI_STATE</type>
<position>82,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4763 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6566</ID>
<type>AE_DFF_LOW</type>
<position>120,-1925</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4659 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6567</ID>
<type>BA_TRI_STATE</type>
<position>153,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4746 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6568</ID>
<type>BA_TRI_STATE</type>
<position>130,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4659 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6569</ID>
<type>AE_DFF_LOW</type>
<position>166,-2138</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4747 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6570</ID>
<type>AE_DFF_LOW</type>
<position>97,-2100.5</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4764 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6571</ID>
<type>AE_DFF_LOW</type>
<position>143,-1925</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4660 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6572</ID>
<type>BA_TRI_STATE</type>
<position>176,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4747 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6573</ID>
<type>BA_TRI_STATE</type>
<position>153,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4660 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6574</ID>
<type>BA_TRI_STATE</type>
<position>107,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4764 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6575</ID>
<type>AE_DFF_LOW</type>
<position>166,-1925</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4661 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6576</ID>
<type>BA_TRI_STATE</type>
<position>176,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4661 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6577</ID>
<type>AE_DFF_LOW</type>
<position>120,-2100.5</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4765 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6578</ID>
<type>AE_DFF_LOW</type>
<position>191,-1925</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4662 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6579</ID>
<type>BA_TRI_STATE</type>
<position>201,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4662 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6580</ID>
<type>AE_DFF_LOW</type>
<position>214,-1925</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4663 </output>
<input>
<ID>clock</ID>4664 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6581</ID>
<type>BA_TRI_STATE</type>
<position>224,-1935.5</position>
<input>
<ID>ENABLE_0</ID>4665 </input>
<input>
<ID>IN_0</ID>4663 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6582</ID>
<type>AA_AND2</type>
<position>21.5,-1907.5</position>
<input>
<ID>IN_0</ID>4696 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4674 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6583</ID>
<type>AA_AND2</type>
<position>32.5,-1917</position>
<input>
<ID>IN_0</ID>4696 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4675 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6584</ID>
<type>AE_DFF_LOW</type>
<position>49,-1906.5</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4666 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6585</ID>
<type>BA_TRI_STATE</type>
<position>59,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4666 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6586</ID>
<type>AE_DFF_LOW</type>
<position>72,-1906.5</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4667 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6587</ID>
<type>BA_TRI_STATE</type>
<position>82,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4667 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6588</ID>
<type>AE_DFF_LOW</type>
<position>97,-1906.5</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4668 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6589</ID>
<type>BA_TRI_STATE</type>
<position>107,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4668 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6590</ID>
<type>AE_DFF_LOW</type>
<position>120,-1906.5</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4669 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6591</ID>
<type>BA_TRI_STATE</type>
<position>130,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4669 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6592</ID>
<type>AE_DFF_LOW</type>
<position>143,-1906.5</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4670 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6593</ID>
<type>BA_TRI_STATE</type>
<position>153,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4670 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6594</ID>
<type>AE_DFF_LOW</type>
<position>166,-1906.5</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4671 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6595</ID>
<type>BA_TRI_STATE</type>
<position>176,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4671 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6596</ID>
<type>AE_DFF_LOW</type>
<position>191,-1906.5</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4672 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6597</ID>
<type>BA_TRI_STATE</type>
<position>201,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4672 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6598</ID>
<type>AE_DFF_LOW</type>
<position>214,-1906.5</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4673 </output>
<input>
<ID>clock</ID>4674 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6599</ID>
<type>BA_TRI_STATE</type>
<position>224,-1917</position>
<input>
<ID>ENABLE_0</ID>4675 </input>
<input>
<ID>IN_0</ID>4673 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6600</ID>
<type>HA_JUNC_2</type>
<position>40.5,-1820</position>
<input>
<ID>N_in0</ID>4676 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6601</ID>
<type>HA_JUNC_2</type>
<position>63.5,-1819.5</position>
<input>
<ID>N_in0</ID>4677 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6602</ID>
<type>HA_JUNC_2</type>
<position>66.5,-1820</position>
<input>
<ID>N_in0</ID>4678 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6603</ID>
<type>HA_JUNC_2</type>
<position>86,-1819.5</position>
<input>
<ID>N_in0</ID>4679 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6604</ID>
<type>HA_JUNC_2</type>
<position>89.5,-1819.5</position>
<input>
<ID>N_in0</ID>4680 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6605</ID>
<type>HA_JUNC_2</type>
<position>110.5,-1820</position>
<input>
<ID>N_in0</ID>4681 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6606</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1819.5</position>
<input>
<ID>N_in0</ID>4682 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6607</ID>
<type>HA_JUNC_2</type>
<position>133,-1819.5</position>
<input>
<ID>N_in0</ID>4683 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6608</ID>
<type>HA_JUNC_2</type>
<position>137,-1819.5</position>
<input>
<ID>N_in0</ID>4684 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6609</ID>
<type>HA_JUNC_2</type>
<position>156,-1819.5</position>
<input>
<ID>N_in0</ID>4685 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6610</ID>
<type>HA_JUNC_2</type>
<position>161,-1819.5</position>
<input>
<ID>N_in0</ID>4686 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6611</ID>
<type>HA_JUNC_2</type>
<position>183.5,-1819.5</position>
<input>
<ID>N_in0</ID>4688 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6612</ID>
<type>HA_JUNC_2</type>
<position>179,-1819.5</position>
<input>
<ID>N_in0</ID>4687 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6613</ID>
<type>HA_JUNC_2</type>
<position>204.5,-1820</position>
<input>
<ID>N_in0</ID>4689 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6614</ID>
<type>HA_JUNC_2</type>
<position>229,-1821</position>
<input>
<ID>N_in0</ID>4691 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6615</ID>
<type>HA_JUNC_2</type>
<position>40.5,-1987</position>
<input>
<ID>N_in0</ID>4810 </input>
<input>
<ID>N_in1</ID>4676 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6616</ID>
<type>HA_JUNC_2</type>
<position>63.5,-1986.5</position>
<input>
<ID>N_in0</ID>4811 </input>
<input>
<ID>N_in1</ID>4677 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6617</ID>
<type>HA_JUNC_2</type>
<position>66.5,-1986.5</position>
<input>
<ID>N_in0</ID>4812 </input>
<input>
<ID>N_in1</ID>4678 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6618</ID>
<type>HA_JUNC_2</type>
<position>86,-1986.5</position>
<input>
<ID>N_in0</ID>4813 </input>
<input>
<ID>N_in1</ID>4679 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6619</ID>
<type>HA_JUNC_2</type>
<position>89.5,-1986.5</position>
<input>
<ID>N_in0</ID>4814 </input>
<input>
<ID>N_in1</ID>4680 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6620</ID>
<type>HA_JUNC_2</type>
<position>110.5,-1986.5</position>
<input>
<ID>N_in0</ID>4815 </input>
<input>
<ID>N_in1</ID>4681 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6621</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1986.5</position>
<input>
<ID>N_in0</ID>4816 </input>
<input>
<ID>N_in1</ID>4682 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6622</ID>
<type>HA_JUNC_2</type>
<position>133,-1986.5</position>
<input>
<ID>N_in0</ID>4817 </input>
<input>
<ID>N_in1</ID>4683 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6623</ID>
<type>HA_JUNC_2</type>
<position>137,-1986.5</position>
<input>
<ID>N_in0</ID>4818 </input>
<input>
<ID>N_in1</ID>4684 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6624</ID>
<type>HA_JUNC_2</type>
<position>156,-1986</position>
<input>
<ID>N_in0</ID>4819 </input>
<input>
<ID>N_in1</ID>4685 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6625</ID>
<type>HA_JUNC_2</type>
<position>161,-1986</position>
<input>
<ID>N_in0</ID>4820 </input>
<input>
<ID>N_in1</ID>4686 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6626</ID>
<type>HA_JUNC_2</type>
<position>179,-1985.5</position>
<input>
<ID>N_in0</ID>4821 </input>
<input>
<ID>N_in1</ID>4687 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6627</ID>
<type>HA_JUNC_2</type>
<position>183.5,-1985.5</position>
<input>
<ID>N_in0</ID>4822 </input>
<input>
<ID>N_in1</ID>4688 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6628</ID>
<type>HA_JUNC_2</type>
<position>204.5,-1985</position>
<input>
<ID>N_in0</ID>4823 </input>
<input>
<ID>N_in1</ID>4689 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6629</ID>
<type>HA_JUNC_2</type>
<position>208,-1985</position>
<input>
<ID>N_in0</ID>4824 </input>
<input>
<ID>N_in1</ID>4690 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6630</ID>
<type>HA_JUNC_2</type>
<position>208,-1820</position>
<input>
<ID>N_in0</ID>4690 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6631</ID>
<type>HA_JUNC_2</type>
<position>229,-1985</position>
<input>
<ID>N_in0</ID>4825 </input>
<input>
<ID>N_in1</ID>4691 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6632</ID>
<type>HA_JUNC_2</type>
<position>27.5,-1820</position>
<input>
<ID>N_in0</ID>4701 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6633</ID>
<type>HA_JUNC_2</type>
<position>17.5,-1820</position>
<input>
<ID>N_in0</ID>4700 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6634</ID>
<type>HA_JUNC_2</type>
<position>27.5,-1987</position>
<input>
<ID>N_in0</ID>4809 </input>
<input>
<ID>N_in1</ID>4701 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6635</ID>
<type>HA_JUNC_2</type>
<position>17.5,-1987</position>
<input>
<ID>N_in0</ID>4808 </input>
<input>
<ID>N_in1</ID>4700 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6636</ID>
<type>AA_LABEL</type>
<position>8.5,-1820.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6637</ID>
<type>BI_DECODER_4x16</type>
<position>-131,-1987.5</position>
<output>
<ID>OUT_0</ID>4805 </output>
<output>
<ID>OUT_1</ID>4804 </output>
<output>
<ID>OUT_10</ID>4697 </output>
<output>
<ID>OUT_11</ID>4696 </output>
<output>
<ID>OUT_12</ID>4695 </output>
<output>
<ID>OUT_13</ID>4694 </output>
<output>
<ID>OUT_14</ID>4693 </output>
<output>
<ID>OUT_15</ID>4692 </output>
<output>
<ID>OUT_2</ID>4803 </output>
<output>
<ID>OUT_3</ID>4802 </output>
<output>
<ID>OUT_4</ID>4801 </output>
<output>
<ID>OUT_5</ID>4800 </output>
<output>
<ID>OUT_6</ID>4799 </output>
<output>
<ID>OUT_7</ID>4798 </output>
<output>
<ID>OUT_8</ID>4699 </output>
<output>
<ID>OUT_9</ID>4698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6638</ID>
<type>AE_DFF_LOW</type>
<position>191,-2138</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4748 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6639</ID>
<type>BA_TRI_STATE</type>
<position>201,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4748 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6640</ID>
<type>AE_DFF_LOW</type>
<position>214,-2138</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4749 </output>
<input>
<ID>clock</ID>4750 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6641</ID>
<type>BA_TRI_STATE</type>
<position>224,-2148.5</position>
<input>
<ID>ENABLE_0</ID>4751 </input>
<input>
<ID>IN_0</ID>4749 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6642</ID>
<type>AA_AND2</type>
<position>21.5,-2120.5</position>
<input>
<ID>IN_0</ID>4804 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4760 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6643</ID>
<type>AA_AND2</type>
<position>32.5,-2130</position>
<input>
<ID>IN_0</ID>4804 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4761 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6644</ID>
<type>AE_DFF_LOW</type>
<position>49,-2119.5</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4752 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6645</ID>
<type>BA_TRI_STATE</type>
<position>59,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4752 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6646</ID>
<type>AE_DFF_LOW</type>
<position>72,-2119.5</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4753 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6647</ID>
<type>BA_TRI_STATE</type>
<position>82,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4753 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6648</ID>
<type>AE_DFF_LOW</type>
<position>97,-2119.5</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4754 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6649</ID>
<type>BA_TRI_STATE</type>
<position>107,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4754 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6650</ID>
<type>AE_DFF_LOW</type>
<position>120,-2119.5</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4755 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6651</ID>
<type>BA_TRI_STATE</type>
<position>130,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4755 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6652</ID>
<type>AE_DFF_LOW</type>
<position>143,-2119.5</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4756 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6653</ID>
<type>BA_TRI_STATE</type>
<position>153,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4756 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6654</ID>
<type>AE_DFF_LOW</type>
<position>166,-2119.5</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4757 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6655</ID>
<type>BA_TRI_STATE</type>
<position>176,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4757 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6656</ID>
<type>AE_DFF_LOW</type>
<position>191,-2119.5</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4758 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6657</ID>
<type>BA_TRI_STATE</type>
<position>201,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4758 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6658</ID>
<type>AE_DFF_LOW</type>
<position>214,-2119.5</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4759 </output>
<input>
<ID>clock</ID>4760 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6659</ID>
<type>BA_TRI_STATE</type>
<position>224,-2130</position>
<input>
<ID>ENABLE_0</ID>4761 </input>
<input>
<ID>IN_0</ID>4759 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6660</ID>
<type>AA_AND2</type>
<position>21.5,-2101.5</position>
<input>
<ID>IN_0</ID>4803 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4770 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6661</ID>
<type>BA_TRI_STATE</type>
<position>130,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4765 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6662</ID>
<type>AE_DFF_LOW</type>
<position>143,-2100.5</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4766 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6663</ID>
<type>BA_TRI_STATE</type>
<position>153,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4766 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6664</ID>
<type>AE_DFF_LOW</type>
<position>166,-2100.5</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4767 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6665</ID>
<type>BA_TRI_STATE</type>
<position>176,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4767 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6666</ID>
<type>AE_DFF_LOW</type>
<position>191,-2100.5</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4768 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6667</ID>
<type>BA_TRI_STATE</type>
<position>201,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4768 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6668</ID>
<type>AA_AND2</type>
<position>21.5,-1885.5</position>
<input>
<ID>IN_0</ID>4695 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4604 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6669</ID>
<type>AE_DFF_LOW</type>
<position>214,-2100.5</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4769 </output>
<input>
<ID>clock</ID>4770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6670</ID>
<type>BA_TRI_STATE</type>
<position>224,-2111</position>
<input>
<ID>ENABLE_0</ID>4771 </input>
<input>
<ID>IN_0</ID>4769 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6671</ID>
<type>AA_AND2</type>
<position>21.5,-2083</position>
<input>
<ID>IN_0</ID>4802 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4780 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6672</ID>
<type>AA_AND2</type>
<position>32.5,-2092.5</position>
<input>
<ID>IN_0</ID>4802 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6673</ID>
<type>AA_AND2</type>
<position>33,-1895</position>
<input>
<ID>IN_0</ID>4695 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4605 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6674</ID>
<type>AE_DFF_LOW</type>
<position>49,-2082</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4772 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6675</ID>
<type>BA_TRI_STATE</type>
<position>59,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4772 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6676</ID>
<type>AE_DFF_LOW</type>
<position>72,-2082</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4773 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6677</ID>
<type>BA_TRI_STATE</type>
<position>82,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4773 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6678</ID>
<type>AE_DFF_LOW</type>
<position>49,-1884.5</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4596 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6679</ID>
<type>AE_DFF_LOW</type>
<position>97,-2082</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4774 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6680</ID>
<type>BA_TRI_STATE</type>
<position>107,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4774 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6681</ID>
<type>AE_DFF_LOW</type>
<position>120,-2082</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4775 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6682</ID>
<type>BA_TRI_STATE</type>
<position>130,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4775 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6683</ID>
<type>AE_DFF_LOW</type>
<position>143,-2082</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4776 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6684</ID>
<type>BA_TRI_STATE</type>
<position>59,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4596 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6685</ID>
<type>BA_TRI_STATE</type>
<position>153,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4776 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6686</ID>
<type>AE_DFF_LOW</type>
<position>166,-2082</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4777 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6687</ID>
<type>BA_TRI_STATE</type>
<position>176,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4777 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6688</ID>
<type>AE_DFF_LOW</type>
<position>191,-2082</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4778 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6689</ID>
<type>BA_TRI_STATE</type>
<position>201,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4778 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6690</ID>
<type>AE_DFF_LOW</type>
<position>214,-2082</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4779 </output>
<input>
<ID>clock</ID>4780 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6691</ID>
<type>BA_TRI_STATE</type>
<position>224,-2092.5</position>
<input>
<ID>ENABLE_0</ID>4781 </input>
<input>
<ID>IN_0</ID>4779 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6692</ID>
<type>HA_JUNC_2</type>
<position>40.5,-1995.5</position>
<input>
<ID>N_in0</ID>4782 </input>
<input>
<ID>N_in1</ID>4810 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6693</ID>
<type>HA_JUNC_2</type>
<position>63.5,-1995</position>
<input>
<ID>N_in0</ID>4783 </input>
<input>
<ID>N_in1</ID>4811 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6694</ID>
<type>HA_JUNC_2</type>
<position>66.5,-1995.5</position>
<input>
<ID>N_in0</ID>4784 </input>
<input>
<ID>N_in1</ID>4812 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6695</ID>
<type>HA_JUNC_2</type>
<position>86,-1995</position>
<input>
<ID>N_in0</ID>4785 </input>
<input>
<ID>N_in1</ID>4813 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6696</ID>
<type>HA_JUNC_2</type>
<position>89.5,-1995</position>
<input>
<ID>N_in0</ID>4786 </input>
<input>
<ID>N_in1</ID>4814 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6697</ID>
<type>HA_JUNC_2</type>
<position>110.5,-1995.5</position>
<input>
<ID>N_in0</ID>4787 </input>
<input>
<ID>N_in1</ID>4815 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6698</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1995</position>
<input>
<ID>N_in0</ID>4788 </input>
<input>
<ID>N_in1</ID>4816 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6699</ID>
<type>HA_JUNC_2</type>
<position>133,-1995</position>
<input>
<ID>N_in0</ID>4789 </input>
<input>
<ID>N_in1</ID>4817 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6700</ID>
<type>AE_DFF_LOW</type>
<position>72,-1884.5</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4597 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6701</ID>
<type>HA_JUNC_2</type>
<position>137,-1995</position>
<input>
<ID>N_in0</ID>4790 </input>
<input>
<ID>N_in1</ID>4818 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6702</ID>
<type>BA_TRI_STATE</type>
<position>82,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4597 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6703</ID>
<type>HA_JUNC_2</type>
<position>156,-1995</position>
<input>
<ID>N_in0</ID>4791 </input>
<input>
<ID>N_in1</ID>4819 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6704</ID>
<type>AE_DFF_LOW</type>
<position>97,-1884.5</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4598 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6705</ID>
<type>HA_JUNC_2</type>
<position>161,-1995</position>
<input>
<ID>N_in0</ID>4792 </input>
<input>
<ID>N_in1</ID>4820 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6706</ID>
<type>BA_TRI_STATE</type>
<position>107,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4598 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6707</ID>
<type>HA_JUNC_2</type>
<position>183.5,-1995</position>
<input>
<ID>N_in0</ID>4794 </input>
<input>
<ID>N_in1</ID>4822 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6708</ID>
<type>AE_DFF_LOW</type>
<position>120,-1884.5</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4599 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6709</ID>
<type>HA_JUNC_2</type>
<position>179,-1995</position>
<input>
<ID>N_in0</ID>4793 </input>
<input>
<ID>N_in1</ID>4821 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6710</ID>
<type>BA_TRI_STATE</type>
<position>130,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4599 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6711</ID>
<type>HA_JUNC_2</type>
<position>204.5,-1995.5</position>
<input>
<ID>N_in0</ID>4795 </input>
<input>
<ID>N_in1</ID>4823 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6712</ID>
<type>AE_DFF_LOW</type>
<position>143,-1884.5</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4600 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6713</ID>
<type>HA_JUNC_2</type>
<position>229,-1996.5</position>
<input>
<ID>N_in0</ID>4797 </input>
<input>
<ID>N_in1</ID>4825 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6714</ID>
<type>BA_TRI_STATE</type>
<position>153,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4600 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6715</ID>
<type>AA_AND2</type>
<position>21.5,-2061</position>
<input>
<ID>IN_0</ID>4801 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4710 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6716</ID>
<type>AE_DFF_LOW</type>
<position>166,-1884.5</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4601 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6717</ID>
<type>AA_AND2</type>
<position>33,-2070.5</position>
<input>
<ID>IN_0</ID>4801 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4711 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6718</ID>
<type>BA_TRI_STATE</type>
<position>176,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4601 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6719</ID>
<type>HA_JUNC_2</type>
<position>40.5,-2162.5</position>
<input>
<ID>N_in1</ID>4782 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6720</ID>
<type>AE_DFF_LOW</type>
<position>191,-1884.5</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4602 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6721</ID>
<type>AE_DFF_LOW</type>
<position>49,-2060</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4702 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6722</ID>
<type>BA_TRI_STATE</type>
<position>201,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4602 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6723</ID>
<type>HA_JUNC_2</type>
<position>63.5,-2162</position>
<input>
<ID>N_in1</ID>4783 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6724</ID>
<type>AE_DFF_LOW</type>
<position>214,-1884.5</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4603 </output>
<input>
<ID>clock</ID>4604 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6725</ID>
<type>HA_JUNC_2</type>
<position>66.5,-2162</position>
<input>
<ID>N_in1</ID>4784 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6726</ID>
<type>BA_TRI_STATE</type>
<position>224,-1895</position>
<input>
<ID>ENABLE_0</ID>4605 </input>
<input>
<ID>IN_0</ID>4603 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6727</ID>
<type>HA_JUNC_2</type>
<position>86,-2162</position>
<input>
<ID>N_in1</ID>4785 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6728</ID>
<type>AA_AND2</type>
<position>21.5,-1867</position>
<input>
<ID>IN_0</ID>4694 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4614 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6729</ID>
<type>HA_JUNC_2</type>
<position>89.5,-2162</position>
<input>
<ID>N_in1</ID>4786 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6730</ID>
<type>AA_AND2</type>
<position>33,-1876.5</position>
<input>
<ID>IN_0</ID>4694 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4615 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6731</ID>
<type>HA_JUNC_2</type>
<position>110.5,-2162</position>
<input>
<ID>N_in1</ID>4787 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6732</ID>
<type>AE_DFF_LOW</type>
<position>49,-1866</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4606 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6733</ID>
<type>BA_TRI_STATE</type>
<position>59,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4702 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6734</ID>
<type>BA_TRI_STATE</type>
<position>59,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4606 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6735</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2162</position>
<input>
<ID>N_in1</ID>4788 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6736</ID>
<type>AE_DFF_LOW</type>
<position>72,-1866</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4607 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6737</ID>
<type>HA_JUNC_2</type>
<position>133,-2162</position>
<input>
<ID>N_in1</ID>4789 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6738</ID>
<type>BA_TRI_STATE</type>
<position>82,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4607 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6739</ID>
<type>HA_JUNC_2</type>
<position>137,-2162</position>
<input>
<ID>N_in1</ID>4790 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6740</ID>
<type>AE_DFF_LOW</type>
<position>97,-1866</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4608 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6741</ID>
<type>HA_JUNC_2</type>
<position>156,-2161.5</position>
<input>
<ID>N_in1</ID>4791 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6742</ID>
<type>BA_TRI_STATE</type>
<position>107,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4608 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6743</ID>
<type>HA_JUNC_2</type>
<position>161,-2161.5</position>
<input>
<ID>N_in1</ID>4792 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6744</ID>
<type>AE_DFF_LOW</type>
<position>120,-1866</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4609 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6745</ID>
<type>HA_JUNC_2</type>
<position>179,-2161</position>
<input>
<ID>N_in1</ID>4793 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6746</ID>
<type>BA_TRI_STATE</type>
<position>130,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4609 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6747</ID>
<type>HA_JUNC_2</type>
<position>183.5,-2161</position>
<input>
<ID>N_in1</ID>4794 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6748</ID>
<type>AE_DFF_LOW</type>
<position>143,-1866</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4610 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6749</ID>
<type>HA_JUNC_2</type>
<position>204.5,-2160.5</position>
<input>
<ID>N_in1</ID>4795 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6750</ID>
<type>BA_TRI_STATE</type>
<position>153,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4610 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6751</ID>
<type>HA_JUNC_2</type>
<position>208,-2160.5</position>
<input>
<ID>N_in1</ID>4796 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6752</ID>
<type>AE_DFF_LOW</type>
<position>166,-1866</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4611 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6753</ID>
<type>HA_JUNC_2</type>
<position>208,-1995.5</position>
<input>
<ID>N_in0</ID>4796 </input>
<input>
<ID>N_in1</ID>4824 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6754</ID>
<type>BA_TRI_STATE</type>
<position>176,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4611 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6755</ID>
<type>HA_JUNC_2</type>
<position>229,-2160.5</position>
<input>
<ID>N_in1</ID>4797 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6756</ID>
<type>AE_DFF_LOW</type>
<position>191,-1866</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4612 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6757</ID>
<type>AE_DFF_LOW</type>
<position>72,-2060</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4703 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6758</ID>
<type>BA_TRI_STATE</type>
<position>201,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4612 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6759</ID>
<type>BA_TRI_STATE</type>
<position>82,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4703 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6760</ID>
<type>AE_DFF_LOW</type>
<position>214,-1866</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4613 </output>
<input>
<ID>clock</ID>4614 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6761</ID>
<type>HA_JUNC_2</type>
<position>27.5,-1995.5</position>
<input>
<ID>N_in0</ID>4807 </input>
<input>
<ID>N_in1</ID>4809 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6762</ID>
<type>BA_TRI_STATE</type>
<position>224,-1876.5</position>
<input>
<ID>ENABLE_0</ID>4615 </input>
<input>
<ID>IN_0</ID>4613 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6763</ID>
<type>AE_DFF_LOW</type>
<position>97,-2060</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4704 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6764</ID>
<type>AA_AND2</type>
<position>21.5,-1848</position>
<input>
<ID>IN_0</ID>4693 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4624 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6765</ID>
<type>HA_JUNC_2</type>
<position>17.5,-1995.5</position>
<input>
<ID>N_in0</ID>4806 </input>
<input>
<ID>N_in1</ID>4808 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6766</ID>
<type>AA_AND2</type>
<position>33,-1857.5</position>
<input>
<ID>IN_0</ID>4693 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6767</ID>
<type>BA_TRI_STATE</type>
<position>107,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4704 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6768</ID>
<type>AE_DFF_LOW</type>
<position>49,-1847</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4616 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6769</ID>
<type>HA_JUNC_2</type>
<position>27.5,-2162.5</position>
<input>
<ID>N_in1</ID>4807 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6770</ID>
<type>BA_TRI_STATE</type>
<position>59,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4616 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6771</ID>
<type>AE_DFF_LOW</type>
<position>120,-2060</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4705 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6772</ID>
<type>AE_DFF_LOW</type>
<position>72,-1847</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4617 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6773</ID>
<type>HA_JUNC_2</type>
<position>17.5,-2162.5</position>
<input>
<ID>N_in1</ID>4806 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6774</ID>
<type>BA_TRI_STATE</type>
<position>82,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4617 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6775</ID>
<type>BA_TRI_STATE</type>
<position>130,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4705 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6776</ID>
<type>AE_DFF_LOW</type>
<position>97,-1847</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4618 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6777</ID>
<type>AE_DFF_LOW</type>
<position>143,-2060</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4706 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6778</ID>
<type>BA_TRI_STATE</type>
<position>107,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4618 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6779</ID>
<type>AA_LABEL</type>
<position>8.5,-1996</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6780</ID>
<type>AE_DFF_LOW</type>
<position>120,-1847</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4619 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6781</ID>
<type>BA_TRI_STATE</type>
<position>153,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4706 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6782</ID>
<type>BA_TRI_STATE</type>
<position>130,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4619 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6783</ID>
<type>AE_DFF_LOW</type>
<position>166,-2060</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4707 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6784</ID>
<type>AE_DFF_LOW</type>
<position>143,-1847</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4620 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6785</ID>
<type>BA_TRI_STATE</type>
<position>176,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4707 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6786</ID>
<type>BA_TRI_STATE</type>
<position>153,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4620 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6787</ID>
<type>AE_DFF_LOW</type>
<position>191,-2060</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4708 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6788</ID>
<type>AE_DFF_LOW</type>
<position>166,-1847</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4621 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6789</ID>
<type>BA_TRI_STATE</type>
<position>201,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4708 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6790</ID>
<type>BA_TRI_STATE</type>
<position>176,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4621 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6791</ID>
<type>AE_DFF_LOW</type>
<position>214,-2060</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4709 </output>
<input>
<ID>clock</ID>4710 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6792</ID>
<type>AE_DFF_LOW</type>
<position>191,-1847</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4622 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6793</ID>
<type>BA_TRI_STATE</type>
<position>224,-2070.5</position>
<input>
<ID>ENABLE_0</ID>4711 </input>
<input>
<ID>IN_0</ID>4709 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6794</ID>
<type>BA_TRI_STATE</type>
<position>201,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4622 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6795</ID>
<type>AA_AND2</type>
<position>21.5,-2042.5</position>
<input>
<ID>IN_0</ID>4800 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4720 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6796</ID>
<type>AE_DFF_LOW</type>
<position>214,-1847</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4623 </output>
<input>
<ID>clock</ID>4624 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6797</ID>
<type>AA_AND2</type>
<position>33,-2052</position>
<input>
<ID>IN_0</ID>4800 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4721 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6798</ID>
<type>BA_TRI_STATE</type>
<position>224,-1857.5</position>
<input>
<ID>ENABLE_0</ID>4625 </input>
<input>
<ID>IN_0</ID>4623 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6799</ID>
<type>AE_DFF_LOW</type>
<position>49,-2041.5</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4712 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6800</ID>
<type>AA_AND2</type>
<position>21.5,-1829.5</position>
<input>
<ID>IN_0</ID>4692 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4634 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6801</ID>
<type>BA_TRI_STATE</type>
<position>59,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4712 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6802</ID>
<type>AA_AND2</type>
<position>33,-1839</position>
<input>
<ID>IN_0</ID>4692 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4635 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6803</ID>
<type>AE_DFF_LOW</type>
<position>72,-2041.5</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4713 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6804</ID>
<type>AE_DFF_LOW</type>
<position>49,-1828.5</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4626 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6805</ID>
<type>BA_TRI_STATE</type>
<position>82,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4713 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6806</ID>
<type>BA_TRI_STATE</type>
<position>59,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4626 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6807</ID>
<type>AE_DFF_LOW</type>
<position>97,-2041.5</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4714 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6808</ID>
<type>AE_DFF_LOW</type>
<position>72,-1828.5</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4627 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6809</ID>
<type>BA_TRI_STATE</type>
<position>107,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4714 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6810</ID>
<type>BA_TRI_STATE</type>
<position>82,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4627 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6811</ID>
<type>AE_DFF_LOW</type>
<position>120,-2041.5</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4715 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6812</ID>
<type>AE_DFF_LOW</type>
<position>97,-1828.5</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4628 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6813</ID>
<type>BA_TRI_STATE</type>
<position>130,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4715 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6814</ID>
<type>BA_TRI_STATE</type>
<position>107,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4628 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6815</ID>
<type>AE_DFF_LOW</type>
<position>143,-2041.5</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4716 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6816</ID>
<type>AE_DFF_LOW</type>
<position>120,-1828.5</position>
<input>
<ID>IN_0</ID>4682 </input>
<output>
<ID>OUT_0</ID>4629 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6817</ID>
<type>BA_TRI_STATE</type>
<position>153,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4716 </input>
<output>
<ID>OUT_0</ID>4791 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6818</ID>
<type>BA_TRI_STATE</type>
<position>130,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4629 </input>
<output>
<ID>OUT_0</ID>4683 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6819</ID>
<type>AE_DFF_LOW</type>
<position>166,-2041.5</position>
<input>
<ID>IN_0</ID>4792 </input>
<output>
<ID>OUT_0</ID>4717 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6820</ID>
<type>AE_DFF_LOW</type>
<position>143,-1828.5</position>
<input>
<ID>IN_0</ID>4684 </input>
<output>
<ID>OUT_0</ID>4630 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6821</ID>
<type>BA_TRI_STATE</type>
<position>176,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4717 </input>
<output>
<ID>OUT_0</ID>4793 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6822</ID>
<type>BA_TRI_STATE</type>
<position>153,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4630 </input>
<output>
<ID>OUT_0</ID>4685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6823</ID>
<type>AE_DFF_LOW</type>
<position>191,-2041.5</position>
<input>
<ID>IN_0</ID>4794 </input>
<output>
<ID>OUT_0</ID>4718 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6824</ID>
<type>AE_DFF_LOW</type>
<position>166,-1828.5</position>
<input>
<ID>IN_0</ID>4686 </input>
<output>
<ID>OUT_0</ID>4631 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6825</ID>
<type>BA_TRI_STATE</type>
<position>201,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4718 </input>
<output>
<ID>OUT_0</ID>4795 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6826</ID>
<type>BA_TRI_STATE</type>
<position>176,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4631 </input>
<output>
<ID>OUT_0</ID>4687 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6827</ID>
<type>AE_DFF_LOW</type>
<position>214,-2041.5</position>
<input>
<ID>IN_0</ID>4796 </input>
<output>
<ID>OUT_0</ID>4719 </output>
<input>
<ID>clock</ID>4720 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6828</ID>
<type>AE_DFF_LOW</type>
<position>191,-1828.5</position>
<input>
<ID>IN_0</ID>4688 </input>
<output>
<ID>OUT_0</ID>4632 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6829</ID>
<type>BA_TRI_STATE</type>
<position>224,-2052</position>
<input>
<ID>ENABLE_0</ID>4721 </input>
<input>
<ID>IN_0</ID>4719 </input>
<output>
<ID>OUT_0</ID>4797 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6830</ID>
<type>BA_TRI_STATE</type>
<position>201,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4632 </input>
<output>
<ID>OUT_0</ID>4689 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6831</ID>
<type>AA_AND2</type>
<position>21.5,-2023.5</position>
<input>
<ID>IN_0</ID>4799 </input>
<input>
<ID>IN_1</ID>4806 </input>
<output>
<ID>OUT</ID>4730 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6832</ID>
<type>AE_DFF_LOW</type>
<position>214,-1828.5</position>
<input>
<ID>IN_0</ID>4690 </input>
<output>
<ID>OUT_0</ID>4633 </output>
<input>
<ID>clock</ID>4634 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6833</ID>
<type>AA_AND2</type>
<position>33,-2033</position>
<input>
<ID>IN_0</ID>4799 </input>
<input>
<ID>IN_1</ID>4807 </input>
<output>
<ID>OUT</ID>4731 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6834</ID>
<type>BA_TRI_STATE</type>
<position>224,-1839</position>
<input>
<ID>ENABLE_0</ID>4635 </input>
<input>
<ID>IN_0</ID>4633 </input>
<output>
<ID>OUT_0</ID>4691 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6835</ID>
<type>AE_DFF_LOW</type>
<position>49,-2022.5</position>
<input>
<ID>IN_0</ID>4782 </input>
<output>
<ID>OUT_0</ID>4722 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6836</ID>
<type>AA_AND2</type>
<position>21.5,-1963.5</position>
<input>
<ID>IN_0</ID>4699 </input>
<input>
<ID>IN_1</ID>4700 </input>
<output>
<ID>OUT</ID>4644 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6837</ID>
<type>BA_TRI_STATE</type>
<position>59,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4722 </input>
<output>
<ID>OUT_0</ID>4783 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6838</ID>
<type>AA_AND2</type>
<position>32.5,-1973</position>
<input>
<ID>IN_0</ID>4699 </input>
<input>
<ID>IN_1</ID>4701 </input>
<output>
<ID>OUT</ID>4645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6839</ID>
<type>AE_DFF_LOW</type>
<position>72,-2022.5</position>
<input>
<ID>IN_0</ID>4784 </input>
<output>
<ID>OUT_0</ID>4723 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6840</ID>
<type>AE_DFF_LOW</type>
<position>49,-1962.5</position>
<input>
<ID>IN_0</ID>4676 </input>
<output>
<ID>OUT_0</ID>4636 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6841</ID>
<type>BA_TRI_STATE</type>
<position>82,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4723 </input>
<output>
<ID>OUT_0</ID>4785 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6842</ID>
<type>BA_TRI_STATE</type>
<position>59,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4636 </input>
<output>
<ID>OUT_0</ID>4677 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6843</ID>
<type>AE_DFF_LOW</type>
<position>97,-2022.5</position>
<input>
<ID>IN_0</ID>4786 </input>
<output>
<ID>OUT_0</ID>4724 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6844</ID>
<type>AE_DFF_LOW</type>
<position>72,-1962.5</position>
<input>
<ID>IN_0</ID>4678 </input>
<output>
<ID>OUT_0</ID>4637 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6845</ID>
<type>BA_TRI_STATE</type>
<position>107,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4724 </input>
<output>
<ID>OUT_0</ID>4787 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6846</ID>
<type>BA_TRI_STATE</type>
<position>82,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4637 </input>
<output>
<ID>OUT_0</ID>4679 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6847</ID>
<type>AE_DFF_LOW</type>
<position>120,-2022.5</position>
<input>
<ID>IN_0</ID>4788 </input>
<output>
<ID>OUT_0</ID>4725 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6848</ID>
<type>AE_DFF_LOW</type>
<position>97,-1962.5</position>
<input>
<ID>IN_0</ID>4680 </input>
<output>
<ID>OUT_0</ID>4638 </output>
<input>
<ID>clock</ID>4644 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6849</ID>
<type>BA_TRI_STATE</type>
<position>130,-2033</position>
<input>
<ID>ENABLE_0</ID>4731 </input>
<input>
<ID>IN_0</ID>4725 </input>
<output>
<ID>OUT_0</ID>4789 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6850</ID>
<type>BA_TRI_STATE</type>
<position>107,-1973</position>
<input>
<ID>ENABLE_0</ID>4645 </input>
<input>
<ID>IN_0</ID>4638 </input>
<output>
<ID>OUT_0</ID>4681 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6851</ID>
<type>AE_DFF_LOW</type>
<position>143,-2022.5</position>
<input>
<ID>IN_0</ID>4790 </input>
<output>
<ID>OUT_0</ID>4726 </output>
<input>
<ID>clock</ID>4730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6853</ID>
<type>AA_LABEL</type>
<position>261,-1985.5</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6854</ID>
<type>AE_DFF_LOW</type>
<position>120,-2322.5</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4869 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6855</ID>
<type>BA_TRI_STATE</type>
<position>153,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4956 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6856</ID>
<type>BA_TRI_STATE</type>
<position>130,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4869 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6857</ID>
<type>AE_DFF_LOW</type>
<position>166,-2382.5</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4957 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6858</ID>
<type>AE_DFF_LOW</type>
<position>143,-2322.5</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4870 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6859</ID>
<type>BA_TRI_STATE</type>
<position>176,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4957 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6860</ID>
<type>BA_TRI_STATE</type>
<position>153,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4870 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6861</ID>
<type>AE_DFF_LOW</type>
<position>191,-2382.5</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4958 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6862</ID>
<type>AE_DFF_LOW</type>
<position>166,-2322.5</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4871 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6863</ID>
<type>BA_TRI_STATE</type>
<position>201,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4958 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6864</ID>
<type>BA_TRI_STATE</type>
<position>176,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4871 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6865</ID>
<type>AE_DFF_LOW</type>
<position>214,-2382.5</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4959 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6866</ID>
<type>AE_DFF_LOW</type>
<position>191,-2322.5</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4872 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6867</ID>
<type>BA_TRI_STATE</type>
<position>224,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4959 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6868</ID>
<type>BA_TRI_STATE</type>
<position>201,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4872 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6869</ID>
<type>AA_AND2</type>
<position>21.5,-2365</position>
<input>
<ID>IN_0</ID>5028 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>4970 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6870</ID>
<type>AE_DFF_LOW</type>
<position>214,-2322.5</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4873 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6871</ID>
<type>AA_AND2</type>
<position>33,-2374.5</position>
<input>
<ID>IN_0</ID>5028 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>4971 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6872</ID>
<type>BA_TRI_STATE</type>
<position>224,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4873 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6873</ID>
<type>AE_DFF_LOW</type>
<position>49,-2364</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4962 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6874</ID>
<type>AA_AND2</type>
<position>21.5,-2305</position>
<input>
<ID>IN_0</ID>4928 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6875</ID>
<type>BA_TRI_STATE</type>
<position>59,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4962 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6876</ID>
<type>AA_AND2</type>
<position>32.5,-2314.5</position>
<input>
<ID>IN_0</ID>4928 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4885 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6877</ID>
<type>AE_DFF_LOW</type>
<position>72,-2364</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4963 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6878</ID>
<type>AE_DFF_LOW</type>
<position>49,-2304</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4876 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6879</ID>
<type>BA_TRI_STATE</type>
<position>82,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4963 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6880</ID>
<type>BA_TRI_STATE</type>
<position>59,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4876 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6881</ID>
<type>AE_DFF_LOW</type>
<position>97,-2364</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4964 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6882</ID>
<type>AE_DFF_LOW</type>
<position>72,-2304</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4877 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6883</ID>
<type>BA_TRI_STATE</type>
<position>107,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4964 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6884</ID>
<type>BA_TRI_STATE</type>
<position>82,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4877 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6885</ID>
<type>AE_DFF_LOW</type>
<position>120,-2364</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4965 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6886</ID>
<type>AE_DFF_LOW</type>
<position>97,-2304</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4878 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6887</ID>
<type>BA_TRI_STATE</type>
<position>130,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4965 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6888</ID>
<type>BA_TRI_STATE</type>
<position>107,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4878 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6889</ID>
<type>AE_DFF_LOW</type>
<position>143,-2364</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4966 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6890</ID>
<type>AE_DFF_LOW</type>
<position>120,-2304</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4879 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6891</ID>
<type>BA_TRI_STATE</type>
<position>153,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4966 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6892</ID>
<type>BA_TRI_STATE</type>
<position>130,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4879 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6893</ID>
<type>AE_DFF_LOW</type>
<position>166,-2364</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4967 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6894</ID>
<type>AE_DFF_LOW</type>
<position>143,-2304</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4880 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6895</ID>
<type>BA_TRI_STATE</type>
<position>176,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4967 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6896</ID>
<type>BA_TRI_STATE</type>
<position>153,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4880 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6897</ID>
<type>AE_DFF_LOW</type>
<position>191,-2364</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4968 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6898</ID>
<type>AE_DFF_LOW</type>
<position>166,-2304</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4881 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6899</ID>
<type>BA_TRI_STATE</type>
<position>201,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4968 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6900</ID>
<type>BA_TRI_STATE</type>
<position>176,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4881 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6901</ID>
<type>AE_DFF_LOW</type>
<position>214,-2364</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4969 </output>
<input>
<ID>clock</ID>4970 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6902</ID>
<type>AE_DFF_LOW</type>
<position>191,-2304</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4882 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6903</ID>
<type>BA_TRI_STATE</type>
<position>224,-2374.5</position>
<input>
<ID>ENABLE_0</ID>4971 </input>
<input>
<ID>IN_0</ID>4969 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6904</ID>
<type>BA_TRI_STATE</type>
<position>201,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4882 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6905</ID>
<type>AA_AND2</type>
<position>21.5,-2499</position>
<input>
<ID>IN_0</ID>5035 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>4980 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6906</ID>
<type>AE_DFF_LOW</type>
<position>214,-2304</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4883 </output>
<input>
<ID>clock</ID>4884 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6907</ID>
<type>AA_AND2</type>
<position>32.5,-2508.5</position>
<input>
<ID>IN_0</ID>5035 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>4981 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6908</ID>
<type>BA_TRI_STATE</type>
<position>224,-2314.5</position>
<input>
<ID>ENABLE_0</ID>4885 </input>
<input>
<ID>IN_0</ID>4883 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6909</ID>
<type>AE_DFF_LOW</type>
<position>49,-2498</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4972 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6910</ID>
<type>AA_AND2</type>
<position>32.5,-2471</position>
<input>
<ID>IN_0</ID>5033 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>5001 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6911</ID>
<type>AA_AND2</type>
<position>21.5,-2286</position>
<input>
<ID>IN_0</ID>4927 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4894 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6912</ID>
<type>BA_TRI_STATE</type>
<position>59,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4972 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6913</ID>
<type>AA_AND2</type>
<position>32.5,-2295.5</position>
<input>
<ID>IN_0</ID>4927 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4895 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6914</ID>
<type>AE_DFF_LOW</type>
<position>72,-2498</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4973 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6915</ID>
<type>AE_DFF_LOW</type>
<position>49,-2460.5</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4992 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6916</ID>
<type>AE_DFF_LOW</type>
<position>49,-2285</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4886 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6917</ID>
<type>BA_TRI_STATE</type>
<position>82,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4973 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6918</ID>
<type>BA_TRI_STATE</type>
<position>59,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4886 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6919</ID>
<type>AE_DFF_LOW</type>
<position>97,-2498</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4974 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6920</ID>
<type>BA_TRI_STATE</type>
<position>59,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4992 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6921</ID>
<type>AE_DFF_LOW</type>
<position>72,-2285</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4887 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6922</ID>
<type>BA_TRI_STATE</type>
<position>107,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4974 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6923</ID>
<type>BA_TRI_STATE</type>
<position>82,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4887 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6924</ID>
<type>AE_DFF_LOW</type>
<position>120,-2498</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4975 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6925</ID>
<type>AE_DFF_LOW</type>
<position>72,-2460.5</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4993 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6926</ID>
<type>AE_DFF_LOW</type>
<position>97,-2285</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4888 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6927</ID>
<type>BA_TRI_STATE</type>
<position>130,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4975 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6928</ID>
<type>BA_TRI_STATE</type>
<position>107,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4888 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6929</ID>
<type>AE_DFF_LOW</type>
<position>143,-2498</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4976 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6930</ID>
<type>BA_TRI_STATE</type>
<position>82,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4993 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6931</ID>
<type>AE_DFF_LOW</type>
<position>120,-2285</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4889 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6932</ID>
<type>BA_TRI_STATE</type>
<position>153,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4976 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6933</ID>
<type>BA_TRI_STATE</type>
<position>130,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4889 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6934</ID>
<type>AE_DFF_LOW</type>
<position>166,-2498</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4977 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6935</ID>
<type>AE_DFF_LOW</type>
<position>97,-2460.5</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4994 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6936</ID>
<type>AE_DFF_LOW</type>
<position>143,-2285</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4890 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6937</ID>
<type>BA_TRI_STATE</type>
<position>176,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4977 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6938</ID>
<type>BA_TRI_STATE</type>
<position>153,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4890 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6939</ID>
<type>BA_TRI_STATE</type>
<position>107,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4994 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6940</ID>
<type>AE_DFF_LOW</type>
<position>166,-2285</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4891 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6941</ID>
<type>BA_TRI_STATE</type>
<position>176,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4891 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6942</ID>
<type>AE_DFF_LOW</type>
<position>120,-2460.5</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4995 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6943</ID>
<type>AE_DFF_LOW</type>
<position>191,-2285</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4892 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6944</ID>
<type>BA_TRI_STATE</type>
<position>201,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4892 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6945</ID>
<type>AE_DFF_LOW</type>
<position>214,-2285</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4893 </output>
<input>
<ID>clock</ID>4894 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6946</ID>
<type>BA_TRI_STATE</type>
<position>224,-2295.5</position>
<input>
<ID>ENABLE_0</ID>4895 </input>
<input>
<ID>IN_0</ID>4893 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6947</ID>
<type>AA_AND2</type>
<position>21.5,-2267.5</position>
<input>
<ID>IN_0</ID>4926 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4904 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6948</ID>
<type>AA_AND2</type>
<position>32.5,-2277</position>
<input>
<ID>IN_0</ID>4926 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4905 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6949</ID>
<type>AE_DFF_LOW</type>
<position>49,-2266.5</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4896 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6950</ID>
<type>BA_TRI_STATE</type>
<position>59,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4896 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6951</ID>
<type>AE_DFF_LOW</type>
<position>72,-2266.5</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4897 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6952</ID>
<type>BA_TRI_STATE</type>
<position>82,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4897 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6953</ID>
<type>AE_DFF_LOW</type>
<position>97,-2266.5</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4898 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6954</ID>
<type>BA_TRI_STATE</type>
<position>107,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4898 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6955</ID>
<type>AE_DFF_LOW</type>
<position>120,-2266.5</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4899 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6956</ID>
<type>BA_TRI_STATE</type>
<position>130,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4899 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6957</ID>
<type>AE_DFF_LOW</type>
<position>143,-2266.5</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4900 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6958</ID>
<type>BA_TRI_STATE</type>
<position>153,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4900 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6959</ID>
<type>AE_DFF_LOW</type>
<position>166,-2266.5</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4901 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6960</ID>
<type>BA_TRI_STATE</type>
<position>176,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4901 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6961</ID>
<type>AE_DFF_LOW</type>
<position>191,-2266.5</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4902 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6962</ID>
<type>BA_TRI_STATE</type>
<position>201,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4902 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6963</ID>
<type>AE_DFF_LOW</type>
<position>214,-2266.5</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4903 </output>
<input>
<ID>clock</ID>4904 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6964</ID>
<type>BA_TRI_STATE</type>
<position>224,-2277</position>
<input>
<ID>ENABLE_0</ID>4905 </input>
<input>
<ID>IN_0</ID>4903 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6965</ID>
<type>HA_JUNC_2</type>
<position>40.5,-2180</position>
<input>
<ID>N_in0</ID>4906 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6966</ID>
<type>HA_JUNC_2</type>
<position>63.5,-2179.5</position>
<input>
<ID>N_in0</ID>4907 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6967</ID>
<type>HA_JUNC_2</type>
<position>66.5,-2180</position>
<input>
<ID>N_in0</ID>4908 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6968</ID>
<type>HA_JUNC_2</type>
<position>86,-2179.5</position>
<input>
<ID>N_in0</ID>4909 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6969</ID>
<type>HA_JUNC_2</type>
<position>89.5,-2179.5</position>
<input>
<ID>N_in0</ID>4910 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6970</ID>
<type>HA_JUNC_2</type>
<position>110.5,-2180</position>
<input>
<ID>N_in0</ID>4911 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6971</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2179.5</position>
<input>
<ID>N_in0</ID>4912 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6972</ID>
<type>HA_JUNC_2</type>
<position>133,-2179.5</position>
<input>
<ID>N_in0</ID>4913 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6973</ID>
<type>HA_JUNC_2</type>
<position>137,-2179.5</position>
<input>
<ID>N_in0</ID>4914 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6974</ID>
<type>HA_JUNC_2</type>
<position>156,-2179.5</position>
<input>
<ID>N_in0</ID>4915 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6975</ID>
<type>HA_JUNC_2</type>
<position>161,-2179.5</position>
<input>
<ID>N_in0</ID>4916 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6976</ID>
<type>HA_JUNC_2</type>
<position>183.5,-2179.5</position>
<input>
<ID>N_in0</ID>4918 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6977</ID>
<type>HA_JUNC_2</type>
<position>179,-2179.5</position>
<input>
<ID>N_in0</ID>4917 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6978</ID>
<type>HA_JUNC_2</type>
<position>204.5,-2180</position>
<input>
<ID>N_in0</ID>4919 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6979</ID>
<type>HA_JUNC_2</type>
<position>229,-2181</position>
<input>
<ID>N_in0</ID>4921 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6980</ID>
<type>HA_JUNC_2</type>
<position>40.5,-2347</position>
<input>
<ID>N_in0</ID>5040 </input>
<input>
<ID>N_in1</ID>4906 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6981</ID>
<type>HA_JUNC_2</type>
<position>63.5,-2346.5</position>
<input>
<ID>N_in0</ID>5041 </input>
<input>
<ID>N_in1</ID>4907 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6982</ID>
<type>HA_JUNC_2</type>
<position>66.5,-2346.5</position>
<input>
<ID>N_in0</ID>5042 </input>
<input>
<ID>N_in1</ID>4908 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6983</ID>
<type>HA_JUNC_2</type>
<position>86,-2346.5</position>
<input>
<ID>N_in0</ID>5043 </input>
<input>
<ID>N_in1</ID>4909 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6984</ID>
<type>HA_JUNC_2</type>
<position>89.5,-2346.5</position>
<input>
<ID>N_in0</ID>5044 </input>
<input>
<ID>N_in1</ID>4910 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6985</ID>
<type>HA_JUNC_2</type>
<position>110.5,-2346.5</position>
<input>
<ID>N_in0</ID>5045 </input>
<input>
<ID>N_in1</ID>4911 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6986</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2346.5</position>
<input>
<ID>N_in0</ID>5046 </input>
<input>
<ID>N_in1</ID>4912 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6987</ID>
<type>HA_JUNC_2</type>
<position>133,-2346.5</position>
<input>
<ID>N_in0</ID>5047 </input>
<input>
<ID>N_in1</ID>4913 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6988</ID>
<type>HA_JUNC_2</type>
<position>137,-2346.5</position>
<input>
<ID>N_in0</ID>5048 </input>
<input>
<ID>N_in1</ID>4914 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6989</ID>
<type>HA_JUNC_2</type>
<position>156,-2346</position>
<input>
<ID>N_in0</ID>5049 </input>
<input>
<ID>N_in1</ID>4915 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6990</ID>
<type>HA_JUNC_2</type>
<position>161,-2346</position>
<input>
<ID>N_in0</ID>5050 </input>
<input>
<ID>N_in1</ID>4916 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6991</ID>
<type>HA_JUNC_2</type>
<position>179,-2345.5</position>
<input>
<ID>N_in0</ID>5051 </input>
<input>
<ID>N_in1</ID>4917 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6992</ID>
<type>HA_JUNC_2</type>
<position>183.5,-2345.5</position>
<input>
<ID>N_in0</ID>5052 </input>
<input>
<ID>N_in1</ID>4918 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6993</ID>
<type>HA_JUNC_2</type>
<position>204.5,-2345</position>
<input>
<ID>N_in0</ID>5053 </input>
<input>
<ID>N_in1</ID>4919 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6994</ID>
<type>HA_JUNC_2</type>
<position>208,-2345</position>
<input>
<ID>N_in0</ID>5054 </input>
<input>
<ID>N_in1</ID>4920 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6995</ID>
<type>HA_JUNC_2</type>
<position>208,-2180</position>
<input>
<ID>N_in0</ID>4920 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6996</ID>
<type>HA_JUNC_2</type>
<position>229,-2345</position>
<input>
<ID>N_in0</ID>5055 </input>
<input>
<ID>N_in1</ID>4921 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6997</ID>
<type>HA_JUNC_2</type>
<position>27.5,-2180</position>
<input>
<ID>N_in0</ID>4931 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6998</ID>
<type>HA_JUNC_2</type>
<position>17.5,-2180</position>
<input>
<ID>N_in0</ID>4930 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6999</ID>
<type>HA_JUNC_2</type>
<position>27.5,-2347</position>
<input>
<ID>N_in0</ID>5039 </input>
<input>
<ID>N_in1</ID>4931 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7000</ID>
<type>HA_JUNC_2</type>
<position>17.5,-2347</position>
<input>
<ID>N_in0</ID>5038 </input>
<input>
<ID>N_in1</ID>4930 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7001</ID>
<type>AA_LABEL</type>
<position>8.5,-2180.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7002</ID>
<type>BI_DECODER_4x16</type>
<position>-131,-2347.5</position>
<output>
<ID>OUT_0</ID>5035 </output>
<output>
<ID>OUT_1</ID>5034 </output>
<output>
<ID>OUT_10</ID>4927 </output>
<output>
<ID>OUT_11</ID>4926 </output>
<output>
<ID>OUT_12</ID>4925 </output>
<output>
<ID>OUT_13</ID>4924 </output>
<output>
<ID>OUT_14</ID>4923 </output>
<output>
<ID>OUT_15</ID>4922 </output>
<output>
<ID>OUT_2</ID>5033 </output>
<output>
<ID>OUT_3</ID>5032 </output>
<output>
<ID>OUT_4</ID>5031 </output>
<output>
<ID>OUT_5</ID>5030 </output>
<output>
<ID>OUT_6</ID>5029 </output>
<output>
<ID>OUT_7</ID>5028 </output>
<output>
<ID>OUT_8</ID>4929 </output>
<output>
<ID>OUT_9</ID>4928 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7003</ID>
<type>AE_DFF_LOW</type>
<position>191,-2498</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4978 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7004</ID>
<type>BA_TRI_STATE</type>
<position>201,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4978 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7005</ID>
<type>AE_DFF_LOW</type>
<position>214,-2498</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4979 </output>
<input>
<ID>clock</ID>4980 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7006</ID>
<type>BA_TRI_STATE</type>
<position>224,-2508.5</position>
<input>
<ID>ENABLE_0</ID>4981 </input>
<input>
<ID>IN_0</ID>4979 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7007</ID>
<type>AA_AND2</type>
<position>21.5,-2480.5</position>
<input>
<ID>IN_0</ID>5034 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>4990 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7008</ID>
<type>AA_AND2</type>
<position>32.5,-2490</position>
<input>
<ID>IN_0</ID>5034 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>4991 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7009</ID>
<type>AE_DFF_LOW</type>
<position>49,-2479.5</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4982 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7010</ID>
<type>BA_TRI_STATE</type>
<position>59,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4982 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7011</ID>
<type>AE_DFF_LOW</type>
<position>72,-2479.5</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4983 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7012</ID>
<type>BA_TRI_STATE</type>
<position>82,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4983 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7013</ID>
<type>AE_DFF_LOW</type>
<position>97,-2479.5</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4984 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7014</ID>
<type>BA_TRI_STATE</type>
<position>107,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4984 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7015</ID>
<type>AE_DFF_LOW</type>
<position>120,-2479.5</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4985 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7016</ID>
<type>BA_TRI_STATE</type>
<position>130,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4985 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7017</ID>
<type>AE_DFF_LOW</type>
<position>143,-2479.5</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4986 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7018</ID>
<type>BA_TRI_STATE</type>
<position>153,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4986 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7019</ID>
<type>AE_DFF_LOW</type>
<position>166,-2479.5</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4987 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7020</ID>
<type>BA_TRI_STATE</type>
<position>176,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4987 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7021</ID>
<type>AE_DFF_LOW</type>
<position>191,-2479.5</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4988 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7022</ID>
<type>BA_TRI_STATE</type>
<position>201,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4988 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7023</ID>
<type>AE_DFF_LOW</type>
<position>214,-2479.5</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4989 </output>
<input>
<ID>clock</ID>4990 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7024</ID>
<type>BA_TRI_STATE</type>
<position>224,-2490</position>
<input>
<ID>ENABLE_0</ID>4991 </input>
<input>
<ID>IN_0</ID>4989 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7025</ID>
<type>AA_AND2</type>
<position>21.5,-2461.5</position>
<input>
<ID>IN_0</ID>5033 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>5000 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7026</ID>
<type>BA_TRI_STATE</type>
<position>130,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4995 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7027</ID>
<type>AE_DFF_LOW</type>
<position>143,-2460.5</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4996 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7028</ID>
<type>BA_TRI_STATE</type>
<position>153,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4996 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7029</ID>
<type>AE_DFF_LOW</type>
<position>166,-2460.5</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4997 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7030</ID>
<type>BA_TRI_STATE</type>
<position>176,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4997 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7031</ID>
<type>AE_DFF_LOW</type>
<position>191,-2460.5</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4998 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7032</ID>
<type>BA_TRI_STATE</type>
<position>201,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4998 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7033</ID>
<type>AA_AND2</type>
<position>21.5,-2245.5</position>
<input>
<ID>IN_0</ID>4925 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4834 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7034</ID>
<type>AE_DFF_LOW</type>
<position>214,-2460.5</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4999 </output>
<input>
<ID>clock</ID>5000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7035</ID>
<type>BA_TRI_STATE</type>
<position>224,-2471</position>
<input>
<ID>ENABLE_0</ID>5001 </input>
<input>
<ID>IN_0</ID>4999 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7036</ID>
<type>AA_AND2</type>
<position>21.5,-2443</position>
<input>
<ID>IN_0</ID>5032 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>5010 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7037</ID>
<type>AA_AND2</type>
<position>32.5,-2452.5</position>
<input>
<ID>IN_0</ID>5032 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>5011 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7038</ID>
<type>AA_AND2</type>
<position>33,-2255</position>
<input>
<ID>IN_0</ID>4925 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4835 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7039</ID>
<type>AE_DFF_LOW</type>
<position>49,-2442</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>5002 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7040</ID>
<type>BA_TRI_STATE</type>
<position>59,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5002 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7041</ID>
<type>AE_DFF_LOW</type>
<position>72,-2442</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>5003 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7042</ID>
<type>BA_TRI_STATE</type>
<position>82,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5003 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7043</ID>
<type>AE_DFF_LOW</type>
<position>49,-2244.5</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4826 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7044</ID>
<type>AE_DFF_LOW</type>
<position>97,-2442</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>5004 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7045</ID>
<type>BA_TRI_STATE</type>
<position>107,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5004 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7046</ID>
<type>AE_DFF_LOW</type>
<position>120,-2442</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>5005 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7047</ID>
<type>BA_TRI_STATE</type>
<position>130,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5005 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7048</ID>
<type>AE_DFF_LOW</type>
<position>143,-2442</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>5006 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7049</ID>
<type>BA_TRI_STATE</type>
<position>59,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4826 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7050</ID>
<type>BA_TRI_STATE</type>
<position>153,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5006 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7051</ID>
<type>AE_DFF_LOW</type>
<position>166,-2442</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>5007 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7052</ID>
<type>BA_TRI_STATE</type>
<position>176,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5007 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7053</ID>
<type>AE_DFF_LOW</type>
<position>191,-2442</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>5008 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7054</ID>
<type>BA_TRI_STATE</type>
<position>201,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5008 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7055</ID>
<type>AE_DFF_LOW</type>
<position>214,-2442</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>5009 </output>
<input>
<ID>clock</ID>5010 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7056</ID>
<type>BA_TRI_STATE</type>
<position>224,-2452.5</position>
<input>
<ID>ENABLE_0</ID>5011 </input>
<input>
<ID>IN_0</ID>5009 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7057</ID>
<type>HA_JUNC_2</type>
<position>40.5,-2355.5</position>
<input>
<ID>N_in0</ID>5012 </input>
<input>
<ID>N_in1</ID>5040 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7058</ID>
<type>HA_JUNC_2</type>
<position>63.5,-2355</position>
<input>
<ID>N_in0</ID>5013 </input>
<input>
<ID>N_in1</ID>5041 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7059</ID>
<type>HA_JUNC_2</type>
<position>66.5,-2355.5</position>
<input>
<ID>N_in0</ID>5014 </input>
<input>
<ID>N_in1</ID>5042 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7060</ID>
<type>HA_JUNC_2</type>
<position>86,-2355</position>
<input>
<ID>N_in0</ID>5015 </input>
<input>
<ID>N_in1</ID>5043 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7061</ID>
<type>HA_JUNC_2</type>
<position>89.5,-2355</position>
<input>
<ID>N_in0</ID>5016 </input>
<input>
<ID>N_in1</ID>5044 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7062</ID>
<type>HA_JUNC_2</type>
<position>110.5,-2355.5</position>
<input>
<ID>N_in0</ID>5017 </input>
<input>
<ID>N_in1</ID>5045 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7063</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2355</position>
<input>
<ID>N_in0</ID>5018 </input>
<input>
<ID>N_in1</ID>5046 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7064</ID>
<type>HA_JUNC_2</type>
<position>133,-2355</position>
<input>
<ID>N_in0</ID>5019 </input>
<input>
<ID>N_in1</ID>5047 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7065</ID>
<type>AE_DFF_LOW</type>
<position>72,-2244.5</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4827 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7066</ID>
<type>HA_JUNC_2</type>
<position>137,-2355</position>
<input>
<ID>N_in0</ID>5020 </input>
<input>
<ID>N_in1</ID>5048 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7067</ID>
<type>BA_TRI_STATE</type>
<position>82,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4827 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7068</ID>
<type>HA_JUNC_2</type>
<position>156,-2355</position>
<input>
<ID>N_in0</ID>5021 </input>
<input>
<ID>N_in1</ID>5049 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7069</ID>
<type>AE_DFF_LOW</type>
<position>97,-2244.5</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4828 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7070</ID>
<type>HA_JUNC_2</type>
<position>161,-2355</position>
<input>
<ID>N_in0</ID>5022 </input>
<input>
<ID>N_in1</ID>5050 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7071</ID>
<type>BA_TRI_STATE</type>
<position>107,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4828 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7072</ID>
<type>HA_JUNC_2</type>
<position>183.5,-2355</position>
<input>
<ID>N_in0</ID>5024 </input>
<input>
<ID>N_in1</ID>5052 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7073</ID>
<type>AE_DFF_LOW</type>
<position>120,-2244.5</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4829 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7074</ID>
<type>HA_JUNC_2</type>
<position>179,-2355</position>
<input>
<ID>N_in0</ID>5023 </input>
<input>
<ID>N_in1</ID>5051 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7075</ID>
<type>BA_TRI_STATE</type>
<position>130,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4829 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7076</ID>
<type>HA_JUNC_2</type>
<position>204.5,-2355.5</position>
<input>
<ID>N_in0</ID>5025 </input>
<input>
<ID>N_in1</ID>5053 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7077</ID>
<type>AE_DFF_LOW</type>
<position>143,-2244.5</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4830 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7078</ID>
<type>HA_JUNC_2</type>
<position>229,-2356.5</position>
<input>
<ID>N_in0</ID>5027 </input>
<input>
<ID>N_in1</ID>5055 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7079</ID>
<type>BA_TRI_STATE</type>
<position>153,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4830 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7080</ID>
<type>AA_AND2</type>
<position>21.5,-2421</position>
<input>
<ID>IN_0</ID>5031 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>4940 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7081</ID>
<type>AE_DFF_LOW</type>
<position>166,-2244.5</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4831 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7082</ID>
<type>AA_AND2</type>
<position>33,-2430.5</position>
<input>
<ID>IN_0</ID>5031 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>4941 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7083</ID>
<type>BA_TRI_STATE</type>
<position>176,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4831 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7084</ID>
<type>HA_JUNC_2</type>
<position>40.5,-2522.5</position>
<input>
<ID>N_in1</ID>5012 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7085</ID>
<type>AE_DFF_LOW</type>
<position>191,-2244.5</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4832 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7086</ID>
<type>AE_DFF_LOW</type>
<position>49,-2420</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4932 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7087</ID>
<type>BA_TRI_STATE</type>
<position>201,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4832 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7088</ID>
<type>HA_JUNC_2</type>
<position>63.5,-2522</position>
<input>
<ID>N_in1</ID>5013 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7089</ID>
<type>AE_DFF_LOW</type>
<position>214,-2244.5</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4833 </output>
<input>
<ID>clock</ID>4834 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7090</ID>
<type>HA_JUNC_2</type>
<position>66.5,-2522</position>
<input>
<ID>N_in1</ID>5014 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7091</ID>
<type>BA_TRI_STATE</type>
<position>224,-2255</position>
<input>
<ID>ENABLE_0</ID>4835 </input>
<input>
<ID>IN_0</ID>4833 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7092</ID>
<type>HA_JUNC_2</type>
<position>86,-2522</position>
<input>
<ID>N_in1</ID>5015 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7093</ID>
<type>AA_AND2</type>
<position>21.5,-2227</position>
<input>
<ID>IN_0</ID>4924 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4844 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7094</ID>
<type>HA_JUNC_2</type>
<position>89.5,-2522</position>
<input>
<ID>N_in1</ID>5016 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7095</ID>
<type>AA_AND2</type>
<position>33,-2236.5</position>
<input>
<ID>IN_0</ID>4924 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4845 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7096</ID>
<type>HA_JUNC_2</type>
<position>110.5,-2522</position>
<input>
<ID>N_in1</ID>5017 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7097</ID>
<type>AE_DFF_LOW</type>
<position>49,-2226</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4836 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7098</ID>
<type>BA_TRI_STATE</type>
<position>59,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4932 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7099</ID>
<type>BA_TRI_STATE</type>
<position>59,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4836 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7100</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2522</position>
<input>
<ID>N_in1</ID>5018 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7101</ID>
<type>AE_DFF_LOW</type>
<position>72,-2226</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4837 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7102</ID>
<type>HA_JUNC_2</type>
<position>133,-2522</position>
<input>
<ID>N_in1</ID>5019 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7103</ID>
<type>BA_TRI_STATE</type>
<position>82,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4837 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7104</ID>
<type>HA_JUNC_2</type>
<position>137,-2522</position>
<input>
<ID>N_in1</ID>5020 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7105</ID>
<type>AE_DFF_LOW</type>
<position>97,-2226</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4838 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7106</ID>
<type>HA_JUNC_2</type>
<position>156,-2521.5</position>
<input>
<ID>N_in1</ID>5021 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7107</ID>
<type>BA_TRI_STATE</type>
<position>107,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4838 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7108</ID>
<type>HA_JUNC_2</type>
<position>161,-2521.5</position>
<input>
<ID>N_in1</ID>5022 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7109</ID>
<type>AE_DFF_LOW</type>
<position>120,-2226</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4839 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7110</ID>
<type>HA_JUNC_2</type>
<position>179,-2521</position>
<input>
<ID>N_in1</ID>5023 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7111</ID>
<type>BA_TRI_STATE</type>
<position>130,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4839 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7112</ID>
<type>HA_JUNC_2</type>
<position>183.5,-2521</position>
<input>
<ID>N_in1</ID>5024 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7113</ID>
<type>AE_DFF_LOW</type>
<position>143,-2226</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4840 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7114</ID>
<type>HA_JUNC_2</type>
<position>204.5,-2520.5</position>
<input>
<ID>N_in1</ID>5025 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7115</ID>
<type>BA_TRI_STATE</type>
<position>153,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4840 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7116</ID>
<type>HA_JUNC_2</type>
<position>208,-2520.5</position>
<input>
<ID>N_in1</ID>5026 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7117</ID>
<type>AE_DFF_LOW</type>
<position>166,-2226</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4841 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7118</ID>
<type>HA_JUNC_2</type>
<position>208,-2355.5</position>
<input>
<ID>N_in0</ID>5026 </input>
<input>
<ID>N_in1</ID>5054 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7119</ID>
<type>BA_TRI_STATE</type>
<position>176,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4841 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7120</ID>
<type>HA_JUNC_2</type>
<position>229,-2520.5</position>
<input>
<ID>N_in1</ID>5027 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7121</ID>
<type>AE_DFF_LOW</type>
<position>191,-2226</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4842 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7122</ID>
<type>AE_DFF_LOW</type>
<position>72,-2420</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4933 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7123</ID>
<type>BA_TRI_STATE</type>
<position>201,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4842 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7124</ID>
<type>BA_TRI_STATE</type>
<position>82,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4933 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7125</ID>
<type>AE_DFF_LOW</type>
<position>214,-2226</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4843 </output>
<input>
<ID>clock</ID>4844 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7126</ID>
<type>HA_JUNC_2</type>
<position>27.5,-2355.5</position>
<input>
<ID>N_in0</ID>5037 </input>
<input>
<ID>N_in1</ID>5039 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7127</ID>
<type>BA_TRI_STATE</type>
<position>224,-2236.5</position>
<input>
<ID>ENABLE_0</ID>4845 </input>
<input>
<ID>IN_0</ID>4843 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7128</ID>
<type>AE_DFF_LOW</type>
<position>97,-2420</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4934 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7129</ID>
<type>AA_AND2</type>
<position>21.5,-2208</position>
<input>
<ID>IN_0</ID>4923 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4854 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7130</ID>
<type>HA_JUNC_2</type>
<position>17.5,-2355.5</position>
<input>
<ID>N_in0</ID>5036 </input>
<input>
<ID>N_in1</ID>5038 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7131</ID>
<type>AA_AND2</type>
<position>33,-2217.5</position>
<input>
<ID>IN_0</ID>4923 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4855 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7132</ID>
<type>BA_TRI_STATE</type>
<position>107,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4934 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7133</ID>
<type>AE_DFF_LOW</type>
<position>49,-2207</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4846 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7134</ID>
<type>HA_JUNC_2</type>
<position>27.5,-2522.5</position>
<input>
<ID>N_in1</ID>5037 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7135</ID>
<type>BA_TRI_STATE</type>
<position>59,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4846 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7136</ID>
<type>AE_DFF_LOW</type>
<position>120,-2420</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4935 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7137</ID>
<type>AE_DFF_LOW</type>
<position>72,-2207</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4847 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7138</ID>
<type>HA_JUNC_2</type>
<position>17.5,-2522.5</position>
<input>
<ID>N_in1</ID>5036 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7139</ID>
<type>BA_TRI_STATE</type>
<position>82,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4847 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7140</ID>
<type>BA_TRI_STATE</type>
<position>130,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4935 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7141</ID>
<type>AE_DFF_LOW</type>
<position>97,-2207</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4848 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7142</ID>
<type>AE_DFF_LOW</type>
<position>143,-2420</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4936 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7143</ID>
<type>BA_TRI_STATE</type>
<position>107,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4848 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7144</ID>
<type>AA_LABEL</type>
<position>8.5,-2356</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7145</ID>
<type>AE_DFF_LOW</type>
<position>120,-2207</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4849 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7146</ID>
<type>BA_TRI_STATE</type>
<position>153,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4936 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7147</ID>
<type>BA_TRI_STATE</type>
<position>130,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4849 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7148</ID>
<type>AE_DFF_LOW</type>
<position>166,-2420</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4937 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7149</ID>
<type>AE_DFF_LOW</type>
<position>143,-2207</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4850 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7150</ID>
<type>BA_TRI_STATE</type>
<position>176,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4937 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7151</ID>
<type>BA_TRI_STATE</type>
<position>153,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4850 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7152</ID>
<type>AE_DFF_LOW</type>
<position>191,-2420</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4938 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7153</ID>
<type>AE_DFF_LOW</type>
<position>166,-2207</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4851 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7154</ID>
<type>BA_TRI_STATE</type>
<position>201,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4938 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7155</ID>
<type>BA_TRI_STATE</type>
<position>176,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4851 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7156</ID>
<type>AE_DFF_LOW</type>
<position>214,-2420</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4939 </output>
<input>
<ID>clock</ID>4940 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7157</ID>
<type>AE_DFF_LOW</type>
<position>191,-2207</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4852 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7158</ID>
<type>BA_TRI_STATE</type>
<position>224,-2430.5</position>
<input>
<ID>ENABLE_0</ID>4941 </input>
<input>
<ID>IN_0</ID>4939 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7159</ID>
<type>BA_TRI_STATE</type>
<position>201,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4852 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7160</ID>
<type>AA_AND2</type>
<position>21.5,-2402.5</position>
<input>
<ID>IN_0</ID>5030 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>4950 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7161</ID>
<type>AE_DFF_LOW</type>
<position>214,-2207</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4853 </output>
<input>
<ID>clock</ID>4854 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7162</ID>
<type>AA_AND2</type>
<position>33,-2412</position>
<input>
<ID>IN_0</ID>5030 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>4951 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7163</ID>
<type>BA_TRI_STATE</type>
<position>224,-2217.5</position>
<input>
<ID>ENABLE_0</ID>4855 </input>
<input>
<ID>IN_0</ID>4853 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7164</ID>
<type>AE_DFF_LOW</type>
<position>49,-2401.5</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4942 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7165</ID>
<type>AA_AND2</type>
<position>21.5,-2189.5</position>
<input>
<ID>IN_0</ID>4922 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4864 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7166</ID>
<type>BA_TRI_STATE</type>
<position>59,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4942 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7167</ID>
<type>AA_AND2</type>
<position>33,-2199</position>
<input>
<ID>IN_0</ID>4922 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4865 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7168</ID>
<type>AE_DFF_LOW</type>
<position>72,-2401.5</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4943 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7169</ID>
<type>AE_DFF_LOW</type>
<position>49,-2188.5</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4856 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7170</ID>
<type>BA_TRI_STATE</type>
<position>82,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4943 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7171</ID>
<type>BA_TRI_STATE</type>
<position>59,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4856 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7172</ID>
<type>AE_DFF_LOW</type>
<position>97,-2401.5</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4944 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7173</ID>
<type>AE_DFF_LOW</type>
<position>72,-2188.5</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4857 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7174</ID>
<type>BA_TRI_STATE</type>
<position>107,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4944 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7175</ID>
<type>BA_TRI_STATE</type>
<position>82,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4857 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7176</ID>
<type>AE_DFF_LOW</type>
<position>120,-2401.5</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4945 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7177</ID>
<type>AE_DFF_LOW</type>
<position>97,-2188.5</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4858 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7178</ID>
<type>BA_TRI_STATE</type>
<position>130,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4945 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7179</ID>
<type>BA_TRI_STATE</type>
<position>107,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4858 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7180</ID>
<type>AE_DFF_LOW</type>
<position>143,-2401.5</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4946 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7181</ID>
<type>AE_DFF_LOW</type>
<position>120,-2188.5</position>
<input>
<ID>IN_0</ID>4912 </input>
<output>
<ID>OUT_0</ID>4859 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7182</ID>
<type>BA_TRI_STATE</type>
<position>153,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4946 </input>
<output>
<ID>OUT_0</ID>5021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7183</ID>
<type>BA_TRI_STATE</type>
<position>130,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4859 </input>
<output>
<ID>OUT_0</ID>4913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7184</ID>
<type>AE_DFF_LOW</type>
<position>166,-2401.5</position>
<input>
<ID>IN_0</ID>5022 </input>
<output>
<ID>OUT_0</ID>4947 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7185</ID>
<type>AE_DFF_LOW</type>
<position>143,-2188.5</position>
<input>
<ID>IN_0</ID>4914 </input>
<output>
<ID>OUT_0</ID>4860 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7186</ID>
<type>BA_TRI_STATE</type>
<position>176,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4947 </input>
<output>
<ID>OUT_0</ID>5023 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7187</ID>
<type>BA_TRI_STATE</type>
<position>153,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4860 </input>
<output>
<ID>OUT_0</ID>4915 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7188</ID>
<type>AE_DFF_LOW</type>
<position>191,-2401.5</position>
<input>
<ID>IN_0</ID>5024 </input>
<output>
<ID>OUT_0</ID>4948 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7189</ID>
<type>AE_DFF_LOW</type>
<position>166,-2188.5</position>
<input>
<ID>IN_0</ID>4916 </input>
<output>
<ID>OUT_0</ID>4861 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7190</ID>
<type>BA_TRI_STATE</type>
<position>201,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4948 </input>
<output>
<ID>OUT_0</ID>5025 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7191</ID>
<type>BA_TRI_STATE</type>
<position>176,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4861 </input>
<output>
<ID>OUT_0</ID>4917 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7192</ID>
<type>AE_DFF_LOW</type>
<position>214,-2401.5</position>
<input>
<ID>IN_0</ID>5026 </input>
<output>
<ID>OUT_0</ID>4949 </output>
<input>
<ID>clock</ID>4950 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7193</ID>
<type>AE_DFF_LOW</type>
<position>191,-2188.5</position>
<input>
<ID>IN_0</ID>4918 </input>
<output>
<ID>OUT_0</ID>4862 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7194</ID>
<type>BA_TRI_STATE</type>
<position>224,-2412</position>
<input>
<ID>ENABLE_0</ID>4951 </input>
<input>
<ID>IN_0</ID>4949 </input>
<output>
<ID>OUT_0</ID>5027 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7195</ID>
<type>BA_TRI_STATE</type>
<position>201,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4862 </input>
<output>
<ID>OUT_0</ID>4919 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7196</ID>
<type>AA_AND2</type>
<position>21.5,-2383.5</position>
<input>
<ID>IN_0</ID>5029 </input>
<input>
<ID>IN_1</ID>5036 </input>
<output>
<ID>OUT</ID>4960 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7197</ID>
<type>AE_DFF_LOW</type>
<position>214,-2188.5</position>
<input>
<ID>IN_0</ID>4920 </input>
<output>
<ID>OUT_0</ID>4863 </output>
<input>
<ID>clock</ID>4864 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7198</ID>
<type>AA_AND2</type>
<position>33,-2393</position>
<input>
<ID>IN_0</ID>5029 </input>
<input>
<ID>IN_1</ID>5037 </input>
<output>
<ID>OUT</ID>4961 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7199</ID>
<type>BA_TRI_STATE</type>
<position>224,-2199</position>
<input>
<ID>ENABLE_0</ID>4865 </input>
<input>
<ID>IN_0</ID>4863 </input>
<output>
<ID>OUT_0</ID>4921 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7200</ID>
<type>AE_DFF_LOW</type>
<position>49,-2382.5</position>
<input>
<ID>IN_0</ID>5012 </input>
<output>
<ID>OUT_0</ID>4952 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7201</ID>
<type>AA_AND2</type>
<position>21.5,-2323.5</position>
<input>
<ID>IN_0</ID>4929 </input>
<input>
<ID>IN_1</ID>4930 </input>
<output>
<ID>OUT</ID>4874 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7202</ID>
<type>BA_TRI_STATE</type>
<position>59,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4952 </input>
<output>
<ID>OUT_0</ID>5013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7203</ID>
<type>AA_AND2</type>
<position>32.5,-2333</position>
<input>
<ID>IN_0</ID>4929 </input>
<input>
<ID>IN_1</ID>4931 </input>
<output>
<ID>OUT</ID>4875 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7204</ID>
<type>AE_DFF_LOW</type>
<position>72,-2382.5</position>
<input>
<ID>IN_0</ID>5014 </input>
<output>
<ID>OUT_0</ID>4953 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7205</ID>
<type>AE_DFF_LOW</type>
<position>49,-2322.5</position>
<input>
<ID>IN_0</ID>4906 </input>
<output>
<ID>OUT_0</ID>4866 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7206</ID>
<type>BA_TRI_STATE</type>
<position>82,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4953 </input>
<output>
<ID>OUT_0</ID>5015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7207</ID>
<type>BA_TRI_STATE</type>
<position>59,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4866 </input>
<output>
<ID>OUT_0</ID>4907 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7208</ID>
<type>AE_DFF_LOW</type>
<position>97,-2382.5</position>
<input>
<ID>IN_0</ID>5016 </input>
<output>
<ID>OUT_0</ID>4954 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7209</ID>
<type>AE_DFF_LOW</type>
<position>72,-2322.5</position>
<input>
<ID>IN_0</ID>4908 </input>
<output>
<ID>OUT_0</ID>4867 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7210</ID>
<type>BA_TRI_STATE</type>
<position>107,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4954 </input>
<output>
<ID>OUT_0</ID>5017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7211</ID>
<type>BA_TRI_STATE</type>
<position>82,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4867 </input>
<output>
<ID>OUT_0</ID>4909 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7212</ID>
<type>AE_DFF_LOW</type>
<position>120,-2382.5</position>
<input>
<ID>IN_0</ID>5018 </input>
<output>
<ID>OUT_0</ID>4955 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7213</ID>
<type>AE_DFF_LOW</type>
<position>97,-2322.5</position>
<input>
<ID>IN_0</ID>4910 </input>
<output>
<ID>OUT_0</ID>4868 </output>
<input>
<ID>clock</ID>4874 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7214</ID>
<type>BA_TRI_STATE</type>
<position>130,-2393</position>
<input>
<ID>ENABLE_0</ID>4961 </input>
<input>
<ID>IN_0</ID>4955 </input>
<output>
<ID>OUT_0</ID>5019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7215</ID>
<type>BA_TRI_STATE</type>
<position>107,-2333</position>
<input>
<ID>ENABLE_0</ID>4875 </input>
<input>
<ID>IN_0</ID>4868 </input>
<output>
<ID>OUT_0</ID>4911 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7216</ID>
<type>AE_DFF_LOW</type>
<position>143,-2382.5</position>
<input>
<ID>IN_0</ID>5020 </input>
<output>
<ID>OUT_0</ID>4956 </output>
<input>
<ID>clock</ID>4960 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7218</ID>
<type>AA_LABEL</type>
<position>263,-2348.5</position>
<gparam>LABEL_TEXT 7</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7219</ID>
<type>AE_DFF_LOW</type>
<position>124,-2712.5</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5099 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7220</ID>
<type>BA_TRI_STATE</type>
<position>157,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5186 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7221</ID>
<type>BA_TRI_STATE</type>
<position>134,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5099 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7222</ID>
<type>AE_DFF_LOW</type>
<position>170,-2772.5</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5187 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7223</ID>
<type>AE_DFF_LOW</type>
<position>147,-2712.5</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5100 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7224</ID>
<type>BA_TRI_STATE</type>
<position>180,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5187 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7225</ID>
<type>BA_TRI_STATE</type>
<position>157,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5100 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7226</ID>
<type>AE_DFF_LOW</type>
<position>195,-2772.5</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5188 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7227</ID>
<type>AE_DFF_LOW</type>
<position>170,-2712.5</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5101 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7228</ID>
<type>BA_TRI_STATE</type>
<position>205,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5188 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7229</ID>
<type>BA_TRI_STATE</type>
<position>180,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5101 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7230</ID>
<type>AE_DFF_LOW</type>
<position>218,-2772.5</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5189 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7231</ID>
<type>AE_DFF_LOW</type>
<position>195,-2712.5</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5102 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7232</ID>
<type>BA_TRI_STATE</type>
<position>228,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5189 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7233</ID>
<type>BA_TRI_STATE</type>
<position>205,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5102 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7234</ID>
<type>AA_AND2</type>
<position>25.5,-2755</position>
<input>
<ID>IN_0</ID>5258 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7235</ID>
<type>AE_DFF_LOW</type>
<position>218,-2712.5</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5103 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7236</ID>
<type>AA_AND2</type>
<position>37,-2764.5</position>
<input>
<ID>IN_0</ID>5258 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7237</ID>
<type>BA_TRI_STATE</type>
<position>228,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5103 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7238</ID>
<type>AE_DFF_LOW</type>
<position>53,-2754</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5192 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7239</ID>
<type>AA_AND2</type>
<position>25.5,-2695</position>
<input>
<ID>IN_0</ID>5158 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7240</ID>
<type>BA_TRI_STATE</type>
<position>63,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5192 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7241</ID>
<type>AA_AND2</type>
<position>36.5,-2704.5</position>
<input>
<ID>IN_0</ID>5158 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7242</ID>
<type>AE_DFF_LOW</type>
<position>76,-2754</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5193 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7243</ID>
<type>AE_DFF_LOW</type>
<position>53,-2694</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5106 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7244</ID>
<type>BA_TRI_STATE</type>
<position>86,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5193 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7245</ID>
<type>BA_TRI_STATE</type>
<position>63,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5106 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7246</ID>
<type>AE_DFF_LOW</type>
<position>101,-2754</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5194 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7247</ID>
<type>AE_DFF_LOW</type>
<position>76,-2694</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5107 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7248</ID>
<type>BA_TRI_STATE</type>
<position>111,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5194 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7249</ID>
<type>BA_TRI_STATE</type>
<position>86,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5107 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7250</ID>
<type>AE_DFF_LOW</type>
<position>124,-2754</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5195 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7251</ID>
<type>AE_DFF_LOW</type>
<position>101,-2694</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5108 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7252</ID>
<type>BA_TRI_STATE</type>
<position>134,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5195 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7253</ID>
<type>BA_TRI_STATE</type>
<position>111,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5108 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7254</ID>
<type>AE_DFF_LOW</type>
<position>147,-2754</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5196 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7255</ID>
<type>AE_DFF_LOW</type>
<position>124,-2694</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5109 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7256</ID>
<type>BA_TRI_STATE</type>
<position>157,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5196 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7257</ID>
<type>BA_TRI_STATE</type>
<position>134,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5109 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7258</ID>
<type>AE_DFF_LOW</type>
<position>170,-2754</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5197 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7259</ID>
<type>AE_DFF_LOW</type>
<position>147,-2694</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5110 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7260</ID>
<type>BA_TRI_STATE</type>
<position>180,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5197 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7261</ID>
<type>BA_TRI_STATE</type>
<position>157,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5110 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7262</ID>
<type>AE_DFF_LOW</type>
<position>195,-2754</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5198 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7263</ID>
<type>AE_DFF_LOW</type>
<position>170,-2694</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5111 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7264</ID>
<type>BA_TRI_STATE</type>
<position>205,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5198 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7265</ID>
<type>BA_TRI_STATE</type>
<position>180,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5111 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7266</ID>
<type>AE_DFF_LOW</type>
<position>218,-2754</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5199 </output>
<input>
<ID>clock</ID>5200 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7267</ID>
<type>AE_DFF_LOW</type>
<position>195,-2694</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5112 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7268</ID>
<type>BA_TRI_STATE</type>
<position>228,-2764.5</position>
<input>
<ID>ENABLE_0</ID>5201 </input>
<input>
<ID>IN_0</ID>5199 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7269</ID>
<type>BA_TRI_STATE</type>
<position>205,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5112 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7270</ID>
<type>AA_AND2</type>
<position>25.5,-2889</position>
<input>
<ID>IN_0</ID>5265 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7271</ID>
<type>AE_DFF_LOW</type>
<position>218,-2694</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5113 </output>
<input>
<ID>clock</ID>5114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7272</ID>
<type>AA_AND2</type>
<position>36.5,-2898.5</position>
<input>
<ID>IN_0</ID>5265 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7273</ID>
<type>BA_TRI_STATE</type>
<position>228,-2704.5</position>
<input>
<ID>ENABLE_0</ID>5115 </input>
<input>
<ID>IN_0</ID>5113 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7274</ID>
<type>AE_DFF_LOW</type>
<position>53,-2888</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5202 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7275</ID>
<type>AA_AND2</type>
<position>36.5,-2861</position>
<input>
<ID>IN_0</ID>5263 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7276</ID>
<type>AA_AND2</type>
<position>25.5,-2676</position>
<input>
<ID>IN_0</ID>5157 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7277</ID>
<type>BA_TRI_STATE</type>
<position>63,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5202 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7278</ID>
<type>AA_AND2</type>
<position>36.5,-2685.5</position>
<input>
<ID>IN_0</ID>5157 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7279</ID>
<type>AE_DFF_LOW</type>
<position>76,-2888</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5203 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7280</ID>
<type>AE_DFF_LOW</type>
<position>53,-2850.5</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5222 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7281</ID>
<type>AE_DFF_LOW</type>
<position>53,-2675</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5116 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7282</ID>
<type>BA_TRI_STATE</type>
<position>86,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5203 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7283</ID>
<type>BA_TRI_STATE</type>
<position>63,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5116 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7284</ID>
<type>AE_DFF_LOW</type>
<position>101,-2888</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5204 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7285</ID>
<type>BA_TRI_STATE</type>
<position>63,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5222 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7286</ID>
<type>AE_DFF_LOW</type>
<position>76,-2675</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5117 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7287</ID>
<type>BA_TRI_STATE</type>
<position>111,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5204 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7288</ID>
<type>BA_TRI_STATE</type>
<position>86,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5117 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7289</ID>
<type>AE_DFF_LOW</type>
<position>124,-2888</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5205 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7290</ID>
<type>AE_DFF_LOW</type>
<position>76,-2850.5</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5223 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7291</ID>
<type>AE_DFF_LOW</type>
<position>101,-2675</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5118 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7292</ID>
<type>BA_TRI_STATE</type>
<position>134,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5205 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7293</ID>
<type>BA_TRI_STATE</type>
<position>111,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5118 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7294</ID>
<type>AE_DFF_LOW</type>
<position>147,-2888</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5206 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7295</ID>
<type>BA_TRI_STATE</type>
<position>86,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5223 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7296</ID>
<type>AE_DFF_LOW</type>
<position>124,-2675</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5119 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7297</ID>
<type>BA_TRI_STATE</type>
<position>157,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5206 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7298</ID>
<type>BA_TRI_STATE</type>
<position>134,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5119 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7299</ID>
<type>AE_DFF_LOW</type>
<position>170,-2888</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5207 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7300</ID>
<type>AE_DFF_LOW</type>
<position>101,-2850.5</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5224 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7301</ID>
<type>AE_DFF_LOW</type>
<position>147,-2675</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5120 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7302</ID>
<type>BA_TRI_STATE</type>
<position>180,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5207 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7303</ID>
<type>BA_TRI_STATE</type>
<position>157,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5120 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7304</ID>
<type>BA_TRI_STATE</type>
<position>111,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5224 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7305</ID>
<type>AE_DFF_LOW</type>
<position>170,-2675</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5121 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7306</ID>
<type>BA_TRI_STATE</type>
<position>180,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5121 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7307</ID>
<type>AE_DFF_LOW</type>
<position>124,-2850.5</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5225 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7308</ID>
<type>AE_DFF_LOW</type>
<position>195,-2675</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5122 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7309</ID>
<type>BA_TRI_STATE</type>
<position>205,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5122 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7310</ID>
<type>AE_DFF_LOW</type>
<position>218,-2675</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5123 </output>
<input>
<ID>clock</ID>5124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7311</ID>
<type>BA_TRI_STATE</type>
<position>228,-2685.5</position>
<input>
<ID>ENABLE_0</ID>5125 </input>
<input>
<ID>IN_0</ID>5123 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7312</ID>
<type>AA_AND2</type>
<position>25.5,-2657.5</position>
<input>
<ID>IN_0</ID>5156 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7313</ID>
<type>AA_AND2</type>
<position>36.5,-2667</position>
<input>
<ID>IN_0</ID>5156 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7314</ID>
<type>AE_DFF_LOW</type>
<position>53,-2656.5</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5126 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7315</ID>
<type>BA_TRI_STATE</type>
<position>63,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5126 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7316</ID>
<type>AE_DFF_LOW</type>
<position>76,-2656.5</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5127 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7317</ID>
<type>BA_TRI_STATE</type>
<position>86,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5127 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7318</ID>
<type>AE_DFF_LOW</type>
<position>101,-2656.5</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5128 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7319</ID>
<type>BA_TRI_STATE</type>
<position>111,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5128 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7320</ID>
<type>AE_DFF_LOW</type>
<position>124,-2656.5</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5129 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7321</ID>
<type>BA_TRI_STATE</type>
<position>134,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5129 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7322</ID>
<type>AE_DFF_LOW</type>
<position>147,-2656.5</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5130 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7323</ID>
<type>BA_TRI_STATE</type>
<position>157,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5130 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7324</ID>
<type>AE_DFF_LOW</type>
<position>170,-2656.5</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5131 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7325</ID>
<type>BA_TRI_STATE</type>
<position>180,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5131 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7326</ID>
<type>AE_DFF_LOW</type>
<position>195,-2656.5</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5132 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7327</ID>
<type>BA_TRI_STATE</type>
<position>205,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5132 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7328</ID>
<type>AE_DFF_LOW</type>
<position>218,-2656.5</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5133 </output>
<input>
<ID>clock</ID>5134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7329</ID>
<type>BA_TRI_STATE</type>
<position>228,-2667</position>
<input>
<ID>ENABLE_0</ID>5135 </input>
<input>
<ID>IN_0</ID>5133 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7330</ID>
<type>HA_JUNC_2</type>
<position>44.5,-2570</position>
<input>
<ID>N_in0</ID>5136 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7331</ID>
<type>HA_JUNC_2</type>
<position>67.5,-2569.5</position>
<input>
<ID>N_in0</ID>5137 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7332</ID>
<type>HA_JUNC_2</type>
<position>70.5,-2570</position>
<input>
<ID>N_in0</ID>5138 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7333</ID>
<type>HA_JUNC_2</type>
<position>90,-2569.5</position>
<input>
<ID>N_in0</ID>5139 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7334</ID>
<type>HA_JUNC_2</type>
<position>93.5,-2569.5</position>
<input>
<ID>N_in0</ID>5140 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7335</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2570</position>
<input>
<ID>N_in0</ID>5141 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7336</ID>
<type>HA_JUNC_2</type>
<position>118.5,-2569.5</position>
<input>
<ID>N_in0</ID>5142 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7337</ID>
<type>HA_JUNC_2</type>
<position>137,-2569.5</position>
<input>
<ID>N_in0</ID>5143 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7338</ID>
<type>HA_JUNC_2</type>
<position>141,-2569.5</position>
<input>
<ID>N_in0</ID>5144 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7339</ID>
<type>HA_JUNC_2</type>
<position>160,-2569.5</position>
<input>
<ID>N_in0</ID>5145 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7340</ID>
<type>HA_JUNC_2</type>
<position>165,-2569.5</position>
<input>
<ID>N_in0</ID>5146 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7341</ID>
<type>HA_JUNC_2</type>
<position>187.5,-2569.5</position>
<input>
<ID>N_in0</ID>5148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7342</ID>
<type>HA_JUNC_2</type>
<position>183,-2569.5</position>
<input>
<ID>N_in0</ID>5147 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7343</ID>
<type>HA_JUNC_2</type>
<position>208.5,-2570</position>
<input>
<ID>N_in0</ID>5149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7344</ID>
<type>HA_JUNC_2</type>
<position>233,-2571</position>
<input>
<ID>N_in0</ID>5151 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7345</ID>
<type>HA_JUNC_2</type>
<position>44.5,-2737</position>
<input>
<ID>N_in0</ID>5270 </input>
<input>
<ID>N_in1</ID>5136 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7346</ID>
<type>HA_JUNC_2</type>
<position>67.5,-2736.5</position>
<input>
<ID>N_in0</ID>5271 </input>
<input>
<ID>N_in1</ID>5137 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7347</ID>
<type>HA_JUNC_2</type>
<position>70.5,-2736.5</position>
<input>
<ID>N_in0</ID>5272 </input>
<input>
<ID>N_in1</ID>5138 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7348</ID>
<type>HA_JUNC_2</type>
<position>90,-2736.5</position>
<input>
<ID>N_in0</ID>5273 </input>
<input>
<ID>N_in1</ID>5139 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7349</ID>
<type>HA_JUNC_2</type>
<position>93.5,-2736.5</position>
<input>
<ID>N_in0</ID>5274 </input>
<input>
<ID>N_in1</ID>5140 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7350</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2736.5</position>
<input>
<ID>N_in0</ID>5275 </input>
<input>
<ID>N_in1</ID>5141 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7351</ID>
<type>HA_JUNC_2</type>
<position>118.5,-2736.5</position>
<input>
<ID>N_in0</ID>5276 </input>
<input>
<ID>N_in1</ID>5142 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7352</ID>
<type>HA_JUNC_2</type>
<position>137,-2736.5</position>
<input>
<ID>N_in0</ID>5277 </input>
<input>
<ID>N_in1</ID>5143 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7353</ID>
<type>HA_JUNC_2</type>
<position>141,-2736.5</position>
<input>
<ID>N_in0</ID>5278 </input>
<input>
<ID>N_in1</ID>5144 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7354</ID>
<type>HA_JUNC_2</type>
<position>160,-2736</position>
<input>
<ID>N_in0</ID>5279 </input>
<input>
<ID>N_in1</ID>5145 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7355</ID>
<type>HA_JUNC_2</type>
<position>165,-2736</position>
<input>
<ID>N_in0</ID>5280 </input>
<input>
<ID>N_in1</ID>5146 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7356</ID>
<type>HA_JUNC_2</type>
<position>183,-2735.5</position>
<input>
<ID>N_in0</ID>5281 </input>
<input>
<ID>N_in1</ID>5147 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7357</ID>
<type>HA_JUNC_2</type>
<position>187.5,-2735.5</position>
<input>
<ID>N_in0</ID>5282 </input>
<input>
<ID>N_in1</ID>5148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7358</ID>
<type>HA_JUNC_2</type>
<position>208.5,-2735</position>
<input>
<ID>N_in0</ID>5283 </input>
<input>
<ID>N_in1</ID>5149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7359</ID>
<type>HA_JUNC_2</type>
<position>212,-2735</position>
<input>
<ID>N_in0</ID>5284 </input>
<input>
<ID>N_in1</ID>5150 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7360</ID>
<type>HA_JUNC_2</type>
<position>212,-2570</position>
<input>
<ID>N_in0</ID>5150 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7361</ID>
<type>HA_JUNC_2</type>
<position>233,-2735</position>
<input>
<ID>N_in0</ID>5285 </input>
<input>
<ID>N_in1</ID>5151 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7362</ID>
<type>HA_JUNC_2</type>
<position>31.5,-2570</position>
<input>
<ID>N_in0</ID>5161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7363</ID>
<type>HA_JUNC_2</type>
<position>21.5,-2570</position>
<input>
<ID>N_in0</ID>5160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7364</ID>
<type>HA_JUNC_2</type>
<position>31.5,-2737</position>
<input>
<ID>N_in0</ID>5269 </input>
<input>
<ID>N_in1</ID>5161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7365</ID>
<type>HA_JUNC_2</type>
<position>21.5,-2737</position>
<input>
<ID>N_in0</ID>5268 </input>
<input>
<ID>N_in1</ID>5160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7366</ID>
<type>AA_LABEL</type>
<position>12.5,-2570.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7367</ID>
<type>BI_DECODER_4x16</type>
<position>-127,-2737.5</position>
<output>
<ID>OUT_0</ID>5265 </output>
<output>
<ID>OUT_1</ID>5264 </output>
<output>
<ID>OUT_10</ID>5157 </output>
<output>
<ID>OUT_11</ID>5156 </output>
<output>
<ID>OUT_12</ID>5155 </output>
<output>
<ID>OUT_13</ID>5154 </output>
<output>
<ID>OUT_14</ID>5153 </output>
<output>
<ID>OUT_15</ID>5152 </output>
<output>
<ID>OUT_2</ID>5263 </output>
<output>
<ID>OUT_3</ID>5262 </output>
<output>
<ID>OUT_4</ID>5261 </output>
<output>
<ID>OUT_5</ID>5260 </output>
<output>
<ID>OUT_6</ID>5259 </output>
<output>
<ID>OUT_7</ID>5258 </output>
<output>
<ID>OUT_8</ID>5159 </output>
<output>
<ID>OUT_9</ID>5158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7368</ID>
<type>AE_DFF_LOW</type>
<position>195,-2888</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5208 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7369</ID>
<type>BA_TRI_STATE</type>
<position>205,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5208 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7370</ID>
<type>AE_DFF_LOW</type>
<position>218,-2888</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5209 </output>
<input>
<ID>clock</ID>5210 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7371</ID>
<type>BA_TRI_STATE</type>
<position>228,-2898.5</position>
<input>
<ID>ENABLE_0</ID>5211 </input>
<input>
<ID>IN_0</ID>5209 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7372</ID>
<type>AA_AND2</type>
<position>25.5,-2870.5</position>
<input>
<ID>IN_0</ID>5264 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7373</ID>
<type>AA_AND2</type>
<position>36.5,-2880</position>
<input>
<ID>IN_0</ID>5264 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7374</ID>
<type>AE_DFF_LOW</type>
<position>53,-2869.5</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5212 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7375</ID>
<type>BA_TRI_STATE</type>
<position>63,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5212 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7376</ID>
<type>AE_DFF_LOW</type>
<position>76,-2869.5</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5213 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7377</ID>
<type>BA_TRI_STATE</type>
<position>86,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5213 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7378</ID>
<type>AE_DFF_LOW</type>
<position>101,-2869.5</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5214 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7379</ID>
<type>BA_TRI_STATE</type>
<position>111,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5214 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7380</ID>
<type>AE_DFF_LOW</type>
<position>124,-2869.5</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5215 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7381</ID>
<type>BA_TRI_STATE</type>
<position>134,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5215 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7382</ID>
<type>AE_DFF_LOW</type>
<position>147,-2869.5</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5216 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7383</ID>
<type>BA_TRI_STATE</type>
<position>157,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5216 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7384</ID>
<type>AE_DFF_LOW</type>
<position>170,-2869.5</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5217 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7385</ID>
<type>BA_TRI_STATE</type>
<position>180,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5217 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7386</ID>
<type>AE_DFF_LOW</type>
<position>195,-2869.5</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5218 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7387</ID>
<type>BA_TRI_STATE</type>
<position>205,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5218 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7388</ID>
<type>AE_DFF_LOW</type>
<position>218,-2869.5</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5219 </output>
<input>
<ID>clock</ID>5220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7389</ID>
<type>BA_TRI_STATE</type>
<position>228,-2880</position>
<input>
<ID>ENABLE_0</ID>5221 </input>
<input>
<ID>IN_0</ID>5219 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7390</ID>
<type>AA_AND2</type>
<position>25.5,-2851.5</position>
<input>
<ID>IN_0</ID>5263 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7391</ID>
<type>BA_TRI_STATE</type>
<position>134,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5225 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7392</ID>
<type>AE_DFF_LOW</type>
<position>147,-2850.5</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5226 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7393</ID>
<type>BA_TRI_STATE</type>
<position>157,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5226 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7394</ID>
<type>AE_DFF_LOW</type>
<position>170,-2850.5</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5227 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7395</ID>
<type>BA_TRI_STATE</type>
<position>180,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5227 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7396</ID>
<type>AE_DFF_LOW</type>
<position>195,-2850.5</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5228 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7397</ID>
<type>BA_TRI_STATE</type>
<position>205,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5228 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7398</ID>
<type>AA_AND2</type>
<position>25.5,-2635.5</position>
<input>
<ID>IN_0</ID>5155 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7399</ID>
<type>AE_DFF_LOW</type>
<position>218,-2850.5</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5229 </output>
<input>
<ID>clock</ID>5230 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7400</ID>
<type>BA_TRI_STATE</type>
<position>228,-2861</position>
<input>
<ID>ENABLE_0</ID>5231 </input>
<input>
<ID>IN_0</ID>5229 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7401</ID>
<type>AA_AND2</type>
<position>25.5,-2833</position>
<input>
<ID>IN_0</ID>5262 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7402</ID>
<type>AA_AND2</type>
<position>36.5,-2842.5</position>
<input>
<ID>IN_0</ID>5262 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7403</ID>
<type>AA_AND2</type>
<position>37,-2645</position>
<input>
<ID>IN_0</ID>5155 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5065 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7404</ID>
<type>AE_DFF_LOW</type>
<position>53,-2832</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5232 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7405</ID>
<type>BA_TRI_STATE</type>
<position>63,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5232 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7406</ID>
<type>AE_DFF_LOW</type>
<position>76,-2832</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5233 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7407</ID>
<type>BA_TRI_STATE</type>
<position>86,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5233 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7408</ID>
<type>AE_DFF_LOW</type>
<position>53,-2634.5</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5056 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7409</ID>
<type>AE_DFF_LOW</type>
<position>101,-2832</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5234 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7410</ID>
<type>BA_TRI_STATE</type>
<position>111,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5234 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7411</ID>
<type>AE_DFF_LOW</type>
<position>124,-2832</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5235 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7412</ID>
<type>BA_TRI_STATE</type>
<position>134,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5235 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7413</ID>
<type>AE_DFF_LOW</type>
<position>147,-2832</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5236 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7414</ID>
<type>BA_TRI_STATE</type>
<position>63,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5056 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7415</ID>
<type>BA_TRI_STATE</type>
<position>157,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5236 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7416</ID>
<type>AE_DFF_LOW</type>
<position>170,-2832</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5237 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7417</ID>
<type>BA_TRI_STATE</type>
<position>180,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5237 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7418</ID>
<type>AE_DFF_LOW</type>
<position>195,-2832</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5238 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7419</ID>
<type>BA_TRI_STATE</type>
<position>205,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5238 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7420</ID>
<type>AE_DFF_LOW</type>
<position>218,-2832</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5239 </output>
<input>
<ID>clock</ID>5240 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7421</ID>
<type>BA_TRI_STATE</type>
<position>228,-2842.5</position>
<input>
<ID>ENABLE_0</ID>5241 </input>
<input>
<ID>IN_0</ID>5239 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7422</ID>
<type>HA_JUNC_2</type>
<position>44.5,-2745.5</position>
<input>
<ID>N_in0</ID>5242 </input>
<input>
<ID>N_in1</ID>5270 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7423</ID>
<type>HA_JUNC_2</type>
<position>67.5,-2745</position>
<input>
<ID>N_in0</ID>5243 </input>
<input>
<ID>N_in1</ID>5271 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7424</ID>
<type>HA_JUNC_2</type>
<position>70.5,-2745.5</position>
<input>
<ID>N_in0</ID>5244 </input>
<input>
<ID>N_in1</ID>5272 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7425</ID>
<type>HA_JUNC_2</type>
<position>90,-2745</position>
<input>
<ID>N_in0</ID>5245 </input>
<input>
<ID>N_in1</ID>5273 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7426</ID>
<type>HA_JUNC_2</type>
<position>93.5,-2745</position>
<input>
<ID>N_in0</ID>5246 </input>
<input>
<ID>N_in1</ID>5274 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7427</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2745.5</position>
<input>
<ID>N_in0</ID>5247 </input>
<input>
<ID>N_in1</ID>5275 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7428</ID>
<type>HA_JUNC_2</type>
<position>118.5,-2745</position>
<input>
<ID>N_in0</ID>5248 </input>
<input>
<ID>N_in1</ID>5276 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7429</ID>
<type>HA_JUNC_2</type>
<position>137,-2745</position>
<input>
<ID>N_in0</ID>5249 </input>
<input>
<ID>N_in1</ID>5277 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7430</ID>
<type>AE_DFF_LOW</type>
<position>76,-2634.5</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5057 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7431</ID>
<type>HA_JUNC_2</type>
<position>141,-2745</position>
<input>
<ID>N_in0</ID>5250 </input>
<input>
<ID>N_in1</ID>5278 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7432</ID>
<type>BA_TRI_STATE</type>
<position>86,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5057 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7433</ID>
<type>HA_JUNC_2</type>
<position>160,-2745</position>
<input>
<ID>N_in0</ID>5251 </input>
<input>
<ID>N_in1</ID>5279 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7434</ID>
<type>AE_DFF_LOW</type>
<position>101,-2634.5</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5058 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7435</ID>
<type>HA_JUNC_2</type>
<position>165,-2745</position>
<input>
<ID>N_in0</ID>5252 </input>
<input>
<ID>N_in1</ID>5280 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7436</ID>
<type>BA_TRI_STATE</type>
<position>111,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5058 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7437</ID>
<type>HA_JUNC_2</type>
<position>187.5,-2745</position>
<input>
<ID>N_in0</ID>5254 </input>
<input>
<ID>N_in1</ID>5282 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7438</ID>
<type>AE_DFF_LOW</type>
<position>124,-2634.5</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5059 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7439</ID>
<type>HA_JUNC_2</type>
<position>183,-2745</position>
<input>
<ID>N_in0</ID>5253 </input>
<input>
<ID>N_in1</ID>5281 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7440</ID>
<type>BA_TRI_STATE</type>
<position>134,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5059 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7441</ID>
<type>HA_JUNC_2</type>
<position>208.5,-2745.5</position>
<input>
<ID>N_in0</ID>5255 </input>
<input>
<ID>N_in1</ID>5283 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7442</ID>
<type>AE_DFF_LOW</type>
<position>147,-2634.5</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5060 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7443</ID>
<type>HA_JUNC_2</type>
<position>233,-2746.5</position>
<input>
<ID>N_in0</ID>5257 </input>
<input>
<ID>N_in1</ID>5285 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7444</ID>
<type>BA_TRI_STATE</type>
<position>157,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5060 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7445</ID>
<type>AA_AND2</type>
<position>25.5,-2811</position>
<input>
<ID>IN_0</ID>5261 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7446</ID>
<type>AE_DFF_LOW</type>
<position>170,-2634.5</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5061 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7447</ID>
<type>AA_AND2</type>
<position>37,-2820.5</position>
<input>
<ID>IN_0</ID>5261 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7448</ID>
<type>BA_TRI_STATE</type>
<position>180,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5061 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7449</ID>
<type>HA_JUNC_2</type>
<position>44.5,-2912.5</position>
<input>
<ID>N_in1</ID>5242 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7450</ID>
<type>AE_DFF_LOW</type>
<position>195,-2634.5</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5062 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7451</ID>
<type>AE_DFF_LOW</type>
<position>53,-2810</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5162 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7452</ID>
<type>BA_TRI_STATE</type>
<position>205,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5062 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7453</ID>
<type>HA_JUNC_2</type>
<position>67.5,-2912</position>
<input>
<ID>N_in1</ID>5243 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7454</ID>
<type>AE_DFF_LOW</type>
<position>218,-2634.5</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5063 </output>
<input>
<ID>clock</ID>5064 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7455</ID>
<type>HA_JUNC_2</type>
<position>70.5,-2912</position>
<input>
<ID>N_in1</ID>5244 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7456</ID>
<type>BA_TRI_STATE</type>
<position>228,-2645</position>
<input>
<ID>ENABLE_0</ID>5065 </input>
<input>
<ID>IN_0</ID>5063 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7457</ID>
<type>HA_JUNC_2</type>
<position>90,-2912</position>
<input>
<ID>N_in1</ID>5245 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7458</ID>
<type>AA_AND2</type>
<position>25.5,-2617</position>
<input>
<ID>IN_0</ID>5154 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7459</ID>
<type>HA_JUNC_2</type>
<position>93.5,-2912</position>
<input>
<ID>N_in1</ID>5246 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7460</ID>
<type>AA_AND2</type>
<position>37,-2626.5</position>
<input>
<ID>IN_0</ID>5154 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7461</ID>
<type>HA_JUNC_2</type>
<position>114.5,-2912</position>
<input>
<ID>N_in1</ID>5247 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7462</ID>
<type>AE_DFF_LOW</type>
<position>53,-2616</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5066 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7463</ID>
<type>BA_TRI_STATE</type>
<position>63,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5162 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7464</ID>
<type>BA_TRI_STATE</type>
<position>63,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5066 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7465</ID>
<type>HA_JUNC_2</type>
<position>118.5,-2912</position>
<input>
<ID>N_in1</ID>5248 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7466</ID>
<type>AE_DFF_LOW</type>
<position>76,-2616</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5067 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7467</ID>
<type>HA_JUNC_2</type>
<position>137,-2912</position>
<input>
<ID>N_in1</ID>5249 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7468</ID>
<type>BA_TRI_STATE</type>
<position>86,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5067 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7469</ID>
<type>HA_JUNC_2</type>
<position>141,-2912</position>
<input>
<ID>N_in1</ID>5250 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7470</ID>
<type>AE_DFF_LOW</type>
<position>101,-2616</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5068 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7471</ID>
<type>HA_JUNC_2</type>
<position>160,-2911.5</position>
<input>
<ID>N_in1</ID>5251 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7472</ID>
<type>BA_TRI_STATE</type>
<position>111,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5068 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7473</ID>
<type>HA_JUNC_2</type>
<position>165,-2911.5</position>
<input>
<ID>N_in1</ID>5252 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7474</ID>
<type>AE_DFF_LOW</type>
<position>124,-2616</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5069 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7475</ID>
<type>HA_JUNC_2</type>
<position>183,-2911</position>
<input>
<ID>N_in1</ID>5253 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7476</ID>
<type>BA_TRI_STATE</type>
<position>134,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5069 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7477</ID>
<type>HA_JUNC_2</type>
<position>187.5,-2911</position>
<input>
<ID>N_in1</ID>5254 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7478</ID>
<type>AE_DFF_LOW</type>
<position>147,-2616</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5070 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7479</ID>
<type>HA_JUNC_2</type>
<position>208.5,-2910.5</position>
<input>
<ID>N_in1</ID>5255 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7480</ID>
<type>BA_TRI_STATE</type>
<position>157,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5070 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7481</ID>
<type>HA_JUNC_2</type>
<position>212,-2910.5</position>
<input>
<ID>N_in1</ID>5256 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7482</ID>
<type>AE_DFF_LOW</type>
<position>170,-2616</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5071 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7483</ID>
<type>HA_JUNC_2</type>
<position>212,-2745.5</position>
<input>
<ID>N_in0</ID>5256 </input>
<input>
<ID>N_in1</ID>5284 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7484</ID>
<type>BA_TRI_STATE</type>
<position>180,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5071 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7485</ID>
<type>HA_JUNC_2</type>
<position>233,-2910.5</position>
<input>
<ID>N_in1</ID>5257 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7486</ID>
<type>AE_DFF_LOW</type>
<position>195,-2616</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5072 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7487</ID>
<type>AE_DFF_LOW</type>
<position>76,-2810</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5163 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7488</ID>
<type>BA_TRI_STATE</type>
<position>205,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5072 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7489</ID>
<type>BA_TRI_STATE</type>
<position>86,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5163 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7490</ID>
<type>AE_DFF_LOW</type>
<position>218,-2616</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5073 </output>
<input>
<ID>clock</ID>5074 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7491</ID>
<type>HA_JUNC_2</type>
<position>31.5,-2745.5</position>
<input>
<ID>N_in0</ID>5267 </input>
<input>
<ID>N_in1</ID>5269 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7492</ID>
<type>BA_TRI_STATE</type>
<position>228,-2626.5</position>
<input>
<ID>ENABLE_0</ID>5075 </input>
<input>
<ID>IN_0</ID>5073 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7493</ID>
<type>AE_DFF_LOW</type>
<position>101,-2810</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5164 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7494</ID>
<type>AA_AND2</type>
<position>25.5,-2598</position>
<input>
<ID>IN_0</ID>5153 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5084 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7495</ID>
<type>HA_JUNC_2</type>
<position>21.5,-2745.5</position>
<input>
<ID>N_in0</ID>5266 </input>
<input>
<ID>N_in1</ID>5268 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7496</ID>
<type>AA_AND2</type>
<position>37,-2607.5</position>
<input>
<ID>IN_0</ID>5153 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5085 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7497</ID>
<type>BA_TRI_STATE</type>
<position>111,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5164 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7498</ID>
<type>AE_DFF_LOW</type>
<position>53,-2597</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5076 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7499</ID>
<type>HA_JUNC_2</type>
<position>31.5,-2912.5</position>
<input>
<ID>N_in1</ID>5267 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7500</ID>
<type>BA_TRI_STATE</type>
<position>63,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5076 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7501</ID>
<type>AE_DFF_LOW</type>
<position>124,-2810</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5165 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7502</ID>
<type>AE_DFF_LOW</type>
<position>76,-2597</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5077 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7503</ID>
<type>HA_JUNC_2</type>
<position>21.5,-2912.5</position>
<input>
<ID>N_in1</ID>5266 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7504</ID>
<type>BA_TRI_STATE</type>
<position>86,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5077 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7505</ID>
<type>BA_TRI_STATE</type>
<position>134,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5165 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7506</ID>
<type>AE_DFF_LOW</type>
<position>101,-2597</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5078 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7507</ID>
<type>AE_DFF_LOW</type>
<position>147,-2810</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5166 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7508</ID>
<type>BA_TRI_STATE</type>
<position>111,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5078 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7509</ID>
<type>AA_LABEL</type>
<position>12.5,-2746</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7510</ID>
<type>AE_DFF_LOW</type>
<position>124,-2597</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5079 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7511</ID>
<type>BA_TRI_STATE</type>
<position>157,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5166 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7512</ID>
<type>BA_TRI_STATE</type>
<position>134,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5079 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7513</ID>
<type>AE_DFF_LOW</type>
<position>170,-2810</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5167 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7514</ID>
<type>AE_DFF_LOW</type>
<position>147,-2597</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5080 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7515</ID>
<type>BA_TRI_STATE</type>
<position>180,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5167 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7516</ID>
<type>BA_TRI_STATE</type>
<position>157,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5080 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7517</ID>
<type>AE_DFF_LOW</type>
<position>195,-2810</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5168 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7518</ID>
<type>AE_DFF_LOW</type>
<position>170,-2597</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5081 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7519</ID>
<type>BA_TRI_STATE</type>
<position>205,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5168 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7520</ID>
<type>BA_TRI_STATE</type>
<position>180,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5081 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7521</ID>
<type>AE_DFF_LOW</type>
<position>218,-2810</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5169 </output>
<input>
<ID>clock</ID>5170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7522</ID>
<type>AE_DFF_LOW</type>
<position>195,-2597</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5082 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7523</ID>
<type>BA_TRI_STATE</type>
<position>228,-2820.5</position>
<input>
<ID>ENABLE_0</ID>5171 </input>
<input>
<ID>IN_0</ID>5169 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7524</ID>
<type>BA_TRI_STATE</type>
<position>205,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5082 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7525</ID>
<type>AA_AND2</type>
<position>25.5,-2792.5</position>
<input>
<ID>IN_0</ID>5260 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7526</ID>
<type>AE_DFF_LOW</type>
<position>218,-2597</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5083 </output>
<input>
<ID>clock</ID>5084 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7527</ID>
<type>AA_AND2</type>
<position>37,-2802</position>
<input>
<ID>IN_0</ID>5260 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7528</ID>
<type>BA_TRI_STATE</type>
<position>228,-2607.5</position>
<input>
<ID>ENABLE_0</ID>5085 </input>
<input>
<ID>IN_0</ID>5083 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7529</ID>
<type>AE_DFF_LOW</type>
<position>53,-2791.5</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5172 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7530</ID>
<type>AA_AND2</type>
<position>25.5,-2579.5</position>
<input>
<ID>IN_0</ID>5152 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5094 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7531</ID>
<type>BA_TRI_STATE</type>
<position>63,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5172 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7532</ID>
<type>AA_AND2</type>
<position>37,-2589</position>
<input>
<ID>IN_0</ID>5152 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5095 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7533</ID>
<type>AE_DFF_LOW</type>
<position>76,-2791.5</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5173 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7534</ID>
<type>AE_DFF_LOW</type>
<position>53,-2578.5</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5086 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7535</ID>
<type>BA_TRI_STATE</type>
<position>86,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5173 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7536</ID>
<type>BA_TRI_STATE</type>
<position>63,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5086 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7537</ID>
<type>AE_DFF_LOW</type>
<position>101,-2791.5</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5174 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7538</ID>
<type>AE_DFF_LOW</type>
<position>76,-2578.5</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5087 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7539</ID>
<type>BA_TRI_STATE</type>
<position>111,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5174 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7540</ID>
<type>BA_TRI_STATE</type>
<position>86,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5087 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7541</ID>
<type>AE_DFF_LOW</type>
<position>124,-2791.5</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5175 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7542</ID>
<type>AE_DFF_LOW</type>
<position>101,-2578.5</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5088 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7543</ID>
<type>BA_TRI_STATE</type>
<position>134,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5175 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7544</ID>
<type>BA_TRI_STATE</type>
<position>111,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5088 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7545</ID>
<type>AE_DFF_LOW</type>
<position>147,-2791.5</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5176 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7546</ID>
<type>AE_DFF_LOW</type>
<position>124,-2578.5</position>
<input>
<ID>IN_0</ID>5142 </input>
<output>
<ID>OUT_0</ID>5089 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7547</ID>
<type>BA_TRI_STATE</type>
<position>157,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5176 </input>
<output>
<ID>OUT_0</ID>5251 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7548</ID>
<type>BA_TRI_STATE</type>
<position>134,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5089 </input>
<output>
<ID>OUT_0</ID>5143 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7549</ID>
<type>AE_DFF_LOW</type>
<position>170,-2791.5</position>
<input>
<ID>IN_0</ID>5252 </input>
<output>
<ID>OUT_0</ID>5177 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7550</ID>
<type>AE_DFF_LOW</type>
<position>147,-2578.5</position>
<input>
<ID>IN_0</ID>5144 </input>
<output>
<ID>OUT_0</ID>5090 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7551</ID>
<type>BA_TRI_STATE</type>
<position>180,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5177 </input>
<output>
<ID>OUT_0</ID>5253 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7552</ID>
<type>BA_TRI_STATE</type>
<position>157,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5090 </input>
<output>
<ID>OUT_0</ID>5145 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7553</ID>
<type>AE_DFF_LOW</type>
<position>195,-2791.5</position>
<input>
<ID>IN_0</ID>5254 </input>
<output>
<ID>OUT_0</ID>5178 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7554</ID>
<type>AE_DFF_LOW</type>
<position>170,-2578.5</position>
<input>
<ID>IN_0</ID>5146 </input>
<output>
<ID>OUT_0</ID>5091 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7555</ID>
<type>BA_TRI_STATE</type>
<position>205,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5178 </input>
<output>
<ID>OUT_0</ID>5255 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7556</ID>
<type>BA_TRI_STATE</type>
<position>180,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5091 </input>
<output>
<ID>OUT_0</ID>5147 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7557</ID>
<type>AE_DFF_LOW</type>
<position>218,-2791.5</position>
<input>
<ID>IN_0</ID>5256 </input>
<output>
<ID>OUT_0</ID>5179 </output>
<input>
<ID>clock</ID>5180 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7558</ID>
<type>AE_DFF_LOW</type>
<position>195,-2578.5</position>
<input>
<ID>IN_0</ID>5148 </input>
<output>
<ID>OUT_0</ID>5092 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7559</ID>
<type>BA_TRI_STATE</type>
<position>228,-2802</position>
<input>
<ID>ENABLE_0</ID>5181 </input>
<input>
<ID>IN_0</ID>5179 </input>
<output>
<ID>OUT_0</ID>5257 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7560</ID>
<type>BA_TRI_STATE</type>
<position>205,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5092 </input>
<output>
<ID>OUT_0</ID>5149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7561</ID>
<type>AA_AND2</type>
<position>25.5,-2773.5</position>
<input>
<ID>IN_0</ID>5259 </input>
<input>
<ID>IN_1</ID>5266 </input>
<output>
<ID>OUT</ID>5190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7562</ID>
<type>AE_DFF_LOW</type>
<position>218,-2578.5</position>
<input>
<ID>IN_0</ID>5150 </input>
<output>
<ID>OUT_0</ID>5093 </output>
<input>
<ID>clock</ID>5094 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7563</ID>
<type>AA_AND2</type>
<position>37,-2783</position>
<input>
<ID>IN_0</ID>5259 </input>
<input>
<ID>IN_1</ID>5267 </input>
<output>
<ID>OUT</ID>5191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7564</ID>
<type>BA_TRI_STATE</type>
<position>228,-2589</position>
<input>
<ID>ENABLE_0</ID>5095 </input>
<input>
<ID>IN_0</ID>5093 </input>
<output>
<ID>OUT_0</ID>5151 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7565</ID>
<type>AE_DFF_LOW</type>
<position>53,-2772.5</position>
<input>
<ID>IN_0</ID>5242 </input>
<output>
<ID>OUT_0</ID>5182 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7566</ID>
<type>AA_AND2</type>
<position>25.5,-2713.5</position>
<input>
<ID>IN_0</ID>5159 </input>
<input>
<ID>IN_1</ID>5160 </input>
<output>
<ID>OUT</ID>5104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7567</ID>
<type>BA_TRI_STATE</type>
<position>63,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5182 </input>
<output>
<ID>OUT_0</ID>5243 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7568</ID>
<type>AA_AND2</type>
<position>36.5,-2723</position>
<input>
<ID>IN_0</ID>5159 </input>
<input>
<ID>IN_1</ID>5161 </input>
<output>
<ID>OUT</ID>5105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7569</ID>
<type>AE_DFF_LOW</type>
<position>76,-2772.5</position>
<input>
<ID>IN_0</ID>5244 </input>
<output>
<ID>OUT_0</ID>5183 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7570</ID>
<type>AE_DFF_LOW</type>
<position>53,-2712.5</position>
<input>
<ID>IN_0</ID>5136 </input>
<output>
<ID>OUT_0</ID>5096 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7571</ID>
<type>BA_TRI_STATE</type>
<position>86,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5183 </input>
<output>
<ID>OUT_0</ID>5245 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7572</ID>
<type>BA_TRI_STATE</type>
<position>63,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5096 </input>
<output>
<ID>OUT_0</ID>5137 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7573</ID>
<type>AE_DFF_LOW</type>
<position>101,-2772.5</position>
<input>
<ID>IN_0</ID>5246 </input>
<output>
<ID>OUT_0</ID>5184 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7574</ID>
<type>AE_DFF_LOW</type>
<position>76,-2712.5</position>
<input>
<ID>IN_0</ID>5138 </input>
<output>
<ID>OUT_0</ID>5097 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7575</ID>
<type>BA_TRI_STATE</type>
<position>111,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5184 </input>
<output>
<ID>OUT_0</ID>5247 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7576</ID>
<type>BA_TRI_STATE</type>
<position>86,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5097 </input>
<output>
<ID>OUT_0</ID>5139 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7577</ID>
<type>AE_DFF_LOW</type>
<position>124,-2772.5</position>
<input>
<ID>IN_0</ID>5248 </input>
<output>
<ID>OUT_0</ID>5185 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7578</ID>
<type>AE_DFF_LOW</type>
<position>101,-2712.5</position>
<input>
<ID>IN_0</ID>5140 </input>
<output>
<ID>OUT_0</ID>5098 </output>
<input>
<ID>clock</ID>5104 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7579</ID>
<type>BA_TRI_STATE</type>
<position>134,-2783</position>
<input>
<ID>ENABLE_0</ID>5191 </input>
<input>
<ID>IN_0</ID>5185 </input>
<output>
<ID>OUT_0</ID>5249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7580</ID>
<type>BA_TRI_STATE</type>
<position>111,-2723</position>
<input>
<ID>ENABLE_0</ID>5105 </input>
<input>
<ID>IN_0</ID>5098 </input>
<output>
<ID>OUT_0</ID>5141 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7581</ID>
<type>AE_DFF_LOW</type>
<position>147,-2772.5</position>
<input>
<ID>IN_0</ID>5250 </input>
<output>
<ID>OUT_0</ID>5186 </output>
<input>
<ID>clock</ID>5190 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7583</ID>
<type>AA_LABEL</type>
<position>274,-2730.5</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7584</ID>
<type>AE_DFF_LOW</type>
<position>115,-3104.5</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5329 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1434</ID>
<type>AA_AND2</type>
<position>30.5,-12.5</position>
<input>
<ID>IN_0</ID>1109 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1018 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7585</ID>
<type>BA_TRI_STATE</type>
<position>148,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5416 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7586</ID>
<type>BA_TRI_STATE</type>
<position>125,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5329 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7587</ID>
<type>AE_DFF_LOW</type>
<position>161,-3164.5</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5417 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7588</ID>
<type>AE_DFF_LOW</type>
<position>138,-3104.5</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5330 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1438</ID>
<type>AA_AND2</type>
<position>42,-22</position>
<input>
<ID>IN_0</ID>1109 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7589</ID>
<type>BA_TRI_STATE</type>
<position>171,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5417 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7590</ID>
<type>BA_TRI_STATE</type>
<position>148,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5330 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7591</ID>
<type>AE_DFF_LOW</type>
<position>186,-3164.5</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5418 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7592</ID>
<type>AE_DFF_LOW</type>
<position>161,-3104.5</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5331 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1442</ID>
<type>AE_DFF_LOW</type>
<position>58,-11.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1010 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7593</ID>
<type>BA_TRI_STATE</type>
<position>196,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5418 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7594</ID>
<type>BA_TRI_STATE</type>
<position>171,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5331 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7595</ID>
<type>AE_DFF_LOW</type>
<position>209,-3164.5</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5419 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7596</ID>
<type>AE_DFF_LOW</type>
<position>186,-3104.5</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5332 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7597</ID>
<type>BA_TRI_STATE</type>
<position>219,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5419 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1447</ID>
<type>BA_TRI_STATE</type>
<position>68,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1010 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7598</ID>
<type>BA_TRI_STATE</type>
<position>196,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5332 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7599</ID>
<type>AA_AND2</type>
<position>16.5,-3147</position>
<input>
<ID>IN_0</ID>5488 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7600</ID>
<type>AE_DFF_LOW</type>
<position>209,-3104.5</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5333 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7601</ID>
<type>AA_AND2</type>
<position>28,-3156.5</position>
<input>
<ID>IN_0</ID>5488 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7602</ID>
<type>BA_TRI_STATE</type>
<position>219,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5333 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7603</ID>
<type>AE_DFF_LOW</type>
<position>44,-3146</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5422 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7604</ID>
<type>AA_AND2</type>
<position>16.5,-3087</position>
<input>
<ID>IN_0</ID>5388 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5344 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7605</ID>
<type>BA_TRI_STATE</type>
<position>54,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5422 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7606</ID>
<type>AA_AND2</type>
<position>27.5,-3096.5</position>
<input>
<ID>IN_0</ID>5388 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7607</ID>
<type>AE_DFF_LOW</type>
<position>67,-3146</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5423 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7608</ID>
<type>AE_DFF_LOW</type>
<position>44,-3086</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5336 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7609</ID>
<type>BA_TRI_STATE</type>
<position>77,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5423 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7610</ID>
<type>BA_TRI_STATE</type>
<position>54,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5336 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7611</ID>
<type>AE_DFF_LOW</type>
<position>92,-3146</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5424 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7612</ID>
<type>AE_DFF_LOW</type>
<position>67,-3086</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5337 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1462</ID>
<type>AE_DFF_LOW</type>
<position>81,-11.5</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1011 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7613</ID>
<type>BA_TRI_STATE</type>
<position>102,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5424 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1463</ID>
<type>BA_TRI_STATE</type>
<position>91,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1011 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7614</ID>
<type>BA_TRI_STATE</type>
<position>77,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5337 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1464</ID>
<type>AE_DFF_LOW</type>
<position>106,-11.5</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1012 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7615</ID>
<type>AE_DFF_LOW</type>
<position>115,-3146</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5425 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1465</ID>
<type>BA_TRI_STATE</type>
<position>116,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1012 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7616</ID>
<type>AE_DFF_LOW</type>
<position>92,-3086</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5338 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1466</ID>
<type>AE_DFF_LOW</type>
<position>129,-11.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1013 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7617</ID>
<type>BA_TRI_STATE</type>
<position>125,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5425 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1467</ID>
<type>BA_TRI_STATE</type>
<position>139,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1013 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7618</ID>
<type>BA_TRI_STATE</type>
<position>102,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5338 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1468</ID>
<type>AE_DFF_LOW</type>
<position>152,-11.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1014 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7619</ID>
<type>AE_DFF_LOW</type>
<position>138,-3146</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5426 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1469</ID>
<type>BA_TRI_STATE</type>
<position>162,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1014 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7620</ID>
<type>AE_DFF_LOW</type>
<position>115,-3086</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5339 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1470</ID>
<type>AE_DFF_LOW</type>
<position>175,-11.5</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1015 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7621</ID>
<type>BA_TRI_STATE</type>
<position>148,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5426 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1471</ID>
<type>BA_TRI_STATE</type>
<position>185,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1015 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7622</ID>
<type>BA_TRI_STATE</type>
<position>125,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5339 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1472</ID>
<type>AE_DFF_LOW</type>
<position>200,-11.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1016 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7623</ID>
<type>AE_DFF_LOW</type>
<position>161,-3146</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5427 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1473</ID>
<type>BA_TRI_STATE</type>
<position>210,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1016 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7624</ID>
<type>AE_DFF_LOW</type>
<position>138,-3086</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5340 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1474</ID>
<type>AE_DFF_LOW</type>
<position>223,-11.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1017 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7625</ID>
<type>BA_TRI_STATE</type>
<position>171,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5427 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1475</ID>
<type>BA_TRI_STATE</type>
<position>233,-22</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1017 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7626</ID>
<type>BA_TRI_STATE</type>
<position>148,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5340 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1476</ID>
<type>AA_AND2</type>
<position>30.5,6</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1028 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7627</ID>
<type>AE_DFF_LOW</type>
<position>186,-3146</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5428 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1477</ID>
<type>AA_AND2</type>
<position>42,-3.5</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1029 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7628</ID>
<type>AE_DFF_LOW</type>
<position>161,-3086</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5341 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1478</ID>
<type>AE_DFF_LOW</type>
<position>58,7</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1020 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7629</ID>
<type>BA_TRI_STATE</type>
<position>196,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5428 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1479</ID>
<type>BA_TRI_STATE</type>
<position>68,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1020 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7630</ID>
<type>BA_TRI_STATE</type>
<position>171,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5341 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1480</ID>
<type>AE_DFF_LOW</type>
<position>81,7</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1021 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7631</ID>
<type>AE_DFF_LOW</type>
<position>209,-3146</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5429 </output>
<input>
<ID>clock</ID>5430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1481</ID>
<type>BA_TRI_STATE</type>
<position>91,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1021 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7632</ID>
<type>AE_DFF_LOW</type>
<position>186,-3086</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5342 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1482</ID>
<type>AE_DFF_LOW</type>
<position>106,7</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1022 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7633</ID>
<type>BA_TRI_STATE</type>
<position>219,-3156.5</position>
<input>
<ID>ENABLE_0</ID>5431 </input>
<input>
<ID>IN_0</ID>5429 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1483</ID>
<type>BA_TRI_STATE</type>
<position>116,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1022 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7634</ID>
<type>BA_TRI_STATE</type>
<position>196,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5342 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1484</ID>
<type>AE_DFF_LOW</type>
<position>129,7</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1023 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7635</ID>
<type>AA_AND2</type>
<position>16.5,-3281</position>
<input>
<ID>IN_0</ID>5495 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5440 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1485</ID>
<type>BA_TRI_STATE</type>
<position>139,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1023 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7636</ID>
<type>AE_DFF_LOW</type>
<position>209,-3086</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5343 </output>
<input>
<ID>clock</ID>5344 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1486</ID>
<type>AE_DFF_LOW</type>
<position>152,7</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1024 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7637</ID>
<type>AA_AND2</type>
<position>27.5,-3290.5</position>
<input>
<ID>IN_0</ID>5495 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5441 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1487</ID>
<type>BA_TRI_STATE</type>
<position>162,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1024 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7638</ID>
<type>BA_TRI_STATE</type>
<position>219,-3096.5</position>
<input>
<ID>ENABLE_0</ID>5345 </input>
<input>
<ID>IN_0</ID>5343 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1488</ID>
<type>AE_DFF_LOW</type>
<position>175,7</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1025 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7639</ID>
<type>AE_DFF_LOW</type>
<position>44,-3280</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5432 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1489</ID>
<type>BA_TRI_STATE</type>
<position>185,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1025 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7640</ID>
<type>AA_AND2</type>
<position>27.5,-3253</position>
<input>
<ID>IN_0</ID>5493 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5461 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1490</ID>
<type>AE_DFF_LOW</type>
<position>200,7</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1026 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7641</ID>
<type>AA_AND2</type>
<position>16.5,-3068</position>
<input>
<ID>IN_0</ID>5387 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1491</ID>
<type>BA_TRI_STATE</type>
<position>210,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1026 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7642</ID>
<type>BA_TRI_STATE</type>
<position>54,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5432 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1492</ID>
<type>AE_DFF_LOW</type>
<position>223,7</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1027 </output>
<input>
<ID>clock</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7643</ID>
<type>AA_AND2</type>
<position>27.5,-3077.5</position>
<input>
<ID>IN_0</ID>5387 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1493</ID>
<type>BA_TRI_STATE</type>
<position>233,-3.5</position>
<input>
<ID>ENABLE_0</ID>1029 </input>
<input>
<ID>IN_0</ID>1027 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7644</ID>
<type>AE_DFF_LOW</type>
<position>67,-3280</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5433 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1494</ID>
<type>AA_AND2</type>
<position>30.5,25</position>
<input>
<ID>IN_0</ID>1107 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1038 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7645</ID>
<type>AE_DFF_LOW</type>
<position>44,-3242.5</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5452 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1495</ID>
<type>AA_AND2</type>
<position>42,15.5</position>
<input>
<ID>IN_0</ID>1107 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1039 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7646</ID>
<type>AE_DFF_LOW</type>
<position>44,-3067</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5346 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1496</ID>
<type>AE_DFF_LOW</type>
<position>58,26</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1030 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7647</ID>
<type>BA_TRI_STATE</type>
<position>77,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5433 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1497</ID>
<type>BA_TRI_STATE</type>
<position>68,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1030 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7648</ID>
<type>BA_TRI_STATE</type>
<position>54,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5346 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1498</ID>
<type>AE_DFF_LOW</type>
<position>81,26</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1031 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7649</ID>
<type>AE_DFF_LOW</type>
<position>92,-3280</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5434 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1499</ID>
<type>BA_TRI_STATE</type>
<position>91,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1031 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7650</ID>
<type>BA_TRI_STATE</type>
<position>54,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5452 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1500</ID>
<type>AE_DFF_LOW</type>
<position>106,26</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1032 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7651</ID>
<type>AE_DFF_LOW</type>
<position>67,-3067</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5347 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1501</ID>
<type>BA_TRI_STATE</type>
<position>116,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1032 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7652</ID>
<type>BA_TRI_STATE</type>
<position>102,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5434 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1502</ID>
<type>AE_DFF_LOW</type>
<position>129,26</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1033 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7653</ID>
<type>BA_TRI_STATE</type>
<position>77,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5347 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1503</ID>
<type>BA_TRI_STATE</type>
<position>139,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1033 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7654</ID>
<type>AE_DFF_LOW</type>
<position>115,-3280</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5435 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1504</ID>
<type>AE_DFF_LOW</type>
<position>152,26</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1034 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7655</ID>
<type>AE_DFF_LOW</type>
<position>67,-3242.5</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5453 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1505</ID>
<type>BA_TRI_STATE</type>
<position>162,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1034 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7656</ID>
<type>AE_DFF_LOW</type>
<position>92,-3067</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5348 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1506</ID>
<type>AE_DFF_LOW</type>
<position>175,26</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1035 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7657</ID>
<type>BA_TRI_STATE</type>
<position>125,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5435 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1507</ID>
<type>BA_TRI_STATE</type>
<position>185,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1035 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7658</ID>
<type>BA_TRI_STATE</type>
<position>102,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5348 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1508</ID>
<type>AE_DFF_LOW</type>
<position>200,26</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1036 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7659</ID>
<type>AE_DFF_LOW</type>
<position>138,-3280</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5436 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1509</ID>
<type>BA_TRI_STATE</type>
<position>210,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1036 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7660</ID>
<type>BA_TRI_STATE</type>
<position>77,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5453 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1510</ID>
<type>AE_DFF_LOW</type>
<position>223,26</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1037 </output>
<input>
<ID>clock</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7661</ID>
<type>AE_DFF_LOW</type>
<position>115,-3067</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5349 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1511</ID>
<type>BA_TRI_STATE</type>
<position>233,15.5</position>
<input>
<ID>ENABLE_0</ID>1039 </input>
<input>
<ID>IN_0</ID>1037 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7662</ID>
<type>BA_TRI_STATE</type>
<position>148,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5436 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1512</ID>
<type>AA_AND2</type>
<position>30.5,43.5</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1048 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7663</ID>
<type>BA_TRI_STATE</type>
<position>125,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5349 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1513</ID>
<type>AA_AND2</type>
<position>42,34</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1049 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7664</ID>
<type>AE_DFF_LOW</type>
<position>161,-3280</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5437 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1514</ID>
<type>AE_DFF_LOW</type>
<position>58,44.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1040 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7665</ID>
<type>AE_DFF_LOW</type>
<position>92,-3242.5</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5454 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1515</ID>
<type>BA_TRI_STATE</type>
<position>68,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1040 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7666</ID>
<type>AE_DFF_LOW</type>
<position>138,-3067</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5350 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1516</ID>
<type>AE_DFF_LOW</type>
<position>81,44.5</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1041 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7667</ID>
<type>BA_TRI_STATE</type>
<position>171,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5437 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1517</ID>
<type>BA_TRI_STATE</type>
<position>91,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1041 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7668</ID>
<type>BA_TRI_STATE</type>
<position>148,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5350 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1518</ID>
<type>AE_DFF_LOW</type>
<position>106,44.5</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1042 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7669</ID>
<type>BA_TRI_STATE</type>
<position>102,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5454 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1519</ID>
<type>BA_TRI_STATE</type>
<position>116,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1042 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7670</ID>
<type>AE_DFF_LOW</type>
<position>161,-3067</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5351 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1520</ID>
<type>AE_DFF_LOW</type>
<position>129,44.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1043 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7671</ID>
<type>BA_TRI_STATE</type>
<position>171,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5351 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1521</ID>
<type>BA_TRI_STATE</type>
<position>139,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1043 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7672</ID>
<type>AE_DFF_LOW</type>
<position>115,-3242.5</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5455 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1522</ID>
<type>AE_DFF_LOW</type>
<position>152,44.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1044 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7673</ID>
<type>AE_DFF_LOW</type>
<position>186,-3067</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5352 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1523</ID>
<type>BA_TRI_STATE</type>
<position>162,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1044 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7674</ID>
<type>BA_TRI_STATE</type>
<position>196,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5352 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1524</ID>
<type>AE_DFF_LOW</type>
<position>175,44.5</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1045 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7675</ID>
<type>AE_DFF_LOW</type>
<position>209,-3067</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5353 </output>
<input>
<ID>clock</ID>5354 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1525</ID>
<type>BA_TRI_STATE</type>
<position>185,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1045 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7676</ID>
<type>BA_TRI_STATE</type>
<position>219,-3077.5</position>
<input>
<ID>ENABLE_0</ID>5355 </input>
<input>
<ID>IN_0</ID>5353 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1526</ID>
<type>AE_DFF_LOW</type>
<position>200,44.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1046 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7677</ID>
<type>AA_AND2</type>
<position>16.5,-3049.5</position>
<input>
<ID>IN_0</ID>5386 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1527</ID>
<type>BA_TRI_STATE</type>
<position>210,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1046 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7678</ID>
<type>AA_AND2</type>
<position>27.5,-3059</position>
<input>
<ID>IN_0</ID>5386 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5365 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1528</ID>
<type>AE_DFF_LOW</type>
<position>223,44.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1047 </output>
<input>
<ID>clock</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7679</ID>
<type>AE_DFF_LOW</type>
<position>44,-3048.5</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5356 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1529</ID>
<type>BA_TRI_STATE</type>
<position>233,34</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1047 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7680</ID>
<type>BA_TRI_STATE</type>
<position>54,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5356 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1530</ID>
<type>AA_AND2</type>
<position>30.5,-90.5</position>
<input>
<ID>IN_0</ID>1114 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1058 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7681</ID>
<type>AE_DFF_LOW</type>
<position>67,-3048.5</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5357 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1531</ID>
<type>AA_AND2</type>
<position>41.5,-100</position>
<input>
<ID>IN_0</ID>1114 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1059 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7682</ID>
<type>BA_TRI_STATE</type>
<position>77,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5357 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1532</ID>
<type>AE_DFF_LOW</type>
<position>58,-89.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1050 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7683</ID>
<type>AE_DFF_LOW</type>
<position>92,-3048.5</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5358 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1533</ID>
<type>BA_TRI_STATE</type>
<position>68,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1050 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7684</ID>
<type>BA_TRI_STATE</type>
<position>102,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5358 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1534</ID>
<type>AE_DFF_LOW</type>
<position>81,-89.5</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1051 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7685</ID>
<type>AE_DFF_LOW</type>
<position>115,-3048.5</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5359 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1535</ID>
<type>BA_TRI_STATE</type>
<position>91,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1051 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7686</ID>
<type>BA_TRI_STATE</type>
<position>125,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5359 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1536</ID>
<type>AE_DFF_LOW</type>
<position>106,-89.5</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1052 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7687</ID>
<type>AE_DFF_LOW</type>
<position>138,-3048.5</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5360 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1537</ID>
<type>BA_TRI_STATE</type>
<position>116,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1052 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7688</ID>
<type>BA_TRI_STATE</type>
<position>148,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5360 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1538</ID>
<type>AE_DFF_LOW</type>
<position>129,-89.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1053 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7689</ID>
<type>AE_DFF_LOW</type>
<position>161,-3048.5</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5361 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1539</ID>
<type>BA_TRI_STATE</type>
<position>139,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1053 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7690</ID>
<type>BA_TRI_STATE</type>
<position>171,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5361 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1540</ID>
<type>AE_DFF_LOW</type>
<position>152,-89.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1054 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7691</ID>
<type>AE_DFF_LOW</type>
<position>186,-3048.5</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5362 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1541</ID>
<type>BA_TRI_STATE</type>
<position>162,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1054 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7692</ID>
<type>BA_TRI_STATE</type>
<position>196,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5362 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1542</ID>
<type>AE_DFF_LOW</type>
<position>175,-89.5</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1055 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7693</ID>
<type>AE_DFF_LOW</type>
<position>209,-3048.5</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5363 </output>
<input>
<ID>clock</ID>5364 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1543</ID>
<type>BA_TRI_STATE</type>
<position>185,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1055 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7694</ID>
<type>BA_TRI_STATE</type>
<position>219,-3059</position>
<input>
<ID>ENABLE_0</ID>5365 </input>
<input>
<ID>IN_0</ID>5363 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1544</ID>
<type>AE_DFF_LOW</type>
<position>200,-89.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1056 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7695</ID>
<type>HA_JUNC_2</type>
<position>35.5,-2962</position>
<input>
<ID>N_in0</ID>5366 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1545</ID>
<type>BA_TRI_STATE</type>
<position>210,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1056 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7696</ID>
<type>HA_JUNC_2</type>
<position>58.5,-2961.5</position>
<input>
<ID>N_in0</ID>5367 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1546</ID>
<type>AE_DFF_LOW</type>
<position>223,-89.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1057 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7697</ID>
<type>HA_JUNC_2</type>
<position>61.5,-2962</position>
<input>
<ID>N_in0</ID>5368 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1547</ID>
<type>BA_TRI_STATE</type>
<position>233,-100</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1057 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7698</ID>
<type>HA_JUNC_2</type>
<position>81,-2961.5</position>
<input>
<ID>N_in0</ID>5369 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1548</ID>
<type>AA_AND2</type>
<position>30.5,-72</position>
<input>
<ID>IN_0</ID>1113 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7699</ID>
<type>HA_JUNC_2</type>
<position>84.5,-2961.5</position>
<input>
<ID>N_in0</ID>5370 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1549</ID>
<type>AA_AND2</type>
<position>41.5,-81.5</position>
<input>
<ID>IN_0</ID>1113 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1069 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7700</ID>
<type>HA_JUNC_2</type>
<position>105.5,-2962</position>
<input>
<ID>N_in0</ID>5371 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1550</ID>
<type>AE_DFF_LOW</type>
<position>58,-71</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1060 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7701</ID>
<type>HA_JUNC_2</type>
<position>109.5,-2961.5</position>
<input>
<ID>N_in0</ID>5372 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1551</ID>
<type>BA_TRI_STATE</type>
<position>68,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1060 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7702</ID>
<type>HA_JUNC_2</type>
<position>128,-2961.5</position>
<input>
<ID>N_in0</ID>5373 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1552</ID>
<type>AE_DFF_LOW</type>
<position>81,-71</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1061 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7703</ID>
<type>HA_JUNC_2</type>
<position>132,-2961.5</position>
<input>
<ID>N_in0</ID>5374 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1553</ID>
<type>BA_TRI_STATE</type>
<position>91,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1061 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7704</ID>
<type>HA_JUNC_2</type>
<position>151,-2961.5</position>
<input>
<ID>N_in0</ID>5375 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1554</ID>
<type>AE_DFF_LOW</type>
<position>106,-71</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1062 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7705</ID>
<type>HA_JUNC_2</type>
<position>156,-2961.5</position>
<input>
<ID>N_in0</ID>5376 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1555</ID>
<type>BA_TRI_STATE</type>
<position>116,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1062 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7706</ID>
<type>HA_JUNC_2</type>
<position>178.5,-2961.5</position>
<input>
<ID>N_in0</ID>5378 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1556</ID>
<type>AE_DFF_LOW</type>
<position>129,-71</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1063 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7707</ID>
<type>HA_JUNC_2</type>
<position>174,-2961.5</position>
<input>
<ID>N_in0</ID>5377 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1557</ID>
<type>BA_TRI_STATE</type>
<position>139,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1063 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7708</ID>
<type>HA_JUNC_2</type>
<position>199.5,-2962</position>
<input>
<ID>N_in0</ID>5379 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1558</ID>
<type>AE_DFF_LOW</type>
<position>152,-71</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1064 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7709</ID>
<type>HA_JUNC_2</type>
<position>224,-2963</position>
<input>
<ID>N_in0</ID>5381 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1559</ID>
<type>BA_TRI_STATE</type>
<position>162,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1064 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7710</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3129</position>
<input>
<ID>N_in0</ID>5500 </input>
<input>
<ID>N_in1</ID>5366 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1560</ID>
<type>AE_DFF_LOW</type>
<position>175,-71</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1065 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7711</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3128.5</position>
<input>
<ID>N_in0</ID>5501 </input>
<input>
<ID>N_in1</ID>5367 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1561</ID>
<type>BA_TRI_STATE</type>
<position>185,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1065 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7712</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3128.5</position>
<input>
<ID>N_in0</ID>5502 </input>
<input>
<ID>N_in1</ID>5368 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1562</ID>
<type>AE_DFF_LOW</type>
<position>200,-71</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1066 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7713</ID>
<type>HA_JUNC_2</type>
<position>81,-3128.5</position>
<input>
<ID>N_in0</ID>5503 </input>
<input>
<ID>N_in1</ID>5369 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1563</ID>
<type>BA_TRI_STATE</type>
<position>210,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1066 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7714</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3128.5</position>
<input>
<ID>N_in0</ID>5504 </input>
<input>
<ID>N_in1</ID>5370 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1564</ID>
<type>AE_DFF_LOW</type>
<position>223,-71</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1067 </output>
<input>
<ID>clock</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7715</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3128.5</position>
<input>
<ID>N_in0</ID>5505 </input>
<input>
<ID>N_in1</ID>5371 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1565</ID>
<type>BA_TRI_STATE</type>
<position>233,-81.5</position>
<input>
<ID>ENABLE_0</ID>1069 </input>
<input>
<ID>IN_0</ID>1067 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7716</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3128.5</position>
<input>
<ID>N_in0</ID>5506 </input>
<input>
<ID>N_in1</ID>5372 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1566</ID>
<type>AA_AND2</type>
<position>30.5,-53</position>
<input>
<ID>IN_0</ID>1112 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1078 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7717</ID>
<type>HA_JUNC_2</type>
<position>128,-3128.5</position>
<input>
<ID>N_in0</ID>5507 </input>
<input>
<ID>N_in1</ID>5373 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1567</ID>
<type>AA_AND2</type>
<position>41.5,-62.5</position>
<input>
<ID>IN_0</ID>1112 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1079 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7718</ID>
<type>HA_JUNC_2</type>
<position>132,-3128.5</position>
<input>
<ID>N_in0</ID>5508 </input>
<input>
<ID>N_in1</ID>5374 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1568</ID>
<type>AE_DFF_LOW</type>
<position>58,-52</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1070 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7719</ID>
<type>HA_JUNC_2</type>
<position>151,-3128</position>
<input>
<ID>N_in0</ID>5509 </input>
<input>
<ID>N_in1</ID>5375 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1569</ID>
<type>BA_TRI_STATE</type>
<position>68,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1070 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7720</ID>
<type>HA_JUNC_2</type>
<position>156,-3128</position>
<input>
<ID>N_in0</ID>5510 </input>
<input>
<ID>N_in1</ID>5376 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1570</ID>
<type>AE_DFF_LOW</type>
<position>81,-52</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1071 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7721</ID>
<type>HA_JUNC_2</type>
<position>174,-3127.5</position>
<input>
<ID>N_in0</ID>5511 </input>
<input>
<ID>N_in1</ID>5377 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1571</ID>
<type>BA_TRI_STATE</type>
<position>91,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1071 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7722</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3127.5</position>
<input>
<ID>N_in0</ID>5512 </input>
<input>
<ID>N_in1</ID>5378 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1572</ID>
<type>AE_DFF_LOW</type>
<position>106,-52</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1072 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7723</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3127</position>
<input>
<ID>N_in0</ID>5513 </input>
<input>
<ID>N_in1</ID>5379 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1573</ID>
<type>BA_TRI_STATE</type>
<position>116,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1072 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7724</ID>
<type>HA_JUNC_2</type>
<position>203,-3127</position>
<input>
<ID>N_in0</ID>5514 </input>
<input>
<ID>N_in1</ID>5380 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1574</ID>
<type>AE_DFF_LOW</type>
<position>129,-52</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1073 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7725</ID>
<type>HA_JUNC_2</type>
<position>203,-2962</position>
<input>
<ID>N_in0</ID>5380 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1575</ID>
<type>BA_TRI_STATE</type>
<position>139,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1073 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7726</ID>
<type>HA_JUNC_2</type>
<position>224,-3127</position>
<input>
<ID>N_in0</ID>5515 </input>
<input>
<ID>N_in1</ID>5381 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1576</ID>
<type>AE_DFF_LOW</type>
<position>152,-52</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1074 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7727</ID>
<type>HA_JUNC_2</type>
<position>22.5,-2962</position>
<input>
<ID>N_in0</ID>5391 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1577</ID>
<type>BA_TRI_STATE</type>
<position>162,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1074 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7728</ID>
<type>HA_JUNC_2</type>
<position>12.5,-2962</position>
<input>
<ID>N_in0</ID>5390 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1578</ID>
<type>AE_DFF_LOW</type>
<position>175,-52</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1075 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7729</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3129</position>
<input>
<ID>N_in0</ID>5499 </input>
<input>
<ID>N_in1</ID>5391 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1579</ID>
<type>BA_TRI_STATE</type>
<position>185,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1075 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7730</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3129</position>
<input>
<ID>N_in0</ID>5498 </input>
<input>
<ID>N_in1</ID>5390 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1580</ID>
<type>AE_DFF_LOW</type>
<position>200,-52</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1076 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7731</ID>
<type>AA_LABEL</type>
<position>3.5,-2962.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1581</ID>
<type>BA_TRI_STATE</type>
<position>210,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1076 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7732</ID>
<type>BI_DECODER_4x16</type>
<position>-136,-3129.5</position>
<output>
<ID>OUT_0</ID>5495 </output>
<output>
<ID>OUT_1</ID>5494 </output>
<output>
<ID>OUT_10</ID>5387 </output>
<output>
<ID>OUT_11</ID>5386 </output>
<output>
<ID>OUT_12</ID>5385 </output>
<output>
<ID>OUT_13</ID>5384 </output>
<output>
<ID>OUT_14</ID>5383 </output>
<output>
<ID>OUT_15</ID>5382 </output>
<output>
<ID>OUT_2</ID>5493 </output>
<output>
<ID>OUT_3</ID>5492 </output>
<output>
<ID>OUT_4</ID>5491 </output>
<output>
<ID>OUT_5</ID>5490 </output>
<output>
<ID>OUT_6</ID>5489 </output>
<output>
<ID>OUT_7</ID>5488 </output>
<output>
<ID>OUT_8</ID>5389 </output>
<output>
<ID>OUT_9</ID>5388 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1582</ID>
<type>AE_DFF_LOW</type>
<position>223,-52</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1077 </output>
<input>
<ID>clock</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7733</ID>
<type>AE_DFF_LOW</type>
<position>186,-3280</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5438 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1583</ID>
<type>BA_TRI_STATE</type>
<position>233,-62.5</position>
<input>
<ID>ENABLE_0</ID>1079 </input>
<input>
<ID>IN_0</ID>1077 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7734</ID>
<type>BA_TRI_STATE</type>
<position>196,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5438 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1584</ID>
<type>AA_AND2</type>
<position>30.5,-34.5</position>
<input>
<ID>IN_0</ID>1111 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1088 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7735</ID>
<type>AE_DFF_LOW</type>
<position>209,-3280</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5439 </output>
<input>
<ID>clock</ID>5440 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1585</ID>
<type>AA_AND2</type>
<position>41.5,-44</position>
<input>
<ID>IN_0</ID>1111 </input>
<input>
<ID>IN_1</ID>1118 </input>
<output>
<ID>OUT</ID>1089 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7736</ID>
<type>BA_TRI_STATE</type>
<position>219,-3290.5</position>
<input>
<ID>ENABLE_0</ID>5441 </input>
<input>
<ID>IN_0</ID>5439 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1586</ID>
<type>AE_DFF_LOW</type>
<position>58,-33.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1080 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7737</ID>
<type>AA_AND2</type>
<position>16.5,-3262.5</position>
<input>
<ID>IN_0</ID>5494 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1587</ID>
<type>BA_TRI_STATE</type>
<position>68,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1080 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7738</ID>
<type>AA_AND2</type>
<position>27.5,-3272</position>
<input>
<ID>IN_0</ID>5494 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1588</ID>
<type>AE_DFF_LOW</type>
<position>81,-33.5</position>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1081 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7739</ID>
<type>AE_DFF_LOW</type>
<position>44,-3261.5</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5442 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1589</ID>
<type>BA_TRI_STATE</type>
<position>91,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1081 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7740</ID>
<type>BA_TRI_STATE</type>
<position>54,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5442 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1590</ID>
<type>AE_DFF_LOW</type>
<position>106,-33.5</position>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1082 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7741</ID>
<type>AE_DFF_LOW</type>
<position>67,-3261.5</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5443 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1591</ID>
<type>BA_TRI_STATE</type>
<position>116,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1082 </input>
<output>
<ID>OUT_0</ID>1095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7742</ID>
<type>BA_TRI_STATE</type>
<position>77,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5443 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1592</ID>
<type>AE_DFF_LOW</type>
<position>129,-33.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1083 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7743</ID>
<type>AE_DFF_LOW</type>
<position>92,-3261.5</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5444 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1593</ID>
<type>BA_TRI_STATE</type>
<position>139,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1083 </input>
<output>
<ID>OUT_0</ID>1097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7744</ID>
<type>BA_TRI_STATE</type>
<position>102,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5444 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1594</ID>
<type>AE_DFF_LOW</type>
<position>152,-33.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1084 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7745</ID>
<type>AE_DFF_LOW</type>
<position>115,-3261.5</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5445 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1595</ID>
<type>BA_TRI_STATE</type>
<position>162,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1084 </input>
<output>
<ID>OUT_0</ID>1099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7746</ID>
<type>BA_TRI_STATE</type>
<position>125,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5445 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1596</ID>
<type>AE_DFF_LOW</type>
<position>175,-33.5</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1085 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7747</ID>
<type>AE_DFF_LOW</type>
<position>138,-3261.5</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5446 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1597</ID>
<type>BA_TRI_STATE</type>
<position>185,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1085 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7748</ID>
<type>BA_TRI_STATE</type>
<position>148,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5446 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1598</ID>
<type>AE_DFF_LOW</type>
<position>200,-33.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<output>
<ID>OUT_0</ID>1086 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7749</ID>
<type>AE_DFF_LOW</type>
<position>161,-3261.5</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5447 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1599</ID>
<type>BA_TRI_STATE</type>
<position>210,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1086 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7750</ID>
<type>BA_TRI_STATE</type>
<position>171,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5447 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1600</ID>
<type>AE_DFF_LOW</type>
<position>223,-33.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<output>
<ID>OUT_0</ID>1087 </output>
<input>
<ID>clock</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7751</ID>
<type>AE_DFF_LOW</type>
<position>186,-3261.5</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5448 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1601</ID>
<type>BA_TRI_STATE</type>
<position>233,-44</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1087 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7752</ID>
<type>BA_TRI_STATE</type>
<position>196,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5448 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7753</ID>
<type>AE_DFF_LOW</type>
<position>209,-3261.5</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5449 </output>
<input>
<ID>clock</ID>5450 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1603</ID>
<type>HA_JUNC_2</type>
<position>49.5,53</position>
<input>
<ID>N_in0</ID>1090 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7754</ID>
<type>BA_TRI_STATE</type>
<position>219,-3272</position>
<input>
<ID>ENABLE_0</ID>5451 </input>
<input>
<ID>IN_0</ID>5449 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7755</ID>
<type>AA_AND2</type>
<position>16.5,-3243.5</position>
<input>
<ID>IN_0</ID>5493 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5460 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1605</ID>
<type>HA_JUNC_2</type>
<position>72.5,53.5</position>
<input>
<ID>N_in0</ID>1091 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7756</ID>
<type>BA_TRI_STATE</type>
<position>125,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5455 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1606</ID>
<type>HA_JUNC_2</type>
<position>75.5,53</position>
<input>
<ID>N_in0</ID>1092 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7757</ID>
<type>AE_DFF_LOW</type>
<position>138,-3242.5</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5456 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1607</ID>
<type>HA_JUNC_2</type>
<position>95,53.5</position>
<input>
<ID>N_in0</ID>1093 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7758</ID>
<type>BA_TRI_STATE</type>
<position>148,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5456 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1608</ID>
<type>HA_JUNC_2</type>
<position>98.5,53.5</position>
<input>
<ID>N_in0</ID>1094 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7759</ID>
<type>AE_DFF_LOW</type>
<position>161,-3242.5</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5457 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1609</ID>
<type>HA_JUNC_2</type>
<position>119.5,53</position>
<input>
<ID>N_in0</ID>1095 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7760</ID>
<type>BA_TRI_STATE</type>
<position>171,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5457 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1610</ID>
<type>HA_JUNC_2</type>
<position>123.5,53.5</position>
<input>
<ID>N_in0</ID>1096 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7761</ID>
<type>AE_DFF_LOW</type>
<position>186,-3242.5</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5458 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1611</ID>
<type>HA_JUNC_2</type>
<position>142,53.5</position>
<input>
<ID>N_in0</ID>1097 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7762</ID>
<type>BA_TRI_STATE</type>
<position>196,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5458 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1612</ID>
<type>HA_JUNC_2</type>
<position>146,53.5</position>
<input>
<ID>N_in0</ID>1098 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7763</ID>
<type>AA_AND2</type>
<position>16.5,-3027.5</position>
<input>
<ID>IN_0</ID>5385 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5294 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1613</ID>
<type>HA_JUNC_2</type>
<position>165,53.5</position>
<input>
<ID>N_in0</ID>1099 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7764</ID>
<type>AE_DFF_LOW</type>
<position>209,-3242.5</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5459 </output>
<input>
<ID>clock</ID>5460 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1614</ID>
<type>HA_JUNC_2</type>
<position>170,53.5</position>
<input>
<ID>N_in0</ID>1100 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7765</ID>
<type>BA_TRI_STATE</type>
<position>219,-3253</position>
<input>
<ID>ENABLE_0</ID>5461 </input>
<input>
<ID>IN_0</ID>5459 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1615</ID>
<type>HA_JUNC_2</type>
<position>192.5,53.5</position>
<input>
<ID>N_in0</ID>1102 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7766</ID>
<type>AA_AND2</type>
<position>16.5,-3225</position>
<input>
<ID>IN_0</ID>5492 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5470 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1616</ID>
<type>HA_JUNC_2</type>
<position>188,53.5</position>
<input>
<ID>N_in0</ID>1101 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7767</ID>
<type>AA_AND2</type>
<position>27.5,-3234.5</position>
<input>
<ID>IN_0</ID>5492 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5471 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1617</ID>
<type>HA_JUNC_2</type>
<position>213.5,53</position>
<input>
<ID>N_in0</ID>1103 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7768</ID>
<type>AA_AND2</type>
<position>28,-3037</position>
<input>
<ID>IN_0</ID>5385 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5295 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1618</ID>
<type>HA_JUNC_2</type>
<position>238,52</position>
<input>
<ID>N_in0</ID>1105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7769</ID>
<type>AE_DFF_LOW</type>
<position>44,-3224</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5462 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7770</ID>
<type>BA_TRI_STATE</type>
<position>54,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5462 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7771</ID>
<type>AE_DFF_LOW</type>
<position>67,-3224</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5463 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7772</ID>
<type>BA_TRI_STATE</type>
<position>77,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5463 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7773</ID>
<type>AE_DFF_LOW</type>
<position>44,-3026.5</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5286 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7774</ID>
<type>AE_DFF_LOW</type>
<position>92,-3224</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5464 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7775</ID>
<type>BA_TRI_STATE</type>
<position>102,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5464 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7776</ID>
<type>AE_DFF_LOW</type>
<position>115,-3224</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5465 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7777</ID>
<type>BA_TRI_STATE</type>
<position>125,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5465 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7778</ID>
<type>AE_DFF_LOW</type>
<position>138,-3224</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5466 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7779</ID>
<type>BA_TRI_STATE</type>
<position>54,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5286 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7780</ID>
<type>BA_TRI_STATE</type>
<position>148,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5466 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7781</ID>
<type>AE_DFF_LOW</type>
<position>161,-3224</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5467 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7782</ID>
<type>BA_TRI_STATE</type>
<position>171,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5467 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7783</ID>
<type>AE_DFF_LOW</type>
<position>186,-3224</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5468 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7784</ID>
<type>BA_TRI_STATE</type>
<position>196,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5468 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7785</ID>
<type>AE_DFF_LOW</type>
<position>209,-3224</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5469 </output>
<input>
<ID>clock</ID>5470 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1635</ID>
<type>HA_JUNC_2</type>
<position>49.5,-114</position>
<input>
<ID>N_in0</ID>3200 </input>
<input>
<ID>N_in1</ID>1090 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7786</ID>
<type>BA_TRI_STATE</type>
<position>219,-3234.5</position>
<input>
<ID>ENABLE_0</ID>5471 </input>
<input>
<ID>IN_0</ID>5469 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1636</ID>
<type>HA_JUNC_2</type>
<position>72.5,-113.5</position>
<input>
<ID>N_in0</ID>3201 </input>
<input>
<ID>N_in1</ID>1091 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7787</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3137.5</position>
<input>
<ID>N_in0</ID>5472 </input>
<input>
<ID>N_in1</ID>5500 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1637</ID>
<type>HA_JUNC_2</type>
<position>75.5,-113.5</position>
<input>
<ID>N_in0</ID>3202 </input>
<input>
<ID>N_in1</ID>1092 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7788</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3137</position>
<input>
<ID>N_in0</ID>5473 </input>
<input>
<ID>N_in1</ID>5501 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1638</ID>
<type>HA_JUNC_2</type>
<position>95,-113.5</position>
<input>
<ID>N_in0</ID>3203 </input>
<input>
<ID>N_in1</ID>1093 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7789</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3137.5</position>
<input>
<ID>N_in0</ID>5474 </input>
<input>
<ID>N_in1</ID>5502 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1639</ID>
<type>HA_JUNC_2</type>
<position>98.5,-113.5</position>
<input>
<ID>N_in0</ID>3204 </input>
<input>
<ID>N_in1</ID>1094 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7790</ID>
<type>HA_JUNC_2</type>
<position>81,-3137</position>
<input>
<ID>N_in0</ID>5475 </input>
<input>
<ID>N_in1</ID>5503 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1640</ID>
<type>HA_JUNC_2</type>
<position>119.5,-113.5</position>
<input>
<ID>N_in0</ID>3205 </input>
<input>
<ID>N_in1</ID>1095 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7791</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3137</position>
<input>
<ID>N_in0</ID>5476 </input>
<input>
<ID>N_in1</ID>5504 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1641</ID>
<type>HA_JUNC_2</type>
<position>123.5,-113.5</position>
<input>
<ID>N_in0</ID>3206 </input>
<input>
<ID>N_in1</ID>1096 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7792</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3137.5</position>
<input>
<ID>N_in0</ID>5477 </input>
<input>
<ID>N_in1</ID>5505 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1642</ID>
<type>HA_JUNC_2</type>
<position>142,-113.5</position>
<input>
<ID>N_in0</ID>3207 </input>
<input>
<ID>N_in1</ID>1097 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7793</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3137</position>
<input>
<ID>N_in0</ID>5478 </input>
<input>
<ID>N_in1</ID>5506 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1643</ID>
<type>HA_JUNC_2</type>
<position>146,-113.5</position>
<input>
<ID>N_in0</ID>3208 </input>
<input>
<ID>N_in1</ID>1098 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7794</ID>
<type>HA_JUNC_2</type>
<position>128,-3137</position>
<input>
<ID>N_in0</ID>5479 </input>
<input>
<ID>N_in1</ID>5507 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1644</ID>
<type>HA_JUNC_2</type>
<position>165,-113</position>
<input>
<ID>N_in0</ID>3209 </input>
<input>
<ID>N_in1</ID>1099 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7795</ID>
<type>AE_DFF_LOW</type>
<position>67,-3026.5</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5287 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1645</ID>
<type>HA_JUNC_2</type>
<position>170,-113</position>
<input>
<ID>N_in0</ID>3210 </input>
<input>
<ID>N_in1</ID>1100 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7796</ID>
<type>HA_JUNC_2</type>
<position>132,-3137</position>
<input>
<ID>N_in0</ID>5480 </input>
<input>
<ID>N_in1</ID>5508 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1646</ID>
<type>HA_JUNC_2</type>
<position>188,-112.5</position>
<input>
<ID>N_in0</ID>3211 </input>
<input>
<ID>N_in1</ID>1101 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7797</ID>
<type>BA_TRI_STATE</type>
<position>77,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5287 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1647</ID>
<type>HA_JUNC_2</type>
<position>192.5,-112.5</position>
<input>
<ID>N_in0</ID>3212 </input>
<input>
<ID>N_in1</ID>1102 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7798</ID>
<type>HA_JUNC_2</type>
<position>151,-3137</position>
<input>
<ID>N_in0</ID>5481 </input>
<input>
<ID>N_in1</ID>5509 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1648</ID>
<type>HA_JUNC_2</type>
<position>213.5,-112</position>
<input>
<ID>N_in0</ID>3213 </input>
<input>
<ID>N_in1</ID>1103 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7799</ID>
<type>AE_DFF_LOW</type>
<position>92,-3026.5</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5288 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1649</ID>
<type>HA_JUNC_2</type>
<position>217,-112</position>
<input>
<ID>N_in0</ID>3214 </input>
<input>
<ID>N_in1</ID>1104 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7800</ID>
<type>HA_JUNC_2</type>
<position>156,-3137</position>
<input>
<ID>N_in0</ID>5482 </input>
<input>
<ID>N_in1</ID>5510 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7801</ID>
<type>BA_TRI_STATE</type>
<position>102,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5288 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1651</ID>
<type>HA_JUNC_2</type>
<position>217,53</position>
<input>
<ID>N_in0</ID>1104 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7802</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3137</position>
<input>
<ID>N_in0</ID>5484 </input>
<input>
<ID>N_in1</ID>5512 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7803</ID>
<type>AE_DFF_LOW</type>
<position>115,-3026.5</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5289 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1653</ID>
<type>HA_JUNC_2</type>
<position>238,-112</position>
<input>
<ID>N_in0</ID>3215 </input>
<input>
<ID>N_in1</ID>1105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7804</ID>
<type>HA_JUNC_2</type>
<position>174,-3137</position>
<input>
<ID>N_in0</ID>5483 </input>
<input>
<ID>N_in1</ID>5511 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7805</ID>
<type>BA_TRI_STATE</type>
<position>125,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5289 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7806</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3137.5</position>
<input>
<ID>N_in0</ID>5485 </input>
<input>
<ID>N_in1</ID>5513 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7807</ID>
<type>AE_DFF_LOW</type>
<position>138,-3026.5</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5290 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1657</ID>
<type>HA_JUNC_2</type>
<position>36.5,53</position>
<input>
<ID>N_in0</ID>1118 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7808</ID>
<type>HA_JUNC_2</type>
<position>224,-3138.5</position>
<input>
<ID>N_in0</ID>5487 </input>
<input>
<ID>N_in1</ID>5515 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1658</ID>
<type>HA_JUNC_2</type>
<position>26.5,53</position>
<input>
<ID>N_in0</ID>1117 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7809</ID>
<type>BA_TRI_STATE</type>
<position>148,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5290 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1659</ID>
<type>HA_JUNC_2</type>
<position>36.5,-114</position>
<input>
<ID>N_in0</ID>3199 </input>
<input>
<ID>N_in1</ID>1118 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7810</ID>
<type>AA_AND2</type>
<position>16.5,-3203</position>
<input>
<ID>IN_0</ID>5491 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5400 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1660</ID>
<type>HA_JUNC_2</type>
<position>26.5,-114</position>
<input>
<ID>N_in0</ID>3198 </input>
<input>
<ID>N_in1</ID>1117 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7811</ID>
<type>AE_DFF_LOW</type>
<position>161,-3026.5</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5291 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7812</ID>
<type>AA_AND2</type>
<position>28,-3212.5</position>
<input>
<ID>IN_0</ID>5491 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1662</ID>
<type>AA_LABEL</type>
<position>17.5,52.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7813</ID>
<type>BA_TRI_STATE</type>
<position>171,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5291 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7814</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3304.5</position>
<input>
<ID>N_in1</ID>5472 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1664</ID>
<type>BI_DECODER_4x16</type>
<position>-122,-114.5</position>
<output>
<ID>OUT_0</ID>3195 </output>
<output>
<ID>OUT_1</ID>3194 </output>
<output>
<ID>OUT_10</ID>1112 </output>
<output>
<ID>OUT_11</ID>1111 </output>
<output>
<ID>OUT_12</ID>1109 </output>
<output>
<ID>OUT_13</ID>1108 </output>
<output>
<ID>OUT_14</ID>1107 </output>
<output>
<ID>OUT_15</ID>1106 </output>
<output>
<ID>OUT_2</ID>3193 </output>
<output>
<ID>OUT_3</ID>3192 </output>
<output>
<ID>OUT_4</ID>3191 </output>
<output>
<ID>OUT_5</ID>3190 </output>
<output>
<ID>OUT_6</ID>3189 </output>
<output>
<ID>OUT_7</ID>3188 </output>
<output>
<ID>OUT_8</ID>1114 </output>
<output>
<ID>OUT_9</ID>1113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7815</ID>
<type>AE_DFF_LOW</type>
<position>186,-3026.5</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5292 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1665</ID>
<type>AE_DFF_LOW</type>
<position>200,-265</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>1165 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7816</ID>
<type>AE_DFF_LOW</type>
<position>44,-3202</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5392 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1666</ID>
<type>BA_TRI_STATE</type>
<position>210,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1165 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7817</ID>
<type>BA_TRI_STATE</type>
<position>196,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5292 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1667</ID>
<type>AE_DFF_LOW</type>
<position>223,-265</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>1166 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7818</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3304</position>
<input>
<ID>N_in1</ID>5473 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1668</ID>
<type>BA_TRI_STATE</type>
<position>233,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1166 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7819</ID>
<type>AE_DFF_LOW</type>
<position>209,-3026.5</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5293 </output>
<input>
<ID>clock</ID>5294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1669</ID>
<type>AA_AND2</type>
<position>30.5,-247.5</position>
<input>
<ID>IN_0</ID>3194 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>1642 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7820</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3304</position>
<input>
<ID>N_in1</ID>5474 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1670</ID>
<type>AA_AND2</type>
<position>41.5,-257</position>
<input>
<ID>IN_0</ID>3194 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>1643 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7821</ID>
<type>BA_TRI_STATE</type>
<position>219,-3037</position>
<input>
<ID>ENABLE_0</ID>5295 </input>
<input>
<ID>IN_0</ID>5293 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1671</ID>
<type>AE_DFF_LOW</type>
<position>58,-246.5</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1169 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7822</ID>
<type>HA_JUNC_2</type>
<position>81,-3304</position>
<input>
<ID>N_in1</ID>5475 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1672</ID>
<type>BA_TRI_STATE</type>
<position>68,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1169 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7823</ID>
<type>AA_AND2</type>
<position>16.5,-3009</position>
<input>
<ID>IN_0</ID>5384 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5304 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1673</ID>
<type>AE_DFF_LOW</type>
<position>81,-246.5</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1170 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7824</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3304</position>
<input>
<ID>N_in1</ID>5476 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1674</ID>
<type>BA_TRI_STATE</type>
<position>91,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1170 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7825</ID>
<type>AA_AND2</type>
<position>28,-3018.5</position>
<input>
<ID>IN_0</ID>5384 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1675</ID>
<type>AE_DFF_LOW</type>
<position>106,-246.5</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1171 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7826</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3304</position>
<input>
<ID>N_in1</ID>5477 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1676</ID>
<type>BA_TRI_STATE</type>
<position>116,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1171 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7827</ID>
<type>AE_DFF_LOW</type>
<position>44,-3008</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5296 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1677</ID>
<type>AE_DFF_LOW</type>
<position>129,-246.5</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1172 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7828</ID>
<type>BA_TRI_STATE</type>
<position>54,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5392 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1678</ID>
<type>BA_TRI_STATE</type>
<position>139,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1172 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7829</ID>
<type>BA_TRI_STATE</type>
<position>54,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5296 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1679</ID>
<type>AE_DFF_LOW</type>
<position>152,-246.5</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1173 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7830</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3304</position>
<input>
<ID>N_in1</ID>5478 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1680</ID>
<type>BA_TRI_STATE</type>
<position>162,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1173 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7831</ID>
<type>AE_DFF_LOW</type>
<position>67,-3008</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5297 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1681</ID>
<type>AE_DFF_LOW</type>
<position>175,-246.5</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>1174 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7832</ID>
<type>HA_JUNC_2</type>
<position>128,-3304</position>
<input>
<ID>N_in1</ID>5479 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1682</ID>
<type>BA_TRI_STATE</type>
<position>185,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1174 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7833</ID>
<type>BA_TRI_STATE</type>
<position>77,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5297 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1683</ID>
<type>AE_DFF_LOW</type>
<position>200,-246.5</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>1175 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7834</ID>
<type>HA_JUNC_2</type>
<position>132,-3304</position>
<input>
<ID>N_in1</ID>5480 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1684</ID>
<type>BA_TRI_STATE</type>
<position>210,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1175 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7835</ID>
<type>AE_DFF_LOW</type>
<position>92,-3008</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5298 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1685</ID>
<type>AE_DFF_LOW</type>
<position>223,-246.5</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>1176 </output>
<input>
<ID>clock</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7836</ID>
<type>HA_JUNC_2</type>
<position>151,-3303.5</position>
<input>
<ID>N_in1</ID>5481 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1686</ID>
<type>BA_TRI_STATE</type>
<position>233,-257</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1176 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7837</ID>
<type>BA_TRI_STATE</type>
<position>102,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5298 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1687</ID>
<type>AA_AND2</type>
<position>30.5,-228.5</position>
<input>
<ID>IN_0</ID>3193 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>3160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7838</ID>
<type>HA_JUNC_2</type>
<position>156,-3303.5</position>
<input>
<ID>N_in1</ID>5482 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7839</ID>
<type>AE_DFF_LOW</type>
<position>115,-3008</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5299 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7840</ID>
<type>HA_JUNC_2</type>
<position>174,-3303</position>
<input>
<ID>N_in1</ID>5483 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7841</ID>
<type>BA_TRI_STATE</type>
<position>125,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5299 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7842</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3303</position>
<input>
<ID>N_in1</ID>5484 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7843</ID>
<type>AE_DFF_LOW</type>
<position>138,-3008</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5300 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7844</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3302.5</position>
<input>
<ID>N_in1</ID>5485 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7845</ID>
<type>BA_TRI_STATE</type>
<position>148,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5300 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7846</ID>
<type>HA_JUNC_2</type>
<position>203,-3302.5</position>
<input>
<ID>N_in1</ID>5486 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7847</ID>
<type>AE_DFF_LOW</type>
<position>161,-3008</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5301 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7848</ID>
<type>HA_JUNC_2</type>
<position>203,-3137.5</position>
<input>
<ID>N_in0</ID>5486 </input>
<input>
<ID>N_in1</ID>5514 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7849</ID>
<type>BA_TRI_STATE</type>
<position>171,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5301 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7850</ID>
<type>HA_JUNC_2</type>
<position>224,-3302.5</position>
<input>
<ID>N_in1</ID>5487 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7851</ID>
<type>AE_DFF_LOW</type>
<position>186,-3008</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5302 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7852</ID>
<type>AE_DFF_LOW</type>
<position>67,-3202</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5393 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7853</ID>
<type>BA_TRI_STATE</type>
<position>196,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5302 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7854</ID>
<type>BA_TRI_STATE</type>
<position>77,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5393 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7855</ID>
<type>AE_DFF_LOW</type>
<position>209,-3008</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5303 </output>
<input>
<ID>clock</ID>5304 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7856</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3137.5</position>
<input>
<ID>N_in0</ID>5497 </input>
<input>
<ID>N_in1</ID>5499 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7857</ID>
<type>BA_TRI_STATE</type>
<position>219,-3018.5</position>
<input>
<ID>ENABLE_0</ID>5305 </input>
<input>
<ID>IN_0</ID>5303 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7858</ID>
<type>AE_DFF_LOW</type>
<position>92,-3202</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5394 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7859</ID>
<type>AA_AND2</type>
<position>16.5,-2990</position>
<input>
<ID>IN_0</ID>5383 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7860</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3137.5</position>
<input>
<ID>N_in0</ID>5496 </input>
<input>
<ID>N_in1</ID>5498 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7861</ID>
<type>AA_AND2</type>
<position>28,-2999.5</position>
<input>
<ID>IN_0</ID>5383 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5315 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7862</ID>
<type>BA_TRI_STATE</type>
<position>102,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5394 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7863</ID>
<type>AE_DFF_LOW</type>
<position>44,-2989</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5306 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7864</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3304.5</position>
<input>
<ID>N_in1</ID>5497 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7865</ID>
<type>BA_TRI_STATE</type>
<position>54,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5306 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7866</ID>
<type>AE_DFF_LOW</type>
<position>115,-3202</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5395 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7867</ID>
<type>AE_DFF_LOW</type>
<position>67,-2989</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5307 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7868</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3304.5</position>
<input>
<ID>N_in1</ID>5496 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>7869</ID>
<type>BA_TRI_STATE</type>
<position>77,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5307 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7870</ID>
<type>BA_TRI_STATE</type>
<position>125,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5395 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7871</ID>
<type>AE_DFF_LOW</type>
<position>92,-2989</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5308 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7872</ID>
<type>AE_DFF_LOW</type>
<position>138,-3202</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5396 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7873</ID>
<type>BA_TRI_STATE</type>
<position>102,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5308 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7874</ID>
<type>AA_LABEL</type>
<position>3.5,-3138</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7875</ID>
<type>AE_DFF_LOW</type>
<position>115,-2989</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5309 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7876</ID>
<type>BA_TRI_STATE</type>
<position>148,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5396 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7877</ID>
<type>BA_TRI_STATE</type>
<position>125,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5309 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7878</ID>
<type>AE_DFF_LOW</type>
<position>161,-3202</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5397 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7879</ID>
<type>AE_DFF_LOW</type>
<position>138,-2989</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5310 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7880</ID>
<type>BA_TRI_STATE</type>
<position>171,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5397 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7881</ID>
<type>BA_TRI_STATE</type>
<position>148,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5310 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7882</ID>
<type>AE_DFF_LOW</type>
<position>186,-3202</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5398 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7883</ID>
<type>AE_DFF_LOW</type>
<position>161,-2989</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5311 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7884</ID>
<type>BA_TRI_STATE</type>
<position>196,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5398 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7885</ID>
<type>BA_TRI_STATE</type>
<position>171,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5311 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7886</ID>
<type>AE_DFF_LOW</type>
<position>209,-3202</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5399 </output>
<input>
<ID>clock</ID>5400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7887</ID>
<type>AE_DFF_LOW</type>
<position>186,-2989</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5312 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7888</ID>
<type>BA_TRI_STATE</type>
<position>219,-3212.5</position>
<input>
<ID>ENABLE_0</ID>5401 </input>
<input>
<ID>IN_0</ID>5399 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7889</ID>
<type>BA_TRI_STATE</type>
<position>196,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5312 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7890</ID>
<type>AA_AND2</type>
<position>16.5,-3184.5</position>
<input>
<ID>IN_0</ID>5490 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7891</ID>
<type>AE_DFF_LOW</type>
<position>209,-2989</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5313 </output>
<input>
<ID>clock</ID>5314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7892</ID>
<type>AA_AND2</type>
<position>28,-3194</position>
<input>
<ID>IN_0</ID>5490 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7893</ID>
<type>BA_TRI_STATE</type>
<position>219,-2999.5</position>
<input>
<ID>ENABLE_0</ID>5315 </input>
<input>
<ID>IN_0</ID>5313 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7894</ID>
<type>AE_DFF_LOW</type>
<position>44,-3183.5</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5402 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7895</ID>
<type>AA_AND2</type>
<position>16.5,-2971.5</position>
<input>
<ID>IN_0</ID>5382 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5324 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7896</ID>
<type>BA_TRI_STATE</type>
<position>54,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5402 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7897</ID>
<type>AA_AND2</type>
<position>28,-2981</position>
<input>
<ID>IN_0</ID>5382 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7898</ID>
<type>AE_DFF_LOW</type>
<position>67,-3183.5</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5403 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7899</ID>
<type>AE_DFF_LOW</type>
<position>44,-2970.5</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5316 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7900</ID>
<type>BA_TRI_STATE</type>
<position>77,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5403 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7901</ID>
<type>BA_TRI_STATE</type>
<position>54,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5316 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7902</ID>
<type>AE_DFF_LOW</type>
<position>92,-3183.5</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5404 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7903</ID>
<type>AE_DFF_LOW</type>
<position>67,-2970.5</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5317 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7904</ID>
<type>BA_TRI_STATE</type>
<position>102,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5404 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7905</ID>
<type>BA_TRI_STATE</type>
<position>77,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5317 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7906</ID>
<type>AE_DFF_LOW</type>
<position>115,-3183.5</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5405 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7907</ID>
<type>AE_DFF_LOW</type>
<position>92,-2970.5</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5318 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7908</ID>
<type>BA_TRI_STATE</type>
<position>125,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5405 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7909</ID>
<type>BA_TRI_STATE</type>
<position>102,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5318 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7910</ID>
<type>AE_DFF_LOW</type>
<position>138,-3183.5</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5406 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7911</ID>
<type>AE_DFF_LOW</type>
<position>115,-2970.5</position>
<input>
<ID>IN_0</ID>5372 </input>
<output>
<ID>OUT_0</ID>5319 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7912</ID>
<type>BA_TRI_STATE</type>
<position>148,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5406 </input>
<output>
<ID>OUT_0</ID>5481 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7913</ID>
<type>BA_TRI_STATE</type>
<position>125,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5319 </input>
<output>
<ID>OUT_0</ID>5373 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7914</ID>
<type>AE_DFF_LOW</type>
<position>161,-3183.5</position>
<input>
<ID>IN_0</ID>5482 </input>
<output>
<ID>OUT_0</ID>5407 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7915</ID>
<type>AE_DFF_LOW</type>
<position>138,-2970.5</position>
<input>
<ID>IN_0</ID>5374 </input>
<output>
<ID>OUT_0</ID>5320 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7916</ID>
<type>BA_TRI_STATE</type>
<position>171,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5407 </input>
<output>
<ID>OUT_0</ID>5483 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7917</ID>
<type>BA_TRI_STATE</type>
<position>148,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5320 </input>
<output>
<ID>OUT_0</ID>5375 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7918</ID>
<type>AE_DFF_LOW</type>
<position>186,-3183.5</position>
<input>
<ID>IN_0</ID>5484 </input>
<output>
<ID>OUT_0</ID>5408 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7919</ID>
<type>AE_DFF_LOW</type>
<position>161,-2970.5</position>
<input>
<ID>IN_0</ID>5376 </input>
<output>
<ID>OUT_0</ID>5321 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7920</ID>
<type>BA_TRI_STATE</type>
<position>196,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5408 </input>
<output>
<ID>OUT_0</ID>5485 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7921</ID>
<type>BA_TRI_STATE</type>
<position>171,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5321 </input>
<output>
<ID>OUT_0</ID>5377 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7922</ID>
<type>AE_DFF_LOW</type>
<position>209,-3183.5</position>
<input>
<ID>IN_0</ID>5486 </input>
<output>
<ID>OUT_0</ID>5409 </output>
<input>
<ID>clock</ID>5410 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7923</ID>
<type>AE_DFF_LOW</type>
<position>186,-2970.5</position>
<input>
<ID>IN_0</ID>5378 </input>
<output>
<ID>OUT_0</ID>5322 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7924</ID>
<type>BA_TRI_STATE</type>
<position>219,-3194</position>
<input>
<ID>ENABLE_0</ID>5411 </input>
<input>
<ID>IN_0</ID>5409 </input>
<output>
<ID>OUT_0</ID>5487 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7925</ID>
<type>BA_TRI_STATE</type>
<position>196,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5322 </input>
<output>
<ID>OUT_0</ID>5379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7926</ID>
<type>AA_AND2</type>
<position>16.5,-3165.5</position>
<input>
<ID>IN_0</ID>5489 </input>
<input>
<ID>IN_1</ID>5496 </input>
<output>
<ID>OUT</ID>5420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7927</ID>
<type>AE_DFF_LOW</type>
<position>209,-2970.5</position>
<input>
<ID>IN_0</ID>5380 </input>
<output>
<ID>OUT_0</ID>5323 </output>
<input>
<ID>clock</ID>5324 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7928</ID>
<type>AA_AND2</type>
<position>28,-3175</position>
<input>
<ID>IN_0</ID>5489 </input>
<input>
<ID>IN_1</ID>5497 </input>
<output>
<ID>OUT</ID>5421 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7929</ID>
<type>BA_TRI_STATE</type>
<position>219,-2981</position>
<input>
<ID>ENABLE_0</ID>5325 </input>
<input>
<ID>IN_0</ID>5323 </input>
<output>
<ID>OUT_0</ID>5381 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7930</ID>
<type>AE_DFF_LOW</type>
<position>44,-3164.5</position>
<input>
<ID>IN_0</ID>5472 </input>
<output>
<ID>OUT_0</ID>5412 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7931</ID>
<type>AA_AND2</type>
<position>16.5,-3105.5</position>
<input>
<ID>IN_0</ID>5389 </input>
<input>
<ID>IN_1</ID>5390 </input>
<output>
<ID>OUT</ID>5334 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7932</ID>
<type>BA_TRI_STATE</type>
<position>54,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5412 </input>
<output>
<ID>OUT_0</ID>5473 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7933</ID>
<type>AA_AND2</type>
<position>27.5,-3115</position>
<input>
<ID>IN_0</ID>5389 </input>
<input>
<ID>IN_1</ID>5391 </input>
<output>
<ID>OUT</ID>5335 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7934</ID>
<type>AE_DFF_LOW</type>
<position>67,-3164.5</position>
<input>
<ID>IN_0</ID>5474 </input>
<output>
<ID>OUT_0</ID>5413 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7935</ID>
<type>AE_DFF_LOW</type>
<position>44,-3104.5</position>
<input>
<ID>IN_0</ID>5366 </input>
<output>
<ID>OUT_0</ID>5326 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7936</ID>
<type>BA_TRI_STATE</type>
<position>77,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5413 </input>
<output>
<ID>OUT_0</ID>5475 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7937</ID>
<type>BA_TRI_STATE</type>
<position>54,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5326 </input>
<output>
<ID>OUT_0</ID>5367 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7938</ID>
<type>AE_DFF_LOW</type>
<position>92,-3164.5</position>
<input>
<ID>IN_0</ID>5476 </input>
<output>
<ID>OUT_0</ID>5414 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7939</ID>
<type>AE_DFF_LOW</type>
<position>67,-3104.5</position>
<input>
<ID>IN_0</ID>5368 </input>
<output>
<ID>OUT_0</ID>5327 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7940</ID>
<type>BA_TRI_STATE</type>
<position>102,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5414 </input>
<output>
<ID>OUT_0</ID>5477 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7941</ID>
<type>BA_TRI_STATE</type>
<position>77,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5327 </input>
<output>
<ID>OUT_0</ID>5369 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7942</ID>
<type>AE_DFF_LOW</type>
<position>115,-3164.5</position>
<input>
<ID>IN_0</ID>5478 </input>
<output>
<ID>OUT_0</ID>5415 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7943</ID>
<type>AE_DFF_LOW</type>
<position>92,-3104.5</position>
<input>
<ID>IN_0</ID>5370 </input>
<output>
<ID>OUT_0</ID>5328 </output>
<input>
<ID>clock</ID>5334 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7944</ID>
<type>BA_TRI_STATE</type>
<position>125,-3175</position>
<input>
<ID>ENABLE_0</ID>5421 </input>
<input>
<ID>IN_0</ID>5415 </input>
<output>
<ID>OUT_0</ID>5479 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7945</ID>
<type>BA_TRI_STATE</type>
<position>102,-3115</position>
<input>
<ID>ENABLE_0</ID>5335 </input>
<input>
<ID>IN_0</ID>5328 </input>
<output>
<ID>OUT_0</ID>5371 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7946</ID>
<type>AE_DFF_LOW</type>
<position>138,-3164.5</position>
<input>
<ID>IN_0</ID>5480 </input>
<output>
<ID>OUT_0</ID>5416 </output>
<input>
<ID>clock</ID>5420 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7948</ID>
<type>AA_LABEL</type>
<position>279,-3125.5</position>
<gparam>LABEL_TEXT 9</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7949</ID>
<type>AE_DFF_LOW</type>
<position>115,-3456.5</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5559 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7950</ID>
<type>BA_TRI_STATE</type>
<position>148,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5646 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7951</ID>
<type>BA_TRI_STATE</type>
<position>125,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5559 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7952</ID>
<type>AE_DFF_LOW</type>
<position>161,-3516.5</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5647 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7953</ID>
<type>AE_DFF_LOW</type>
<position>138,-3456.5</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5560 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7954</ID>
<type>BA_TRI_STATE</type>
<position>171,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5647 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7955</ID>
<type>BA_TRI_STATE</type>
<position>148,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5560 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7956</ID>
<type>AE_DFF_LOW</type>
<position>186,-3516.5</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5648 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7957</ID>
<type>AE_DFF_LOW</type>
<position>161,-3456.5</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5561 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7958</ID>
<type>BA_TRI_STATE</type>
<position>196,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5648 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7959</ID>
<type>BA_TRI_STATE</type>
<position>171,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5561 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7960</ID>
<type>AE_DFF_LOW</type>
<position>209,-3516.5</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5649 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7961</ID>
<type>AE_DFF_LOW</type>
<position>186,-3456.5</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5562 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7962</ID>
<type>BA_TRI_STATE</type>
<position>219,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5649 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7963</ID>
<type>BA_TRI_STATE</type>
<position>196,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5562 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7964</ID>
<type>AA_AND2</type>
<position>16.5,-3499</position>
<input>
<ID>IN_0</ID>5718 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5660 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7965</ID>
<type>AE_DFF_LOW</type>
<position>209,-3456.5</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5563 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7966</ID>
<type>AA_AND2</type>
<position>28,-3508.5</position>
<input>
<ID>IN_0</ID>5718 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5661 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7967</ID>
<type>BA_TRI_STATE</type>
<position>219,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5563 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7968</ID>
<type>AE_DFF_LOW</type>
<position>44,-3498</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5652 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7969</ID>
<type>AA_AND2</type>
<position>16.5,-3439</position>
<input>
<ID>IN_0</ID>5618 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5574 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7970</ID>
<type>BA_TRI_STATE</type>
<position>54,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5652 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7971</ID>
<type>AA_AND2</type>
<position>27.5,-3448.5</position>
<input>
<ID>IN_0</ID>5618 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5575 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7972</ID>
<type>AE_DFF_LOW</type>
<position>67,-3498</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5653 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7973</ID>
<type>AE_DFF_LOW</type>
<position>44,-3438</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5566 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7974</ID>
<type>BA_TRI_STATE</type>
<position>77,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5653 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7975</ID>
<type>BA_TRI_STATE</type>
<position>54,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5566 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7976</ID>
<type>AE_DFF_LOW</type>
<position>92,-3498</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5654 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7977</ID>
<type>AE_DFF_LOW</type>
<position>67,-3438</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5567 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7978</ID>
<type>BA_TRI_STATE</type>
<position>102,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5654 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7979</ID>
<type>BA_TRI_STATE</type>
<position>77,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5567 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7980</ID>
<type>AE_DFF_LOW</type>
<position>115,-3498</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5655 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7981</ID>
<type>AE_DFF_LOW</type>
<position>92,-3438</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5568 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7982</ID>
<type>BA_TRI_STATE</type>
<position>125,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5655 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7983</ID>
<type>BA_TRI_STATE</type>
<position>102,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5568 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7984</ID>
<type>AE_DFF_LOW</type>
<position>138,-3498</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5656 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7985</ID>
<type>AE_DFF_LOW</type>
<position>115,-3438</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5569 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7986</ID>
<type>BA_TRI_STATE</type>
<position>148,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5656 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7987</ID>
<type>BA_TRI_STATE</type>
<position>125,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5569 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7988</ID>
<type>AE_DFF_LOW</type>
<position>161,-3498</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5657 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7989</ID>
<type>AE_DFF_LOW</type>
<position>138,-3438</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5570 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7990</ID>
<type>BA_TRI_STATE</type>
<position>171,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5657 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7991</ID>
<type>BA_TRI_STATE</type>
<position>148,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5570 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7992</ID>
<type>AE_DFF_LOW</type>
<position>186,-3498</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5658 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7993</ID>
<type>AE_DFF_LOW</type>
<position>161,-3438</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5571 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7994</ID>
<type>BA_TRI_STATE</type>
<position>196,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5658 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7995</ID>
<type>BA_TRI_STATE</type>
<position>171,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5571 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7996</ID>
<type>AE_DFF_LOW</type>
<position>209,-3498</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5659 </output>
<input>
<ID>clock</ID>5660 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7997</ID>
<type>AE_DFF_LOW</type>
<position>186,-3438</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5572 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7998</ID>
<type>BA_TRI_STATE</type>
<position>219,-3508.5</position>
<input>
<ID>ENABLE_0</ID>5661 </input>
<input>
<ID>IN_0</ID>5659 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7999</ID>
<type>BA_TRI_STATE</type>
<position>196,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5572 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8000</ID>
<type>AA_AND2</type>
<position>16.5,-3633</position>
<input>
<ID>IN_0</ID>5725 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5670 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8001</ID>
<type>AE_DFF_LOW</type>
<position>209,-3438</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5573 </output>
<input>
<ID>clock</ID>5574 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8002</ID>
<type>AA_AND2</type>
<position>27.5,-3642.5</position>
<input>
<ID>IN_0</ID>5725 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5671 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8003</ID>
<type>BA_TRI_STATE</type>
<position>219,-3448.5</position>
<input>
<ID>ENABLE_0</ID>5575 </input>
<input>
<ID>IN_0</ID>5573 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8004</ID>
<type>AE_DFF_LOW</type>
<position>44,-3632</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5662 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8005</ID>
<type>AA_AND2</type>
<position>27.5,-3605</position>
<input>
<ID>IN_0</ID>5723 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5691 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8006</ID>
<type>AA_AND2</type>
<position>16.5,-3420</position>
<input>
<ID>IN_0</ID>5617 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8007</ID>
<type>BA_TRI_STATE</type>
<position>54,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5662 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8008</ID>
<type>AA_AND2</type>
<position>27.5,-3429.5</position>
<input>
<ID>IN_0</ID>5617 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5585 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8009</ID>
<type>AE_DFF_LOW</type>
<position>67,-3632</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5663 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8010</ID>
<type>AE_DFF_LOW</type>
<position>44,-3594.5</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5682 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8011</ID>
<type>AE_DFF_LOW</type>
<position>44,-3419</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5576 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8012</ID>
<type>BA_TRI_STATE</type>
<position>77,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5663 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8013</ID>
<type>BA_TRI_STATE</type>
<position>54,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5576 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8014</ID>
<type>AE_DFF_LOW</type>
<position>92,-3632</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5664 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8015</ID>
<type>BA_TRI_STATE</type>
<position>54,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5682 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8016</ID>
<type>AE_DFF_LOW</type>
<position>67,-3419</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5577 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8017</ID>
<type>BA_TRI_STATE</type>
<position>102,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5664 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8018</ID>
<type>BA_TRI_STATE</type>
<position>77,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5577 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8019</ID>
<type>AE_DFF_LOW</type>
<position>115,-3632</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5665 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8020</ID>
<type>AE_DFF_LOW</type>
<position>67,-3594.5</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5683 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8021</ID>
<type>AE_DFF_LOW</type>
<position>92,-3419</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5578 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8022</ID>
<type>BA_TRI_STATE</type>
<position>125,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5665 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8023</ID>
<type>BA_TRI_STATE</type>
<position>102,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5578 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8024</ID>
<type>AE_DFF_LOW</type>
<position>138,-3632</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5666 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8025</ID>
<type>BA_TRI_STATE</type>
<position>77,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5683 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8026</ID>
<type>AE_DFF_LOW</type>
<position>115,-3419</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5579 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8027</ID>
<type>BA_TRI_STATE</type>
<position>148,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5666 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8028</ID>
<type>BA_TRI_STATE</type>
<position>125,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5579 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8029</ID>
<type>AE_DFF_LOW</type>
<position>161,-3632</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5667 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8030</ID>
<type>AE_DFF_LOW</type>
<position>92,-3594.5</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5684 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8031</ID>
<type>AE_DFF_LOW</type>
<position>138,-3419</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5580 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8032</ID>
<type>BA_TRI_STATE</type>
<position>171,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5667 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8033</ID>
<type>BA_TRI_STATE</type>
<position>148,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5580 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8034</ID>
<type>BA_TRI_STATE</type>
<position>102,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5684 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8035</ID>
<type>AE_DFF_LOW</type>
<position>161,-3419</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5581 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8036</ID>
<type>BA_TRI_STATE</type>
<position>171,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5581 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8037</ID>
<type>AE_DFF_LOW</type>
<position>115,-3594.5</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5685 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8038</ID>
<type>AE_DFF_LOW</type>
<position>186,-3419</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5582 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8039</ID>
<type>BA_TRI_STATE</type>
<position>196,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5582 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8040</ID>
<type>AE_DFF_LOW</type>
<position>209,-3419</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5583 </output>
<input>
<ID>clock</ID>5584 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8041</ID>
<type>BA_TRI_STATE</type>
<position>219,-3429.5</position>
<input>
<ID>ENABLE_0</ID>5585 </input>
<input>
<ID>IN_0</ID>5583 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8042</ID>
<type>AA_AND2</type>
<position>16.5,-3401.5</position>
<input>
<ID>IN_0</ID>5616 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5594 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8043</ID>
<type>AA_AND2</type>
<position>27.5,-3411</position>
<input>
<ID>IN_0</ID>5616 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8044</ID>
<type>AE_DFF_LOW</type>
<position>44,-3400.5</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5586 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8045</ID>
<type>BA_TRI_STATE</type>
<position>54,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5586 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8046</ID>
<type>AE_DFF_LOW</type>
<position>67,-3400.5</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5587 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8047</ID>
<type>BA_TRI_STATE</type>
<position>77,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5587 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8048</ID>
<type>AE_DFF_LOW</type>
<position>92,-3400.5</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5588 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8049</ID>
<type>BA_TRI_STATE</type>
<position>102,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5588 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8050</ID>
<type>AE_DFF_LOW</type>
<position>115,-3400.5</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5589 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8051</ID>
<type>BA_TRI_STATE</type>
<position>125,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5589 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8052</ID>
<type>AE_DFF_LOW</type>
<position>138,-3400.5</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5590 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8053</ID>
<type>BA_TRI_STATE</type>
<position>148,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5590 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8054</ID>
<type>AE_DFF_LOW</type>
<position>161,-3400.5</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5591 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8055</ID>
<type>BA_TRI_STATE</type>
<position>171,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5591 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8056</ID>
<type>AE_DFF_LOW</type>
<position>186,-3400.5</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5592 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8057</ID>
<type>BA_TRI_STATE</type>
<position>196,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5592 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8058</ID>
<type>AE_DFF_LOW</type>
<position>209,-3400.5</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5593 </output>
<input>
<ID>clock</ID>5594 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8059</ID>
<type>BA_TRI_STATE</type>
<position>219,-3411</position>
<input>
<ID>ENABLE_0</ID>5595 </input>
<input>
<ID>IN_0</ID>5593 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8060</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3314</position>
<input>
<ID>N_in0</ID>5596 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8061</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3313.5</position>
<input>
<ID>N_in0</ID>5597 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8062</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3314</position>
<input>
<ID>N_in0</ID>5598 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8063</ID>
<type>HA_JUNC_2</type>
<position>81,-3313.5</position>
<input>
<ID>N_in0</ID>5599 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8064</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3313.5</position>
<input>
<ID>N_in0</ID>5600 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8065</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3314</position>
<input>
<ID>N_in0</ID>5601 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8066</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3313.5</position>
<input>
<ID>N_in0</ID>5602 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8067</ID>
<type>HA_JUNC_2</type>
<position>128,-3313.5</position>
<input>
<ID>N_in0</ID>5603 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8068</ID>
<type>HA_JUNC_2</type>
<position>132,-3313.5</position>
<input>
<ID>N_in0</ID>5604 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8069</ID>
<type>HA_JUNC_2</type>
<position>151,-3313.5</position>
<input>
<ID>N_in0</ID>5605 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8070</ID>
<type>HA_JUNC_2</type>
<position>156,-3313.5</position>
<input>
<ID>N_in0</ID>5606 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8071</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3313.5</position>
<input>
<ID>N_in0</ID>5608 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8072</ID>
<type>HA_JUNC_2</type>
<position>174,-3313.5</position>
<input>
<ID>N_in0</ID>5607 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8073</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3314</position>
<input>
<ID>N_in0</ID>5609 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8074</ID>
<type>HA_JUNC_2</type>
<position>224,-3315</position>
<input>
<ID>N_in0</ID>5611 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8075</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3481</position>
<input>
<ID>N_in0</ID>5730 </input>
<input>
<ID>N_in1</ID>5596 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8076</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3480.5</position>
<input>
<ID>N_in0</ID>5731 </input>
<input>
<ID>N_in1</ID>5597 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8077</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3480.5</position>
<input>
<ID>N_in0</ID>5732 </input>
<input>
<ID>N_in1</ID>5598 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8078</ID>
<type>HA_JUNC_2</type>
<position>81,-3480.5</position>
<input>
<ID>N_in0</ID>5733 </input>
<input>
<ID>N_in1</ID>5599 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8079</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3480.5</position>
<input>
<ID>N_in0</ID>5734 </input>
<input>
<ID>N_in1</ID>5600 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8080</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3480.5</position>
<input>
<ID>N_in0</ID>5735 </input>
<input>
<ID>N_in1</ID>5601 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8081</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3480.5</position>
<input>
<ID>N_in0</ID>5736 </input>
<input>
<ID>N_in1</ID>5602 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8082</ID>
<type>HA_JUNC_2</type>
<position>128,-3480.5</position>
<input>
<ID>N_in0</ID>5737 </input>
<input>
<ID>N_in1</ID>5603 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8083</ID>
<type>HA_JUNC_2</type>
<position>132,-3480.5</position>
<input>
<ID>N_in0</ID>5738 </input>
<input>
<ID>N_in1</ID>5604 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8084</ID>
<type>HA_JUNC_2</type>
<position>151,-3480</position>
<input>
<ID>N_in0</ID>5739 </input>
<input>
<ID>N_in1</ID>5605 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8085</ID>
<type>HA_JUNC_2</type>
<position>156,-3480</position>
<input>
<ID>N_in0</ID>5740 </input>
<input>
<ID>N_in1</ID>5606 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8086</ID>
<type>HA_JUNC_2</type>
<position>174,-3479.5</position>
<input>
<ID>N_in0</ID>5741 </input>
<input>
<ID>N_in1</ID>5607 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8087</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3479.5</position>
<input>
<ID>N_in0</ID>5742 </input>
<input>
<ID>N_in1</ID>5608 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8088</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3479</position>
<input>
<ID>N_in0</ID>5743 </input>
<input>
<ID>N_in1</ID>5609 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8089</ID>
<type>HA_JUNC_2</type>
<position>203,-3479</position>
<input>
<ID>N_in0</ID>5744 </input>
<input>
<ID>N_in1</ID>5610 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8090</ID>
<type>HA_JUNC_2</type>
<position>203,-3314</position>
<input>
<ID>N_in0</ID>5610 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8091</ID>
<type>HA_JUNC_2</type>
<position>224,-3479</position>
<input>
<ID>N_in0</ID>5745 </input>
<input>
<ID>N_in1</ID>5611 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8092</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3314</position>
<input>
<ID>N_in0</ID>5621 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8093</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3314</position>
<input>
<ID>N_in0</ID>5620 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8094</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3481</position>
<input>
<ID>N_in0</ID>5729 </input>
<input>
<ID>N_in1</ID>5621 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8095</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3481</position>
<input>
<ID>N_in0</ID>5728 </input>
<input>
<ID>N_in1</ID>5620 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8096</ID>
<type>AA_LABEL</type>
<position>3.5,-3314.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8097</ID>
<type>BI_DECODER_4x16</type>
<position>-136,-3481.5</position>
<output>
<ID>OUT_0</ID>5725 </output>
<output>
<ID>OUT_1</ID>5724 </output>
<output>
<ID>OUT_10</ID>5617 </output>
<output>
<ID>OUT_11</ID>5616 </output>
<output>
<ID>OUT_12</ID>5615 </output>
<output>
<ID>OUT_13</ID>5614 </output>
<output>
<ID>OUT_14</ID>5613 </output>
<output>
<ID>OUT_15</ID>5612 </output>
<output>
<ID>OUT_2</ID>5723 </output>
<output>
<ID>OUT_3</ID>5722 </output>
<output>
<ID>OUT_4</ID>5721 </output>
<output>
<ID>OUT_5</ID>5720 </output>
<output>
<ID>OUT_6</ID>5719 </output>
<output>
<ID>OUT_7</ID>5718 </output>
<output>
<ID>OUT_8</ID>5619 </output>
<output>
<ID>OUT_9</ID>5618 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8098</ID>
<type>AE_DFF_LOW</type>
<position>186,-3632</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5668 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8099</ID>
<type>BA_TRI_STATE</type>
<position>196,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5668 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8100</ID>
<type>AE_DFF_LOW</type>
<position>209,-3632</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5669 </output>
<input>
<ID>clock</ID>5670 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8101</ID>
<type>BA_TRI_STATE</type>
<position>219,-3642.5</position>
<input>
<ID>ENABLE_0</ID>5671 </input>
<input>
<ID>IN_0</ID>5669 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8102</ID>
<type>AA_AND2</type>
<position>16.5,-3614.5</position>
<input>
<ID>IN_0</ID>5724 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5680 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8103</ID>
<type>AA_AND2</type>
<position>27.5,-3624</position>
<input>
<ID>IN_0</ID>5724 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5681 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8104</ID>
<type>AE_DFF_LOW</type>
<position>44,-3613.5</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5672 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8105</ID>
<type>BA_TRI_STATE</type>
<position>54,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5672 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1955</ID>
<type>AA_AND2</type>
<position>41.5,-238</position>
<input>
<ID>IN_0</ID>3193 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>3161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8106</ID>
<type>AE_DFF_LOW</type>
<position>67,-3613.5</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5673 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8107</ID>
<type>BA_TRI_STATE</type>
<position>77,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5673 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1957</ID>
<type>AE_DFF_LOW</type>
<position>58,-227.5</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1644 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8108</ID>
<type>AE_DFF_LOW</type>
<position>92,-3613.5</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5674 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8109</ID>
<type>BA_TRI_STATE</type>
<position>102,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5674 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1959</ID>
<type>BA_TRI_STATE</type>
<position>68,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>1644 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8110</ID>
<type>AE_DFF_LOW</type>
<position>115,-3613.5</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5675 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8111</ID>
<type>BA_TRI_STATE</type>
<position>125,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5675 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1961</ID>
<type>AE_DFF_LOW</type>
<position>81,-227.5</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1645 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8112</ID>
<type>AE_DFF_LOW</type>
<position>138,-3613.5</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5676 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8113</ID>
<type>BA_TRI_STATE</type>
<position>148,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5676 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1963</ID>
<type>BA_TRI_STATE</type>
<position>91,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>1645 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8114</ID>
<type>AE_DFF_LOW</type>
<position>161,-3613.5</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5677 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8115</ID>
<type>BA_TRI_STATE</type>
<position>171,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5677 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1965</ID>
<type>AE_DFF_LOW</type>
<position>106,-227.5</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1646 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8116</ID>
<type>AE_DFF_LOW</type>
<position>186,-3613.5</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5678 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8117</ID>
<type>BA_TRI_STATE</type>
<position>196,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5678 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1967</ID>
<type>BA_TRI_STATE</type>
<position>116,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>1646 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8118</ID>
<type>AE_DFF_LOW</type>
<position>209,-3613.5</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5679 </output>
<input>
<ID>clock</ID>5680 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8119</ID>
<type>BA_TRI_STATE</type>
<position>219,-3624</position>
<input>
<ID>ENABLE_0</ID>5681 </input>
<input>
<ID>IN_0</ID>5679 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1969</ID>
<type>AE_DFF_LOW</type>
<position>129,-227.5</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1647 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8120</ID>
<type>AA_AND2</type>
<position>16.5,-3595.5</position>
<input>
<ID>IN_0</ID>5723 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5690 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8121</ID>
<type>BA_TRI_STATE</type>
<position>125,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5685 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8122</ID>
<type>AE_DFF_LOW</type>
<position>138,-3594.5</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5686 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8123</ID>
<type>BA_TRI_STATE</type>
<position>148,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5686 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8124</ID>
<type>AE_DFF_LOW</type>
<position>161,-3594.5</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5687 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8125</ID>
<type>BA_TRI_STATE</type>
<position>171,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5687 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8126</ID>
<type>AE_DFF_LOW</type>
<position>186,-3594.5</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5688 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8127</ID>
<type>BA_TRI_STATE</type>
<position>196,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5688 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8128</ID>
<type>AA_AND2</type>
<position>16.5,-3379.5</position>
<input>
<ID>IN_0</ID>5615 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8129</ID>
<type>AE_DFF_LOW</type>
<position>209,-3594.5</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5689 </output>
<input>
<ID>clock</ID>5690 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8130</ID>
<type>BA_TRI_STATE</type>
<position>219,-3605</position>
<input>
<ID>ENABLE_0</ID>5691 </input>
<input>
<ID>IN_0</ID>5689 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8131</ID>
<type>AA_AND2</type>
<position>16.5,-3577</position>
<input>
<ID>IN_0</ID>5722 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5700 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8132</ID>
<type>AA_AND2</type>
<position>27.5,-3586.5</position>
<input>
<ID>IN_0</ID>5722 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5701 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8133</ID>
<type>AA_AND2</type>
<position>28,-3389</position>
<input>
<ID>IN_0</ID>5615 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5525 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8134</ID>
<type>AE_DFF_LOW</type>
<position>44,-3576</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5692 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8135</ID>
<type>BA_TRI_STATE</type>
<position>54,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5692 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8136</ID>
<type>AE_DFF_LOW</type>
<position>67,-3576</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5693 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8137</ID>
<type>BA_TRI_STATE</type>
<position>77,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5693 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8138</ID>
<type>AE_DFF_LOW</type>
<position>44,-3378.5</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5516 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8139</ID>
<type>AE_DFF_LOW</type>
<position>92,-3576</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5694 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8140</ID>
<type>BA_TRI_STATE</type>
<position>102,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5694 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8141</ID>
<type>AE_DFF_LOW</type>
<position>115,-3576</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5695 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8142</ID>
<type>BA_TRI_STATE</type>
<position>125,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5695 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8143</ID>
<type>AE_DFF_LOW</type>
<position>138,-3576</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5696 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8144</ID>
<type>BA_TRI_STATE</type>
<position>54,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5516 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8145</ID>
<type>BA_TRI_STATE</type>
<position>148,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5696 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8146</ID>
<type>AE_DFF_LOW</type>
<position>161,-3576</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5697 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8147</ID>
<type>BA_TRI_STATE</type>
<position>171,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5697 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8148</ID>
<type>AE_DFF_LOW</type>
<position>186,-3576</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5698 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8149</ID>
<type>BA_TRI_STATE</type>
<position>196,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5698 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8150</ID>
<type>AE_DFF_LOW</type>
<position>209,-3576</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5699 </output>
<input>
<ID>clock</ID>5700 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8151</ID>
<type>BA_TRI_STATE</type>
<position>219,-3586.5</position>
<input>
<ID>ENABLE_0</ID>5701 </input>
<input>
<ID>IN_0</ID>5699 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8152</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3489.5</position>
<input>
<ID>N_in0</ID>5702 </input>
<input>
<ID>N_in1</ID>5730 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8153</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3489</position>
<input>
<ID>N_in0</ID>5703 </input>
<input>
<ID>N_in1</ID>5731 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8154</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3489.5</position>
<input>
<ID>N_in0</ID>5704 </input>
<input>
<ID>N_in1</ID>5732 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8155</ID>
<type>HA_JUNC_2</type>
<position>81,-3489</position>
<input>
<ID>N_in0</ID>5705 </input>
<input>
<ID>N_in1</ID>5733 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8156</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3489</position>
<input>
<ID>N_in0</ID>5706 </input>
<input>
<ID>N_in1</ID>5734 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8157</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3489.5</position>
<input>
<ID>N_in0</ID>5707 </input>
<input>
<ID>N_in1</ID>5735 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8158</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3489</position>
<input>
<ID>N_in0</ID>5708 </input>
<input>
<ID>N_in1</ID>5736 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8159</ID>
<type>HA_JUNC_2</type>
<position>128,-3489</position>
<input>
<ID>N_in0</ID>5709 </input>
<input>
<ID>N_in1</ID>5737 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8160</ID>
<type>AE_DFF_LOW</type>
<position>67,-3378.5</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5517 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8161</ID>
<type>HA_JUNC_2</type>
<position>132,-3489</position>
<input>
<ID>N_in0</ID>5710 </input>
<input>
<ID>N_in1</ID>5738 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8162</ID>
<type>BA_TRI_STATE</type>
<position>77,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5517 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8163</ID>
<type>HA_JUNC_2</type>
<position>151,-3489</position>
<input>
<ID>N_in0</ID>5711 </input>
<input>
<ID>N_in1</ID>5739 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8164</ID>
<type>AE_DFF_LOW</type>
<position>92,-3378.5</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5518 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8165</ID>
<type>HA_JUNC_2</type>
<position>156,-3489</position>
<input>
<ID>N_in0</ID>5712 </input>
<input>
<ID>N_in1</ID>5740 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8166</ID>
<type>BA_TRI_STATE</type>
<position>102,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5518 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8167</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3489</position>
<input>
<ID>N_in0</ID>5714 </input>
<input>
<ID>N_in1</ID>5742 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8168</ID>
<type>AE_DFF_LOW</type>
<position>115,-3378.5</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5519 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8169</ID>
<type>HA_JUNC_2</type>
<position>174,-3489</position>
<input>
<ID>N_in0</ID>5713 </input>
<input>
<ID>N_in1</ID>5741 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8170</ID>
<type>BA_TRI_STATE</type>
<position>125,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5519 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8171</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3489.5</position>
<input>
<ID>N_in0</ID>5715 </input>
<input>
<ID>N_in1</ID>5743 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8172</ID>
<type>AE_DFF_LOW</type>
<position>138,-3378.5</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5520 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8173</ID>
<type>HA_JUNC_2</type>
<position>224,-3490.5</position>
<input>
<ID>N_in0</ID>5717 </input>
<input>
<ID>N_in1</ID>5745 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8174</ID>
<type>BA_TRI_STATE</type>
<position>148,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5520 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8175</ID>
<type>AA_AND2</type>
<position>16.5,-3555</position>
<input>
<ID>IN_0</ID>5721 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5630 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8176</ID>
<type>AE_DFF_LOW</type>
<position>161,-3378.5</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5521 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8177</ID>
<type>AA_AND2</type>
<position>28,-3564.5</position>
<input>
<ID>IN_0</ID>5721 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5631 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8178</ID>
<type>BA_TRI_STATE</type>
<position>171,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5521 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8179</ID>
<type>HA_JUNC_2</type>
<position>35.5,-3656.5</position>
<input>
<ID>N_in1</ID>5702 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8180</ID>
<type>AE_DFF_LOW</type>
<position>186,-3378.5</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5522 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8181</ID>
<type>AE_DFF_LOW</type>
<position>44,-3554</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5622 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8182</ID>
<type>BA_TRI_STATE</type>
<position>196,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5522 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8183</ID>
<type>HA_JUNC_2</type>
<position>58.5,-3656</position>
<input>
<ID>N_in1</ID>5703 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8184</ID>
<type>AE_DFF_LOW</type>
<position>209,-3378.5</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5523 </output>
<input>
<ID>clock</ID>5524 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8185</ID>
<type>HA_JUNC_2</type>
<position>61.5,-3656</position>
<input>
<ID>N_in1</ID>5704 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8186</ID>
<type>BA_TRI_STATE</type>
<position>219,-3389</position>
<input>
<ID>ENABLE_0</ID>5525 </input>
<input>
<ID>IN_0</ID>5523 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8187</ID>
<type>HA_JUNC_2</type>
<position>81,-3656</position>
<input>
<ID>N_in1</ID>5705 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8188</ID>
<type>AA_AND2</type>
<position>16.5,-3361</position>
<input>
<ID>IN_0</ID>5614 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5534 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8189</ID>
<type>HA_JUNC_2</type>
<position>84.5,-3656</position>
<input>
<ID>N_in1</ID>5706 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8190</ID>
<type>AA_AND2</type>
<position>28,-3370.5</position>
<input>
<ID>IN_0</ID>5614 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5535 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8191</ID>
<type>HA_JUNC_2</type>
<position>105.5,-3656</position>
<input>
<ID>N_in1</ID>5707 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8192</ID>
<type>AE_DFF_LOW</type>
<position>44,-3360</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5526 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8193</ID>
<type>BA_TRI_STATE</type>
<position>54,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5622 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8194</ID>
<type>BA_TRI_STATE</type>
<position>54,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5526 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8195</ID>
<type>HA_JUNC_2</type>
<position>109.5,-3656</position>
<input>
<ID>N_in1</ID>5708 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8196</ID>
<type>AE_DFF_LOW</type>
<position>67,-3360</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5527 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8197</ID>
<type>HA_JUNC_2</type>
<position>128,-3656</position>
<input>
<ID>N_in1</ID>5709 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8198</ID>
<type>BA_TRI_STATE</type>
<position>77,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5527 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8199</ID>
<type>HA_JUNC_2</type>
<position>132,-3656</position>
<input>
<ID>N_in1</ID>5710 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8200</ID>
<type>AE_DFF_LOW</type>
<position>92,-3360</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5528 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8201</ID>
<type>HA_JUNC_2</type>
<position>151,-3655.5</position>
<input>
<ID>N_in1</ID>5711 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8202</ID>
<type>BA_TRI_STATE</type>
<position>102,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5528 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8203</ID>
<type>HA_JUNC_2</type>
<position>156,-3655.5</position>
<input>
<ID>N_in1</ID>5712 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8204</ID>
<type>AE_DFF_LOW</type>
<position>115,-3360</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5529 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8205</ID>
<type>HA_JUNC_2</type>
<position>174,-3655</position>
<input>
<ID>N_in1</ID>5713 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8206</ID>
<type>BA_TRI_STATE</type>
<position>125,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5529 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8207</ID>
<type>HA_JUNC_2</type>
<position>178.5,-3655</position>
<input>
<ID>N_in1</ID>5714 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8208</ID>
<type>AE_DFF_LOW</type>
<position>138,-3360</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5530 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8209</ID>
<type>HA_JUNC_2</type>
<position>199.5,-3654.5</position>
<input>
<ID>N_in1</ID>5715 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8210</ID>
<type>BA_TRI_STATE</type>
<position>148,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5530 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8211</ID>
<type>HA_JUNC_2</type>
<position>203,-3654.5</position>
<input>
<ID>N_in1</ID>5716 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8212</ID>
<type>AE_DFF_LOW</type>
<position>161,-3360</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5531 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8213</ID>
<type>HA_JUNC_2</type>
<position>203,-3489.5</position>
<input>
<ID>N_in0</ID>5716 </input>
<input>
<ID>N_in1</ID>5744 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8214</ID>
<type>BA_TRI_STATE</type>
<position>171,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5531 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8215</ID>
<type>HA_JUNC_2</type>
<position>224,-3654.5</position>
<input>
<ID>N_in1</ID>5717 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8216</ID>
<type>AE_DFF_LOW</type>
<position>186,-3360</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5532 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8217</ID>
<type>AE_DFF_LOW</type>
<position>67,-3554</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5623 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8218</ID>
<type>BA_TRI_STATE</type>
<position>196,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5532 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8219</ID>
<type>BA_TRI_STATE</type>
<position>77,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5623 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8220</ID>
<type>AE_DFF_LOW</type>
<position>209,-3360</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5533 </output>
<input>
<ID>clock</ID>5534 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8221</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3489.5</position>
<input>
<ID>N_in0</ID>5727 </input>
<input>
<ID>N_in1</ID>5729 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8222</ID>
<type>BA_TRI_STATE</type>
<position>219,-3370.5</position>
<input>
<ID>ENABLE_0</ID>5535 </input>
<input>
<ID>IN_0</ID>5533 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8223</ID>
<type>AE_DFF_LOW</type>
<position>92,-3554</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5624 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8224</ID>
<type>AA_AND2</type>
<position>16.5,-3342</position>
<input>
<ID>IN_0</ID>5613 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5544 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8225</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3489.5</position>
<input>
<ID>N_in0</ID>5726 </input>
<input>
<ID>N_in1</ID>5728 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8226</ID>
<type>AA_AND2</type>
<position>28,-3351.5</position>
<input>
<ID>IN_0</ID>5613 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5545 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8227</ID>
<type>BA_TRI_STATE</type>
<position>102,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5624 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8228</ID>
<type>AE_DFF_LOW</type>
<position>44,-3341</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5536 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8229</ID>
<type>HA_JUNC_2</type>
<position>22.5,-3656.5</position>
<input>
<ID>N_in1</ID>5727 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8230</ID>
<type>BA_TRI_STATE</type>
<position>54,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5536 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8231</ID>
<type>AE_DFF_LOW</type>
<position>115,-3554</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5625 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8232</ID>
<type>AE_DFF_LOW</type>
<position>67,-3341</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5537 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8233</ID>
<type>HA_JUNC_2</type>
<position>12.5,-3656.5</position>
<input>
<ID>N_in1</ID>5726 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>8234</ID>
<type>BA_TRI_STATE</type>
<position>77,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5537 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8235</ID>
<type>BA_TRI_STATE</type>
<position>125,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5625 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8236</ID>
<type>AE_DFF_LOW</type>
<position>92,-3341</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5538 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8237</ID>
<type>AE_DFF_LOW</type>
<position>138,-3554</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5626 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8238</ID>
<type>BA_TRI_STATE</type>
<position>102,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5538 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8239</ID>
<type>AA_LABEL</type>
<position>3.5,-3490</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8240</ID>
<type>AE_DFF_LOW</type>
<position>115,-3341</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5539 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8241</ID>
<type>BA_TRI_STATE</type>
<position>148,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5626 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8242</ID>
<type>BA_TRI_STATE</type>
<position>125,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5539 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8243</ID>
<type>AE_DFF_LOW</type>
<position>161,-3554</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5627 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8244</ID>
<type>AE_DFF_LOW</type>
<position>138,-3341</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5540 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8245</ID>
<type>BA_TRI_STATE</type>
<position>171,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5627 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8246</ID>
<type>BA_TRI_STATE</type>
<position>148,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5540 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8247</ID>
<type>AE_DFF_LOW</type>
<position>186,-3554</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5628 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8248</ID>
<type>AE_DFF_LOW</type>
<position>161,-3341</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5541 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8249</ID>
<type>BA_TRI_STATE</type>
<position>196,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5628 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8250</ID>
<type>BA_TRI_STATE</type>
<position>171,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5541 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8251</ID>
<type>AE_DFF_LOW</type>
<position>209,-3554</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5629 </output>
<input>
<ID>clock</ID>5630 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8252</ID>
<type>AE_DFF_LOW</type>
<position>186,-3341</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5542 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8253</ID>
<type>BA_TRI_STATE</type>
<position>219,-3564.5</position>
<input>
<ID>ENABLE_0</ID>5631 </input>
<input>
<ID>IN_0</ID>5629 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8254</ID>
<type>BA_TRI_STATE</type>
<position>196,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5542 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8255</ID>
<type>AA_AND2</type>
<position>16.5,-3536.5</position>
<input>
<ID>IN_0</ID>5720 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5640 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8256</ID>
<type>AE_DFF_LOW</type>
<position>209,-3341</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5543 </output>
<input>
<ID>clock</ID>5544 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8257</ID>
<type>AA_AND2</type>
<position>28,-3546</position>
<input>
<ID>IN_0</ID>5720 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8258</ID>
<type>BA_TRI_STATE</type>
<position>219,-3351.5</position>
<input>
<ID>ENABLE_0</ID>5545 </input>
<input>
<ID>IN_0</ID>5543 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8259</ID>
<type>AE_DFF_LOW</type>
<position>44,-3535.5</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5632 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8260</ID>
<type>AA_AND2</type>
<position>16.5,-3323.5</position>
<input>
<ID>IN_0</ID>5612 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5554 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8261</ID>
<type>BA_TRI_STATE</type>
<position>54,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5632 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8262</ID>
<type>AA_AND2</type>
<position>28,-3333</position>
<input>
<ID>IN_0</ID>5612 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8263</ID>
<type>AE_DFF_LOW</type>
<position>67,-3535.5</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5633 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8264</ID>
<type>AE_DFF_LOW</type>
<position>44,-3322.5</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5546 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8265</ID>
<type>BA_TRI_STATE</type>
<position>77,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5633 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8266</ID>
<type>BA_TRI_STATE</type>
<position>54,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5546 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8267</ID>
<type>AE_DFF_LOW</type>
<position>92,-3535.5</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5634 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8268</ID>
<type>AE_DFF_LOW</type>
<position>67,-3322.5</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5547 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8269</ID>
<type>BA_TRI_STATE</type>
<position>102,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5634 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8270</ID>
<type>BA_TRI_STATE</type>
<position>77,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5547 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8271</ID>
<type>AE_DFF_LOW</type>
<position>115,-3535.5</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5635 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8272</ID>
<type>AE_DFF_LOW</type>
<position>92,-3322.5</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5548 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8273</ID>
<type>BA_TRI_STATE</type>
<position>125,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5635 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8274</ID>
<type>BA_TRI_STATE</type>
<position>102,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5548 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8275</ID>
<type>AE_DFF_LOW</type>
<position>138,-3535.5</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5636 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8276</ID>
<type>AE_DFF_LOW</type>
<position>115,-3322.5</position>
<input>
<ID>IN_0</ID>5602 </input>
<output>
<ID>OUT_0</ID>5549 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8277</ID>
<type>BA_TRI_STATE</type>
<position>148,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5636 </input>
<output>
<ID>OUT_0</ID>5711 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8278</ID>
<type>BA_TRI_STATE</type>
<position>125,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5549 </input>
<output>
<ID>OUT_0</ID>5603 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8279</ID>
<type>AE_DFF_LOW</type>
<position>161,-3535.5</position>
<input>
<ID>IN_0</ID>5712 </input>
<output>
<ID>OUT_0</ID>5637 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8280</ID>
<type>AE_DFF_LOW</type>
<position>138,-3322.5</position>
<input>
<ID>IN_0</ID>5604 </input>
<output>
<ID>OUT_0</ID>5550 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8281</ID>
<type>BA_TRI_STATE</type>
<position>171,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5637 </input>
<output>
<ID>OUT_0</ID>5713 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8282</ID>
<type>BA_TRI_STATE</type>
<position>148,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5550 </input>
<output>
<ID>OUT_0</ID>5605 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8283</ID>
<type>AE_DFF_LOW</type>
<position>186,-3535.5</position>
<input>
<ID>IN_0</ID>5714 </input>
<output>
<ID>OUT_0</ID>5638 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8284</ID>
<type>AE_DFF_LOW</type>
<position>161,-3322.5</position>
<input>
<ID>IN_0</ID>5606 </input>
<output>
<ID>OUT_0</ID>5551 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8285</ID>
<type>BA_TRI_STATE</type>
<position>196,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5638 </input>
<output>
<ID>OUT_0</ID>5715 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8286</ID>
<type>BA_TRI_STATE</type>
<position>171,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5551 </input>
<output>
<ID>OUT_0</ID>5607 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8287</ID>
<type>AE_DFF_LOW</type>
<position>209,-3535.5</position>
<input>
<ID>IN_0</ID>5716 </input>
<output>
<ID>OUT_0</ID>5639 </output>
<input>
<ID>clock</ID>5640 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8288</ID>
<type>AE_DFF_LOW</type>
<position>186,-3322.5</position>
<input>
<ID>IN_0</ID>5608 </input>
<output>
<ID>OUT_0</ID>5552 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8289</ID>
<type>BA_TRI_STATE</type>
<position>219,-3546</position>
<input>
<ID>ENABLE_0</ID>5641 </input>
<input>
<ID>IN_0</ID>5639 </input>
<output>
<ID>OUT_0</ID>5717 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8290</ID>
<type>BA_TRI_STATE</type>
<position>196,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5552 </input>
<output>
<ID>OUT_0</ID>5609 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8291</ID>
<type>AA_AND2</type>
<position>16.5,-3517.5</position>
<input>
<ID>IN_0</ID>5719 </input>
<input>
<ID>IN_1</ID>5726 </input>
<output>
<ID>OUT</ID>5650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8292</ID>
<type>AE_DFF_LOW</type>
<position>209,-3322.5</position>
<input>
<ID>IN_0</ID>5610 </input>
<output>
<ID>OUT_0</ID>5553 </output>
<input>
<ID>clock</ID>5554 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8293</ID>
<type>AA_AND2</type>
<position>28,-3527</position>
<input>
<ID>IN_0</ID>5719 </input>
<input>
<ID>IN_1</ID>5727 </input>
<output>
<ID>OUT</ID>5651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8294</ID>
<type>BA_TRI_STATE</type>
<position>219,-3333</position>
<input>
<ID>ENABLE_0</ID>5555 </input>
<input>
<ID>IN_0</ID>5553 </input>
<output>
<ID>OUT_0</ID>5611 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8295</ID>
<type>AE_DFF_LOW</type>
<position>44,-3516.5</position>
<input>
<ID>IN_0</ID>5702 </input>
<output>
<ID>OUT_0</ID>5642 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8296</ID>
<type>AA_AND2</type>
<position>16.5,-3457.5</position>
<input>
<ID>IN_0</ID>5619 </input>
<input>
<ID>IN_1</ID>5620 </input>
<output>
<ID>OUT</ID>5564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8297</ID>
<type>BA_TRI_STATE</type>
<position>54,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5642 </input>
<output>
<ID>OUT_0</ID>5703 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8298</ID>
<type>AA_AND2</type>
<position>27.5,-3467</position>
<input>
<ID>IN_0</ID>5619 </input>
<input>
<ID>IN_1</ID>5621 </input>
<output>
<ID>OUT</ID>5565 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8299</ID>
<type>AE_DFF_LOW</type>
<position>67,-3516.5</position>
<input>
<ID>IN_0</ID>5704 </input>
<output>
<ID>OUT_0</ID>5643 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8300</ID>
<type>AE_DFF_LOW</type>
<position>44,-3456.5</position>
<input>
<ID>IN_0</ID>5596 </input>
<output>
<ID>OUT_0</ID>5556 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8301</ID>
<type>BA_TRI_STATE</type>
<position>77,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5643 </input>
<output>
<ID>OUT_0</ID>5705 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8302</ID>
<type>BA_TRI_STATE</type>
<position>54,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5556 </input>
<output>
<ID>OUT_0</ID>5597 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8303</ID>
<type>AE_DFF_LOW</type>
<position>92,-3516.5</position>
<input>
<ID>IN_0</ID>5706 </input>
<output>
<ID>OUT_0</ID>5644 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8304</ID>
<type>AE_DFF_LOW</type>
<position>67,-3456.5</position>
<input>
<ID>IN_0</ID>5598 </input>
<output>
<ID>OUT_0</ID>5557 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8305</ID>
<type>BA_TRI_STATE</type>
<position>102,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5644 </input>
<output>
<ID>OUT_0</ID>5707 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8306</ID>
<type>BA_TRI_STATE</type>
<position>77,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5557 </input>
<output>
<ID>OUT_0</ID>5599 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8307</ID>
<type>AE_DFF_LOW</type>
<position>115,-3516.5</position>
<input>
<ID>IN_0</ID>5708 </input>
<output>
<ID>OUT_0</ID>5645 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8308</ID>
<type>AE_DFF_LOW</type>
<position>92,-3456.5</position>
<input>
<ID>IN_0</ID>5600 </input>
<output>
<ID>OUT_0</ID>5558 </output>
<input>
<ID>clock</ID>5564 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8309</ID>
<type>BA_TRI_STATE</type>
<position>125,-3527</position>
<input>
<ID>ENABLE_0</ID>5651 </input>
<input>
<ID>IN_0</ID>5645 </input>
<output>
<ID>OUT_0</ID>5709 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8310</ID>
<type>BA_TRI_STATE</type>
<position>102,-3467</position>
<input>
<ID>ENABLE_0</ID>5565 </input>
<input>
<ID>IN_0</ID>5558 </input>
<output>
<ID>OUT_0</ID>5601 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8311</ID>
<type>AE_DFF_LOW</type>
<position>138,-3516.5</position>
<input>
<ID>IN_0</ID>5710 </input>
<output>
<ID>OUT_0</ID>5646 </output>
<input>
<ID>clock</ID>5650 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8313</ID>
<type>AA_LABEL</type>
<position>269,-3480.5</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2204</ID>
<type>BA_TRI_STATE</type>
<position>139,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>1647 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2205</ID>
<type>AE_DFF_LOW</type>
<position>152,-227.5</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1648 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2206</ID>
<type>BA_TRI_STATE</type>
<position>162,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>1648 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2207</ID>
<type>AE_DFF_LOW</type>
<position>175,-227.5</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>3157 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2208</ID>
<type>BA_TRI_STATE</type>
<position>185,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>3157 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2209</ID>
<type>AE_DFF_LOW</type>
<position>200,-227.5</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>3158 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2210</ID>
<type>BA_TRI_STATE</type>
<position>210,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>3158 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4158</ID>
<type>AE_DFF_LOW</type>
<position>223,-227.5</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>3159 </output>
<input>
<ID>clock</ID>3160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4159</ID>
<type>BA_TRI_STATE</type>
<position>233,-238</position>
<input>
<ID>ENABLE_0</ID>3161 </input>
<input>
<ID>IN_0</ID>3159 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4160</ID>
<type>AA_AND2</type>
<position>30.5,-210</position>
<input>
<ID>IN_0</ID>3192 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>3170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4161</ID>
<type>AA_AND2</type>
<position>41.5,-219.5</position>
<input>
<ID>IN_0</ID>3192 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>3171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4162</ID>
<type>AE_DFF_LOW</type>
<position>58,-209</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>3162 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4163</ID>
<type>BA_TRI_STATE</type>
<position>68,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3162 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4164</ID>
<type>AE_DFF_LOW</type>
<position>81,-209</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>3163 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4165</ID>
<type>BA_TRI_STATE</type>
<position>91,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3163 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4166</ID>
<type>AE_DFF_LOW</type>
<position>106,-209</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>3164 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4167</ID>
<type>BA_TRI_STATE</type>
<position>116,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3164 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4168</ID>
<type>AE_DFF_LOW</type>
<position>129,-209</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>3165 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4169</ID>
<type>BA_TRI_STATE</type>
<position>139,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3165 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4170</ID>
<type>AE_DFF_LOW</type>
<position>152,-209</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>3166 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4171</ID>
<type>BA_TRI_STATE</type>
<position>162,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3166 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4172</ID>
<type>AE_DFF_LOW</type>
<position>175,-209</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>3167 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4173</ID>
<type>BA_TRI_STATE</type>
<position>185,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3167 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4174</ID>
<type>AE_DFF_LOW</type>
<position>200,-209</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>3168 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4175</ID>
<type>BA_TRI_STATE</type>
<position>210,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3168 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4176</ID>
<type>AE_DFF_LOW</type>
<position>223,-209</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>3169 </output>
<input>
<ID>clock</ID>3170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4177</ID>
<type>BA_TRI_STATE</type>
<position>233,-219.5</position>
<input>
<ID>ENABLE_0</ID>3171 </input>
<input>
<ID>IN_0</ID>3169 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4178</ID>
<type>HA_JUNC_2</type>
<position>49.5,-122.5</position>
<input>
<ID>N_in0</ID>3172 </input>
<input>
<ID>N_in1</ID>3200 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4179</ID>
<type>HA_JUNC_2</type>
<position>72.5,-122</position>
<input>
<ID>N_in0</ID>3173 </input>
<input>
<ID>N_in1</ID>3201 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4180</ID>
<type>HA_JUNC_2</type>
<position>75.5,-122.5</position>
<input>
<ID>N_in0</ID>3174 </input>
<input>
<ID>N_in1</ID>3202 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4181</ID>
<type>HA_JUNC_2</type>
<position>95,-122</position>
<input>
<ID>N_in0</ID>3175 </input>
<input>
<ID>N_in1</ID>3203 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4182</ID>
<type>HA_JUNC_2</type>
<position>98.5,-122</position>
<input>
<ID>N_in0</ID>3176 </input>
<input>
<ID>N_in1</ID>3204 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4183</ID>
<type>HA_JUNC_2</type>
<position>119.5,-122.5</position>
<input>
<ID>N_in0</ID>3177 </input>
<input>
<ID>N_in1</ID>3205 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4184</ID>
<type>HA_JUNC_2</type>
<position>123.5,-122</position>
<input>
<ID>N_in0</ID>3178 </input>
<input>
<ID>N_in1</ID>3206 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4185</ID>
<type>HA_JUNC_2</type>
<position>142,-122</position>
<input>
<ID>N_in0</ID>3179 </input>
<input>
<ID>N_in1</ID>3207 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4186</ID>
<type>HA_JUNC_2</type>
<position>146,-122</position>
<input>
<ID>N_in0</ID>3180 </input>
<input>
<ID>N_in1</ID>3208 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4187</ID>
<type>HA_JUNC_2</type>
<position>165,-122</position>
<input>
<ID>N_in0</ID>3181 </input>
<input>
<ID>N_in1</ID>3209 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4188</ID>
<type>HA_JUNC_2</type>
<position>170,-122</position>
<input>
<ID>N_in0</ID>3182 </input>
<input>
<ID>N_in1</ID>3210 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4189</ID>
<type>HA_JUNC_2</type>
<position>192.5,-122</position>
<input>
<ID>N_in0</ID>3184 </input>
<input>
<ID>N_in1</ID>3212 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4190</ID>
<type>HA_JUNC_2</type>
<position>188,-122</position>
<input>
<ID>N_in0</ID>3183 </input>
<input>
<ID>N_in1</ID>3211 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4191</ID>
<type>HA_JUNC_2</type>
<position>213.5,-122.5</position>
<input>
<ID>N_in0</ID>3185 </input>
<input>
<ID>N_in1</ID>3213 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4192</ID>
<type>HA_JUNC_2</type>
<position>238,-123.5</position>
<input>
<ID>N_in0</ID>3187 </input>
<input>
<ID>N_in1</ID>3215 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4193</ID>
<type>AA_AND2</type>
<position>30.5,-188</position>
<input>
<ID>IN_0</ID>3191 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>1127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4194</ID>
<type>AA_AND2</type>
<position>42,-197.5</position>
<input>
<ID>IN_0</ID>3191 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>1128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4195</ID>
<type>HA_JUNC_2</type>
<position>49.5,-289.5</position>
<input>
<ID>N_in1</ID>3172 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4196</ID>
<type>AE_DFF_LOW</type>
<position>58,-187</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1119 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4197</ID>
<type>HA_JUNC_2</type>
<position>72.5,-289</position>
<input>
<ID>N_in1</ID>3173 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4198</ID>
<type>HA_JUNC_2</type>
<position>75.5,-289</position>
<input>
<ID>N_in1</ID>3174 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4199</ID>
<type>HA_JUNC_2</type>
<position>95,-289</position>
<input>
<ID>N_in1</ID>3175 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4200</ID>
<type>HA_JUNC_2</type>
<position>98.5,-289</position>
<input>
<ID>N_in1</ID>3176 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4201</ID>
<type>HA_JUNC_2</type>
<position>119.5,-289</position>
<input>
<ID>N_in1</ID>3177 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4202</ID>
<type>BA_TRI_STATE</type>
<position>68,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4203</ID>
<type>HA_JUNC_2</type>
<position>123.5,-289</position>
<input>
<ID>N_in1</ID>3178 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4204</ID>
<type>HA_JUNC_2</type>
<position>142,-289</position>
<input>
<ID>N_in1</ID>3179 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4205</ID>
<type>HA_JUNC_2</type>
<position>146,-289</position>
<input>
<ID>N_in1</ID>3180 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4206</ID>
<type>HA_JUNC_2</type>
<position>165,-288.5</position>
<input>
<ID>N_in1</ID>3181 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4207</ID>
<type>HA_JUNC_2</type>
<position>170,-288.5</position>
<input>
<ID>N_in1</ID>3182 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4208</ID>
<type>HA_JUNC_2</type>
<position>188,-288</position>
<input>
<ID>N_in1</ID>3183 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4209</ID>
<type>HA_JUNC_2</type>
<position>192.5,-288</position>
<input>
<ID>N_in1</ID>3184 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4210</ID>
<type>HA_JUNC_2</type>
<position>213.5,-287.5</position>
<input>
<ID>N_in1</ID>3185 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4211</ID>
<type>HA_JUNC_2</type>
<position>217,-287.5</position>
<input>
<ID>N_in1</ID>3186 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4212</ID>
<type>HA_JUNC_2</type>
<position>217,-122.5</position>
<input>
<ID>N_in0</ID>3186 </input>
<input>
<ID>N_in1</ID>3214 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4213</ID>
<type>HA_JUNC_2</type>
<position>238,-287.5</position>
<input>
<ID>N_in1</ID>3187 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4214</ID>
<type>AE_DFF_LOW</type>
<position>81,-187</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1120 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4215</ID>
<type>BA_TRI_STATE</type>
<position>91,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1120 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4216</ID>
<type>HA_JUNC_2</type>
<position>36.5,-122.5</position>
<input>
<ID>N_in0</ID>3197 </input>
<input>
<ID>N_in1</ID>3199 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4217</ID>
<type>AE_DFF_LOW</type>
<position>106,-187</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1121 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4218</ID>
<type>HA_JUNC_2</type>
<position>26.5,-122.5</position>
<input>
<ID>N_in0</ID>3196 </input>
<input>
<ID>N_in1</ID>3198 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4219</ID>
<type>BA_TRI_STATE</type>
<position>116,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1121 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4220</ID>
<type>HA_JUNC_2</type>
<position>36.5,-289.5</position>
<input>
<ID>N_in1</ID>3197 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4221</ID>
<type>AE_DFF_LOW</type>
<position>129,-187</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1122 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4222</ID>
<type>HA_JUNC_2</type>
<position>26.5,-289.5</position>
<input>
<ID>N_in1</ID>3196 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4223</ID>
<type>BA_TRI_STATE</type>
<position>139,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1122 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4224</ID>
<type>AE_DFF_LOW</type>
<position>152,-187</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1123 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4225</ID>
<type>AA_LABEL</type>
<position>17.5,-123</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4226</ID>
<type>BA_TRI_STATE</type>
<position>162,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1123 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4227</ID>
<type>AE_DFF_LOW</type>
<position>175,-187</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>1124 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4228</ID>
<type>BA_TRI_STATE</type>
<position>185,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1124 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4229</ID>
<type>AE_DFF_LOW</type>
<position>200,-187</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>1125 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4230</ID>
<type>BA_TRI_STATE</type>
<position>210,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1125 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4231</ID>
<type>AE_DFF_LOW</type>
<position>223,-187</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>1126 </output>
<input>
<ID>clock</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4232</ID>
<type>BA_TRI_STATE</type>
<position>233,-197.5</position>
<input>
<ID>ENABLE_0</ID>1128 </input>
<input>
<ID>IN_0</ID>1126 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4233</ID>
<type>AA_AND2</type>
<position>30.5,-169.5</position>
<input>
<ID>IN_0</ID>3190 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>1137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4234</ID>
<type>AA_AND2</type>
<position>42,-179</position>
<input>
<ID>IN_0</ID>3190 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>1138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4235</ID>
<type>AE_DFF_LOW</type>
<position>58,-168.5</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1129 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4236</ID>
<type>BA_TRI_STATE</type>
<position>68,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1129 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4237</ID>
<type>AE_DFF_LOW</type>
<position>81,-168.5</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1130 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4238</ID>
<type>BA_TRI_STATE</type>
<position>91,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1130 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4239</ID>
<type>AE_DFF_LOW</type>
<position>106,-168.5</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1131 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4240</ID>
<type>BA_TRI_STATE</type>
<position>116,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1131 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4241</ID>
<type>AE_DFF_LOW</type>
<position>129,-168.5</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1132 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4242</ID>
<type>BA_TRI_STATE</type>
<position>139,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1132 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4243</ID>
<type>AE_DFF_LOW</type>
<position>152,-168.5</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1133 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4244</ID>
<type>BA_TRI_STATE</type>
<position>162,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1133 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4245</ID>
<type>AE_DFF_LOW</type>
<position>175,-168.5</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>1134 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4246</ID>
<type>BA_TRI_STATE</type>
<position>185,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1134 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4247</ID>
<type>AE_DFF_LOW</type>
<position>200,-168.5</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>1135 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4248</ID>
<type>BA_TRI_STATE</type>
<position>210,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1135 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4249</ID>
<type>AE_DFF_LOW</type>
<position>223,-168.5</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>1136 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4250</ID>
<type>BA_TRI_STATE</type>
<position>233,-179</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1136 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4251</ID>
<type>AA_AND2</type>
<position>30.5,-150.5</position>
<input>
<ID>IN_0</ID>3189 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>1147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4252</ID>
<type>AA_AND2</type>
<position>42,-160</position>
<input>
<ID>IN_0</ID>3189 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>1148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4253</ID>
<type>AE_DFF_LOW</type>
<position>58,-149.5</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1139 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4254</ID>
<type>BA_TRI_STATE</type>
<position>68,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1139 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4255</ID>
<type>AE_DFF_LOW</type>
<position>81,-149.5</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1140 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4256</ID>
<type>BA_TRI_STATE</type>
<position>91,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1140 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4257</ID>
<type>AE_DFF_LOW</type>
<position>106,-149.5</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1141 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4258</ID>
<type>BA_TRI_STATE</type>
<position>116,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1141 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4259</ID>
<type>AE_DFF_LOW</type>
<position>129,-149.5</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1142 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4260</ID>
<type>BA_TRI_STATE</type>
<position>139,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1142 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4261</ID>
<type>AE_DFF_LOW</type>
<position>152,-149.5</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1143 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4262</ID>
<type>BA_TRI_STATE</type>
<position>162,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1143 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4263</ID>
<type>AE_DFF_LOW</type>
<position>175,-149.5</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>1144 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4264</ID>
<type>BA_TRI_STATE</type>
<position>185,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1144 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4265</ID>
<type>AE_DFF_LOW</type>
<position>200,-149.5</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>1145 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4266</ID>
<type>BA_TRI_STATE</type>
<position>210,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1145 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4267</ID>
<type>AE_DFF_LOW</type>
<position>223,-149.5</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>1146 </output>
<input>
<ID>clock</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4268</ID>
<type>BA_TRI_STATE</type>
<position>233,-160</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1146 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4269</ID>
<type>AA_AND2</type>
<position>30.5,-132</position>
<input>
<ID>IN_0</ID>3188 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>1157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4270</ID>
<type>AA_AND2</type>
<position>42,-141.5</position>
<input>
<ID>IN_0</ID>3188 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>1158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4271</ID>
<type>AE_DFF_LOW</type>
<position>58,-131</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1149 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4272</ID>
<type>BA_TRI_STATE</type>
<position>68,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1149 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4273</ID>
<type>AE_DFF_LOW</type>
<position>81,-131</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1150 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4274</ID>
<type>BA_TRI_STATE</type>
<position>91,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1150 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4275</ID>
<type>AE_DFF_LOW</type>
<position>106,-131</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1151 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4276</ID>
<type>BA_TRI_STATE</type>
<position>116,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1151 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4277</ID>
<type>AE_DFF_LOW</type>
<position>129,-131</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1152 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4278</ID>
<type>BA_TRI_STATE</type>
<position>139,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1152 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4279</ID>
<type>AE_DFF_LOW</type>
<position>152,-131</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1153 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4280</ID>
<type>BA_TRI_STATE</type>
<position>162,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1153 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4281</ID>
<type>AE_DFF_LOW</type>
<position>175,-131</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>1154 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4282</ID>
<type>BA_TRI_STATE</type>
<position>185,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1154 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4283</ID>
<type>AE_DFF_LOW</type>
<position>200,-131</position>
<input>
<ID>IN_0</ID>3184 </input>
<output>
<ID>OUT_0</ID>1155 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4284</ID>
<type>BA_TRI_STATE</type>
<position>210,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1155 </input>
<output>
<ID>OUT_0</ID>3185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4285</ID>
<type>AE_DFF_LOW</type>
<position>223,-131</position>
<input>
<ID>IN_0</ID>3186 </input>
<output>
<ID>OUT_0</ID>1156 </output>
<input>
<ID>clock</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4286</ID>
<type>BA_TRI_STATE</type>
<position>233,-141.5</position>
<input>
<ID>ENABLE_0</ID>1158 </input>
<input>
<ID>IN_0</ID>1156 </input>
<output>
<ID>OUT_0</ID>3187 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4287</ID>
<type>AA_AND2</type>
<position>30.5,-266</position>
<input>
<ID>IN_0</ID>3195 </input>
<input>
<ID>IN_1</ID>3196 </input>
<output>
<ID>OUT</ID>1167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4288</ID>
<type>AA_AND2</type>
<position>41.5,-275.5</position>
<input>
<ID>IN_0</ID>3195 </input>
<input>
<ID>IN_1</ID>3197 </input>
<output>
<ID>OUT</ID>1168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4289</ID>
<type>AE_DFF_LOW</type>
<position>58,-265</position>
<input>
<ID>IN_0</ID>3172 </input>
<output>
<ID>OUT_0</ID>1159 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4290</ID>
<type>BA_TRI_STATE</type>
<position>68,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1159 </input>
<output>
<ID>OUT_0</ID>3173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4291</ID>
<type>AE_DFF_LOW</type>
<position>81,-265</position>
<input>
<ID>IN_0</ID>3174 </input>
<output>
<ID>OUT_0</ID>1160 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4292</ID>
<type>BA_TRI_STATE</type>
<position>91,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1160 </input>
<output>
<ID>OUT_0</ID>3175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4293</ID>
<type>AE_DFF_LOW</type>
<position>106,-265</position>
<input>
<ID>IN_0</ID>3176 </input>
<output>
<ID>OUT_0</ID>1161 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4294</ID>
<type>BA_TRI_STATE</type>
<position>116,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1161 </input>
<output>
<ID>OUT_0</ID>3177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4295</ID>
<type>AE_DFF_LOW</type>
<position>129,-265</position>
<input>
<ID>IN_0</ID>3178 </input>
<output>
<ID>OUT_0</ID>1162 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4296</ID>
<type>BA_TRI_STATE</type>
<position>139,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1162 </input>
<output>
<ID>OUT_0</ID>3179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4297</ID>
<type>AE_DFF_LOW</type>
<position>152,-265</position>
<input>
<ID>IN_0</ID>3180 </input>
<output>
<ID>OUT_0</ID>1163 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4298</ID>
<type>BA_TRI_STATE</type>
<position>162,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1163 </input>
<output>
<ID>OUT_0</ID>3181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4299</ID>
<type>AE_DFF_LOW</type>
<position>175,-265</position>
<input>
<ID>IN_0</ID>3182 </input>
<output>
<ID>OUT_0</ID>1164 </output>
<input>
<ID>clock</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4300</ID>
<type>BA_TRI_STATE</type>
<position>185,-275.5</position>
<input>
<ID>ENABLE_0</ID>1168 </input>
<input>
<ID>IN_0</ID>1164 </input>
<output>
<ID>OUT_0</ID>3183 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4301</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-491</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3356 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4302</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-431</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3269 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4303</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3356 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4304</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3269 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4305</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-491</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3357 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4306</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-431</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3270 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4307</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3357 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4308</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3270 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4309</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-491</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3358 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4310</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-431</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3271 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4311</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3358 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4312</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3271 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4313</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-491</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3359 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4314</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-431</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3272 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4315</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3359 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4316</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3272 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4317</ID>
<type>AA_AND2</type>
<position>31,-626</position>
<input>
<ID>IN_0</ID>3425 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4318</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-431</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3273 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4319</ID>
<type>AA_AND2</type>
<position>42,-635.5</position>
<input>
<ID>IN_0</ID>3425 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3371 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4320</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3273 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4321</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-625</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3362 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4322</ID>
<type>AA_AND2</type>
<position>42,-598</position>
<input>
<ID>IN_0</ID>3423 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3391 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4323</ID>
<type>AA_AND2</type>
<position>31,-413</position>
<input>
<ID>IN_0</ID>3317 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3284 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4324</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3362 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4325</ID>
<type>AA_AND2</type>
<position>42,-422.5</position>
<input>
<ID>IN_0</ID>3317 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3285 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4326</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-625</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3363 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4327</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-587.5</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3382 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4328</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-412</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3276 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4329</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3363 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4330</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3276 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4331</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-625</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3364 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4332</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3382 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4333</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-412</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3277 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4334</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3364 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4335</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3277 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4336</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-625</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3365 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4337</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-587.5</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3383 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4338</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-412</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3278 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4339</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3365 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4340</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3278 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4341</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-625</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3366 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4342</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3383 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4343</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-412</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3279 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4344</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3366 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4345</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3279 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4346</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-625</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3367 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4347</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-587.5</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3384 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4348</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-412</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3280 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4349</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3367 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4350</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3280 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4351</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3384 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4352</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-412</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3281 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4353</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3281 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4354</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-587.5</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3385 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4355</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-412</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3282 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4356</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3282 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4357</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-412</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3283 </output>
<input>
<ID>clock</ID>3284 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4358</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-422.5</position>
<input>
<ID>ENABLE_0</ID>3285 </input>
<input>
<ID>IN_0</ID>3283 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4359</ID>
<type>AA_AND2</type>
<position>31,-394.5</position>
<input>
<ID>IN_0</ID>3316 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3294 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4360</ID>
<type>AA_AND2</type>
<position>42,-404</position>
<input>
<ID>IN_0</ID>3316 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3295 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4361</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-393.5</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3286 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4362</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3286 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4363</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-393.5</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3287 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4364</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3287 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4365</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-393.5</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3288 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4366</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3288 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4367</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-393.5</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3289 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4368</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3289 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4369</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-393.5</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3290 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4370</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3290 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4371</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-393.5</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3291 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4372</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3291 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4373</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-393.5</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3292 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4374</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3292 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4375</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-393.5</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3293 </output>
<input>
<ID>clock</ID>3294 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4376</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-404</position>
<input>
<ID>ENABLE_0</ID>3295 </input>
<input>
<ID>IN_0</ID>3293 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4377</ID>
<type>HA_JUNC_2</type>
<position>50,-307</position>
<input>
<ID>N_in0</ID>3296 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4378</ID>
<type>HA_JUNC_2</type>
<position>73,-306.5</position>
<input>
<ID>N_in0</ID>3297 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4379</ID>
<type>HA_JUNC_2</type>
<position>76,-307</position>
<input>
<ID>N_in0</ID>3298 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4380</ID>
<type>HA_JUNC_2</type>
<position>95.5,-306.5</position>
<input>
<ID>N_in0</ID>3299 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4381</ID>
<type>HA_JUNC_2</type>
<position>99,-306.5</position>
<input>
<ID>N_in0</ID>3300 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4382</ID>
<type>HA_JUNC_2</type>
<position>120,-307</position>
<input>
<ID>N_in0</ID>3301 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4383</ID>
<type>HA_JUNC_2</type>
<position>124,-306.5</position>
<input>
<ID>N_in0</ID>3302 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4384</ID>
<type>HA_JUNC_2</type>
<position>142.5,-306.5</position>
<input>
<ID>N_in0</ID>3303 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4385</ID>
<type>HA_JUNC_2</type>
<position>146.5,-306.5</position>
<input>
<ID>N_in0</ID>3304 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4386</ID>
<type>HA_JUNC_2</type>
<position>165.5,-306.5</position>
<input>
<ID>N_in0</ID>3305 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4387</ID>
<type>HA_JUNC_2</type>
<position>170.5,-306.5</position>
<input>
<ID>N_in0</ID>3306 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4388</ID>
<type>HA_JUNC_2</type>
<position>193,-306.5</position>
<input>
<ID>N_in0</ID>3308 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4389</ID>
<type>HA_JUNC_2</type>
<position>188.5,-306.5</position>
<input>
<ID>N_in0</ID>3307 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4390</ID>
<type>HA_JUNC_2</type>
<position>214,-307</position>
<input>
<ID>N_in0</ID>3309 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4391</ID>
<type>HA_JUNC_2</type>
<position>238.5,-308</position>
<input>
<ID>N_in0</ID>3311 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4392</ID>
<type>HA_JUNC_2</type>
<position>50,-474</position>
<input>
<ID>N_in0</ID>3430 </input>
<input>
<ID>N_in1</ID>3296 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4393</ID>
<type>HA_JUNC_2</type>
<position>73,-473.5</position>
<input>
<ID>N_in0</ID>3431 </input>
<input>
<ID>N_in1</ID>3297 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4394</ID>
<type>HA_JUNC_2</type>
<position>76,-473.5</position>
<input>
<ID>N_in0</ID>3432 </input>
<input>
<ID>N_in1</ID>3298 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4395</ID>
<type>HA_JUNC_2</type>
<position>95.5,-473.5</position>
<input>
<ID>N_in0</ID>3433 </input>
<input>
<ID>N_in1</ID>3299 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4396</ID>
<type>HA_JUNC_2</type>
<position>99,-473.5</position>
<input>
<ID>N_in0</ID>3434 </input>
<input>
<ID>N_in1</ID>3300 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4397</ID>
<type>HA_JUNC_2</type>
<position>120,-473.5</position>
<input>
<ID>N_in0</ID>3435 </input>
<input>
<ID>N_in1</ID>3301 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4398</ID>
<type>HA_JUNC_2</type>
<position>124,-473.5</position>
<input>
<ID>N_in0</ID>3436 </input>
<input>
<ID>N_in1</ID>3302 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4399</ID>
<type>HA_JUNC_2</type>
<position>142.5,-473.5</position>
<input>
<ID>N_in0</ID>3437 </input>
<input>
<ID>N_in1</ID>3303 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4400</ID>
<type>HA_JUNC_2</type>
<position>146.5,-473.5</position>
<input>
<ID>N_in0</ID>3438 </input>
<input>
<ID>N_in1</ID>3304 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4401</ID>
<type>HA_JUNC_2</type>
<position>165.5,-473</position>
<input>
<ID>N_in0</ID>3439 </input>
<input>
<ID>N_in1</ID>3305 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4402</ID>
<type>HA_JUNC_2</type>
<position>170.5,-473</position>
<input>
<ID>N_in0</ID>3440 </input>
<input>
<ID>N_in1</ID>3306 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4403</ID>
<type>HA_JUNC_2</type>
<position>188.5,-472.5</position>
<input>
<ID>N_in0</ID>3441 </input>
<input>
<ID>N_in1</ID>3307 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4404</ID>
<type>HA_JUNC_2</type>
<position>193,-472.5</position>
<input>
<ID>N_in0</ID>3442 </input>
<input>
<ID>N_in1</ID>3308 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4405</ID>
<type>HA_JUNC_2</type>
<position>214,-472</position>
<input>
<ID>N_in0</ID>3443 </input>
<input>
<ID>N_in1</ID>3309 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4406</ID>
<type>HA_JUNC_2</type>
<position>217.5,-472</position>
<input>
<ID>N_in0</ID>3444 </input>
<input>
<ID>N_in1</ID>3310 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4407</ID>
<type>HA_JUNC_2</type>
<position>217.5,-307</position>
<input>
<ID>N_in0</ID>3310 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4408</ID>
<type>HA_JUNC_2</type>
<position>238.5,-472</position>
<input>
<ID>N_in0</ID>3445 </input>
<input>
<ID>N_in1</ID>3311 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4409</ID>
<type>HA_JUNC_2</type>
<position>37,-307</position>
<input>
<ID>N_in0</ID>3321 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4410</ID>
<type>HA_JUNC_2</type>
<position>27,-307</position>
<input>
<ID>N_in0</ID>3320 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4411</ID>
<type>HA_JUNC_2</type>
<position>37,-474</position>
<input>
<ID>N_in0</ID>3429 </input>
<input>
<ID>N_in1</ID>3321 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4412</ID>
<type>HA_JUNC_2</type>
<position>27,-474</position>
<input>
<ID>N_in0</ID>3428 </input>
<input>
<ID>N_in1</ID>3320 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4413</ID>
<type>AA_LABEL</type>
<position>18,-307.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4414</ID>
<type>BI_DECODER_4x16</type>
<position>-121.5,-474.5</position>
<output>
<ID>OUT_0</ID>3425 </output>
<output>
<ID>OUT_1</ID>3424 </output>
<output>
<ID>OUT_10</ID>3317 </output>
<output>
<ID>OUT_11</ID>3316 </output>
<output>
<ID>OUT_12</ID>3315 </output>
<output>
<ID>OUT_13</ID>3314 </output>
<output>
<ID>OUT_14</ID>3313 </output>
<output>
<ID>OUT_15</ID>3312 </output>
<output>
<ID>OUT_2</ID>3423 </output>
<output>
<ID>OUT_3</ID>3422 </output>
<output>
<ID>OUT_4</ID>3421 </output>
<output>
<ID>OUT_5</ID>3420 </output>
<output>
<ID>OUT_6</ID>3419 </output>
<output>
<ID>OUT_7</ID>3418 </output>
<output>
<ID>OUT_8</ID>3319 </output>
<output>
<ID>OUT_9</ID>3318 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4415</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-625</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3368 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4416</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3368 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4417</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-625</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3369 </output>
<input>
<ID>clock</ID>3370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4418</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-635.5</position>
<input>
<ID>ENABLE_0</ID>3371 </input>
<input>
<ID>IN_0</ID>3369 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4419</ID>
<type>AA_AND2</type>
<position>31,-607.5</position>
<input>
<ID>IN_0</ID>3424 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4420</ID>
<type>AA_AND2</type>
<position>42,-617</position>
<input>
<ID>IN_0</ID>3424 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3381 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4421</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-606.5</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3372 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4422</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3372 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4423</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-606.5</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3373 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4424</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3373 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4425</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-606.5</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3374 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4426</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3374 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4427</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-606.5</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3375 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4428</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3375 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4429</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-606.5</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3376 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4430</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3376 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4431</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-606.5</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3377 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4432</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3377 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4433</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-606.5</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3378 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4434</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3378 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4435</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-606.5</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3379 </output>
<input>
<ID>clock</ID>3380 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4436</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-617</position>
<input>
<ID>ENABLE_0</ID>3381 </input>
<input>
<ID>IN_0</ID>3379 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4437</ID>
<type>AA_AND2</type>
<position>31,-588.5</position>
<input>
<ID>IN_0</ID>3423 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3390 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4438</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3385 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4439</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-587.5</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3386 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4440</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3386 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4441</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-587.5</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3387 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4442</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3387 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4443</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-587.5</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3388 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4444</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3388 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4445</ID>
<type>AA_AND2</type>
<position>31,-372.5</position>
<input>
<ID>IN_0</ID>3315 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4446</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-587.5</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3389 </output>
<input>
<ID>clock</ID>3390 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4447</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-598</position>
<input>
<ID>ENABLE_0</ID>3391 </input>
<input>
<ID>IN_0</ID>3389 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4448</ID>
<type>AA_AND2</type>
<position>31,-570</position>
<input>
<ID>IN_0</ID>3422 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3400 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4449</ID>
<type>AA_AND2</type>
<position>42,-579.5</position>
<input>
<ID>IN_0</ID>3422 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4450</ID>
<type>AA_AND2</type>
<position>42.5,-382</position>
<input>
<ID>IN_0</ID>3315 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4451</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-569</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3392 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4452</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3392 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4453</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-569</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3393 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4454</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3393 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4455</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-371.5</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3216 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4456</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-569</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3394 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4457</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3394 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4458</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-569</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3395 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4459</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3395 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4460</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-569</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3396 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4461</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3216 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4462</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3396 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4463</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-569</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3397 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4464</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3397 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4465</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-569</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3398 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4466</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3398 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4467</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-569</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3399 </output>
<input>
<ID>clock</ID>3400 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4468</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-579.5</position>
<input>
<ID>ENABLE_0</ID>3401 </input>
<input>
<ID>IN_0</ID>3399 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4469</ID>
<type>HA_JUNC_2</type>
<position>50,-482.5</position>
<input>
<ID>N_in0</ID>3402 </input>
<input>
<ID>N_in1</ID>3430 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4470</ID>
<type>HA_JUNC_2</type>
<position>73,-482</position>
<input>
<ID>N_in0</ID>3403 </input>
<input>
<ID>N_in1</ID>3431 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4471</ID>
<type>HA_JUNC_2</type>
<position>76,-482.5</position>
<input>
<ID>N_in0</ID>3404 </input>
<input>
<ID>N_in1</ID>3432 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4472</ID>
<type>HA_JUNC_2</type>
<position>95.5,-482</position>
<input>
<ID>N_in0</ID>3405 </input>
<input>
<ID>N_in1</ID>3433 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4473</ID>
<type>HA_JUNC_2</type>
<position>99,-482</position>
<input>
<ID>N_in0</ID>3406 </input>
<input>
<ID>N_in1</ID>3434 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4474</ID>
<type>HA_JUNC_2</type>
<position>120,-482.5</position>
<input>
<ID>N_in0</ID>3407 </input>
<input>
<ID>N_in1</ID>3435 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4475</ID>
<type>HA_JUNC_2</type>
<position>124,-482</position>
<input>
<ID>N_in0</ID>3408 </input>
<input>
<ID>N_in1</ID>3436 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4476</ID>
<type>HA_JUNC_2</type>
<position>142.5,-482</position>
<input>
<ID>N_in0</ID>3409 </input>
<input>
<ID>N_in1</ID>3437 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4477</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-371.5</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3217 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4478</ID>
<type>HA_JUNC_2</type>
<position>146.5,-482</position>
<input>
<ID>N_in0</ID>3410 </input>
<input>
<ID>N_in1</ID>3438 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4479</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3217 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4480</ID>
<type>HA_JUNC_2</type>
<position>165.5,-482</position>
<input>
<ID>N_in0</ID>3411 </input>
<input>
<ID>N_in1</ID>3439 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4481</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-371.5</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3218 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4482</ID>
<type>HA_JUNC_2</type>
<position>170.5,-482</position>
<input>
<ID>N_in0</ID>3412 </input>
<input>
<ID>N_in1</ID>3440 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4483</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3218 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4484</ID>
<type>HA_JUNC_2</type>
<position>193,-482</position>
<input>
<ID>N_in0</ID>3414 </input>
<input>
<ID>N_in1</ID>3442 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4485</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-371.5</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3219 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4486</ID>
<type>HA_JUNC_2</type>
<position>188.5,-482</position>
<input>
<ID>N_in0</ID>3413 </input>
<input>
<ID>N_in1</ID>3441 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4487</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3219 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4488</ID>
<type>HA_JUNC_2</type>
<position>214,-482.5</position>
<input>
<ID>N_in0</ID>3415 </input>
<input>
<ID>N_in1</ID>3443 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4489</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-371.5</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3220 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4490</ID>
<type>HA_JUNC_2</type>
<position>238.5,-483.5</position>
<input>
<ID>N_in0</ID>3417 </input>
<input>
<ID>N_in1</ID>3445 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4491</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3220 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4492</ID>
<type>AA_AND2</type>
<position>31,-548</position>
<input>
<ID>IN_0</ID>3421 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3330 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4493</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-371.5</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3221 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4494</ID>
<type>AA_AND2</type>
<position>42.5,-557.5</position>
<input>
<ID>IN_0</ID>3421 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3331 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4495</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3221 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4496</ID>
<type>HA_JUNC_2</type>
<position>50,-649.5</position>
<input>
<ID>N_in1</ID>3402 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4497</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-371.5</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3222 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4498</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-547</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3322 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4499</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3222 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4500</ID>
<type>HA_JUNC_2</type>
<position>73,-649</position>
<input>
<ID>N_in1</ID>3403 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4501</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-371.5</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3223 </output>
<input>
<ID>clock</ID>3224 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4502</ID>
<type>HA_JUNC_2</type>
<position>76,-649</position>
<input>
<ID>N_in1</ID>3404 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4503</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-382</position>
<input>
<ID>ENABLE_0</ID>3225 </input>
<input>
<ID>IN_0</ID>3223 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4504</ID>
<type>HA_JUNC_2</type>
<position>95.5,-649</position>
<input>
<ID>N_in1</ID>3405 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4505</ID>
<type>AA_AND2</type>
<position>31,-354</position>
<input>
<ID>IN_0</ID>3314 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4506</ID>
<type>HA_JUNC_2</type>
<position>99,-649</position>
<input>
<ID>N_in1</ID>3406 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4507</ID>
<type>AA_AND2</type>
<position>42.5,-363.5</position>
<input>
<ID>IN_0</ID>3314 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4508</ID>
<type>HA_JUNC_2</type>
<position>120,-649</position>
<input>
<ID>N_in1</ID>3407 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4509</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-353</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3226 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4510</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3322 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4511</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3226 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4512</ID>
<type>HA_JUNC_2</type>
<position>124,-649</position>
<input>
<ID>N_in1</ID>3408 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4513</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-353</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3227 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4514</ID>
<type>HA_JUNC_2</type>
<position>142.5,-649</position>
<input>
<ID>N_in1</ID>3409 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4515</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3227 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4516</ID>
<type>HA_JUNC_2</type>
<position>146.5,-649</position>
<input>
<ID>N_in1</ID>3410 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4517</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-353</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3228 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4518</ID>
<type>HA_JUNC_2</type>
<position>165.5,-648.5</position>
<input>
<ID>N_in1</ID>3411 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4519</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3228 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4520</ID>
<type>HA_JUNC_2</type>
<position>170.5,-648.5</position>
<input>
<ID>N_in1</ID>3412 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4521</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-353</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3229 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4522</ID>
<type>HA_JUNC_2</type>
<position>188.5,-648</position>
<input>
<ID>N_in1</ID>3413 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4523</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3229 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4524</ID>
<type>HA_JUNC_2</type>
<position>193,-648</position>
<input>
<ID>N_in1</ID>3414 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4525</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-353</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3230 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4526</ID>
<type>HA_JUNC_2</type>
<position>214,-647.5</position>
<input>
<ID>N_in1</ID>3415 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4527</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3230 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4528</ID>
<type>HA_JUNC_2</type>
<position>217.5,-647.5</position>
<input>
<ID>N_in1</ID>3416 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4529</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-353</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3231 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4530</ID>
<type>HA_JUNC_2</type>
<position>217.5,-482.5</position>
<input>
<ID>N_in0</ID>3416 </input>
<input>
<ID>N_in1</ID>3444 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4531</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3231 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4532</ID>
<type>HA_JUNC_2</type>
<position>238.5,-647.5</position>
<input>
<ID>N_in1</ID>3417 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4533</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-353</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3232 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4534</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-547</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3323 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4535</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3232 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4536</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3323 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4537</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-353</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3233 </output>
<input>
<ID>clock</ID>3234 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4538</ID>
<type>HA_JUNC_2</type>
<position>37,-482.5</position>
<input>
<ID>N_in0</ID>3427 </input>
<input>
<ID>N_in1</ID>3429 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4539</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-363.5</position>
<input>
<ID>ENABLE_0</ID>3235 </input>
<input>
<ID>IN_0</ID>3233 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4540</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-547</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3324 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4541</ID>
<type>AA_AND2</type>
<position>31,-335</position>
<input>
<ID>IN_0</ID>3313 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4542</ID>
<type>HA_JUNC_2</type>
<position>27,-482.5</position>
<input>
<ID>N_in0</ID>3426 </input>
<input>
<ID>N_in1</ID>3428 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4543</ID>
<type>AA_AND2</type>
<position>42.5,-344.5</position>
<input>
<ID>IN_0</ID>3313 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4544</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3324 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4545</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-334</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3236 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4546</ID>
<type>HA_JUNC_2</type>
<position>37,-649.5</position>
<input>
<ID>N_in1</ID>3427 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4547</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3236 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4548</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-547</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3325 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4549</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-334</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3237 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4550</ID>
<type>HA_JUNC_2</type>
<position>27,-649.5</position>
<input>
<ID>N_in1</ID>3426 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4551</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3237 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4552</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3325 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4553</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-334</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3238 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4554</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-547</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3326 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4555</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3238 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4556</ID>
<type>AA_LABEL</type>
<position>18,-483</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4557</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-334</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3239 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4558</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3326 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4559</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3239 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4560</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-547</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3327 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4561</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-334</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3240 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4562</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3327 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4563</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3240 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4564</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-547</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3328 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4565</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-334</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3241 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4566</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3328 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4567</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3241 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4568</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-547</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3329 </output>
<input>
<ID>clock</ID>3330 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4569</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-334</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3242 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4570</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-557.5</position>
<input>
<ID>ENABLE_0</ID>3331 </input>
<input>
<ID>IN_0</ID>3329 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4571</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3242 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4572</ID>
<type>AA_AND2</type>
<position>31,-529.5</position>
<input>
<ID>IN_0</ID>3420 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4573</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-334</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3243 </output>
<input>
<ID>clock</ID>3244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4574</ID>
<type>AA_AND2</type>
<position>42.5,-539</position>
<input>
<ID>IN_0</ID>3420 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4575</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-344.5</position>
<input>
<ID>ENABLE_0</ID>3245 </input>
<input>
<ID>IN_0</ID>3243 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4576</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-528.5</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3332 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4577</ID>
<type>AA_AND2</type>
<position>31,-316.5</position>
<input>
<ID>IN_0</ID>3312 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4578</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3332 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4579</ID>
<type>AA_AND2</type>
<position>42.5,-326</position>
<input>
<ID>IN_0</ID>3312 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4580</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-528.5</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3333 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4581</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-315.5</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3246 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4582</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3333 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4583</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3246 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4584</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-528.5</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3334 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4585</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-315.5</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3247 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4586</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3334 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4587</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3247 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4588</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-528.5</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3335 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4589</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-315.5</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3248 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4590</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3335 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4591</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3248 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4592</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-528.5</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3336 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4593</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-315.5</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3249 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4594</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3336 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4595</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3249 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4596</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-528.5</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3337 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4597</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-315.5</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3250 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4598</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3337 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4599</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3250 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4600</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-528.5</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3338 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4601</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-315.5</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3251 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4602</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3338 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4603</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3251 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4604</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-528.5</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3339 </output>
<input>
<ID>clock</ID>3340 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4605</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-315.5</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3252 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4606</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-539</position>
<input>
<ID>ENABLE_0</ID>3341 </input>
<input>
<ID>IN_0</ID>3339 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4607</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3252 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4608</ID>
<type>AA_AND2</type>
<position>31,-510.5</position>
<input>
<ID>IN_0</ID>3419 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4609</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-315.5</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3253 </output>
<input>
<ID>clock</ID>3254 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4610</ID>
<type>AA_AND2</type>
<position>42.5,-520</position>
<input>
<ID>IN_0</ID>3419 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3351 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4611</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-326</position>
<input>
<ID>ENABLE_0</ID>3255 </input>
<input>
<ID>IN_0</ID>3253 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4612</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-509.5</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3342 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4613</ID>
<type>AA_AND2</type>
<position>31,-450.5</position>
<input>
<ID>IN_0</ID>3319 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3264 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4614</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3342 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4615</ID>
<type>AA_AND2</type>
<position>42,-460</position>
<input>
<ID>IN_0</ID>3319 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4616</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-509.5</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3343 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4617</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-449.5</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3256 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4618</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3343 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4619</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3256 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4620</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-509.5</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3344 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4621</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-449.5</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3257 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4622</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3344 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4623</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3257 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4624</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-509.5</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3345 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4625</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-449.5</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3258 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4626</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3345 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4627</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3258 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4628</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-509.5</position>
<input>
<ID>IN_0</ID>3410 </input>
<output>
<ID>OUT_0</ID>3346 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4629</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-449.5</position>
<input>
<ID>IN_0</ID>3302 </input>
<output>
<ID>OUT_0</ID>3259 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4630</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3346 </input>
<output>
<ID>OUT_0</ID>3411 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4631</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3259 </input>
<output>
<ID>OUT_0</ID>3303 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4632</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-509.5</position>
<input>
<ID>IN_0</ID>3412 </input>
<output>
<ID>OUT_0</ID>3347 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4633</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-449.5</position>
<input>
<ID>IN_0</ID>3304 </input>
<output>
<ID>OUT_0</ID>3260 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4634</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3347 </input>
<output>
<ID>OUT_0</ID>3413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4635</ID>
<type>BA_TRI_STATE</type>
<position>162.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3260 </input>
<output>
<ID>OUT_0</ID>3305 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4636</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-509.5</position>
<input>
<ID>IN_0</ID>3414 </input>
<output>
<ID>OUT_0</ID>3348 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4637</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-449.5</position>
<input>
<ID>IN_0</ID>3306 </input>
<output>
<ID>OUT_0</ID>3261 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4638</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3348 </input>
<output>
<ID>OUT_0</ID>3415 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4639</ID>
<type>BA_TRI_STATE</type>
<position>185.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3261 </input>
<output>
<ID>OUT_0</ID>3307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4640</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-509.5</position>
<input>
<ID>IN_0</ID>3416 </input>
<output>
<ID>OUT_0</ID>3349 </output>
<input>
<ID>clock</ID>3350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4641</ID>
<type>AE_DFF_LOW</type>
<position>200.5,-449.5</position>
<input>
<ID>IN_0</ID>3308 </input>
<output>
<ID>OUT_0</ID>3262 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4642</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-520</position>
<input>
<ID>ENABLE_0</ID>3351 </input>
<input>
<ID>IN_0</ID>3349 </input>
<output>
<ID>OUT_0</ID>3417 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4643</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3262 </input>
<output>
<ID>OUT_0</ID>3309 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4644</ID>
<type>AA_AND2</type>
<position>31,-492</position>
<input>
<ID>IN_0</ID>3418 </input>
<input>
<ID>IN_1</ID>3426 </input>
<output>
<ID>OUT</ID>3360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4645</ID>
<type>AE_DFF_LOW</type>
<position>223.5,-449.5</position>
<input>
<ID>IN_0</ID>3310 </input>
<output>
<ID>OUT_0</ID>3263 </output>
<input>
<ID>clock</ID>3264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4646</ID>
<type>AA_AND2</type>
<position>42.5,-501.5</position>
<input>
<ID>IN_0</ID>3418 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3361 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4647</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-460</position>
<input>
<ID>ENABLE_0</ID>3265 </input>
<input>
<ID>IN_0</ID>3263 </input>
<output>
<ID>OUT_0</ID>3311 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4648</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-491</position>
<input>
<ID>IN_0</ID>3402 </input>
<output>
<ID>OUT_0</ID>3352 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4649</ID>
<type>AA_AND2</type>
<position>31,-432</position>
<input>
<ID>IN_0</ID>3318 </input>
<input>
<ID>IN_1</ID>3320 </input>
<output>
<ID>OUT</ID>3274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4650</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3352 </input>
<output>
<ID>OUT_0</ID>3403 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4651</ID>
<type>AA_AND2</type>
<position>42,-441.5</position>
<input>
<ID>IN_0</ID>3318 </input>
<input>
<ID>IN_1</ID>3321 </input>
<output>
<ID>OUT</ID>3275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4652</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-491</position>
<input>
<ID>IN_0</ID>3404 </input>
<output>
<ID>OUT_0</ID>3353 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4653</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-431</position>
<input>
<ID>IN_0</ID>3296 </input>
<output>
<ID>OUT_0</ID>3266 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4654</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3353 </input>
<output>
<ID>OUT_0</ID>3405 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4655</ID>
<type>BA_TRI_STATE</type>
<position>68.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3266 </input>
<output>
<ID>OUT_0</ID>3297 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4656</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-491</position>
<input>
<ID>IN_0</ID>3406 </input>
<output>
<ID>OUT_0</ID>3354 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4657</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-431</position>
<input>
<ID>IN_0</ID>3298 </input>
<output>
<ID>OUT_0</ID>3267 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4658</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3354 </input>
<output>
<ID>OUT_0</ID>3407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4659</ID>
<type>BA_TRI_STATE</type>
<position>91.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3267 </input>
<output>
<ID>OUT_0</ID>3299 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4660</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-491</position>
<input>
<ID>IN_0</ID>3408 </input>
<output>
<ID>OUT_0</ID>3355 </output>
<input>
<ID>clock</ID>3360 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4661</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-431</position>
<input>
<ID>IN_0</ID>3300 </input>
<output>
<ID>OUT_0</ID>3268 </output>
<input>
<ID>clock</ID>3274 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4662</ID>
<type>BA_TRI_STATE</type>
<position>139.5,-501.5</position>
<input>
<ID>ENABLE_0</ID>3361 </input>
<input>
<ID>IN_0</ID>3355 </input>
<output>
<ID>OUT_0</ID>3409 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4663</ID>
<type>BA_TRI_STATE</type>
<position>116.5,-441.5</position>
<input>
<ID>ENABLE_0</ID>3275 </input>
<input>
<ID>IN_0</ID>3268 </input>
<output>
<ID>OUT_0</ID>3301 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4665</ID>
<type>AA_LABEL</type>
<position>274.5,-123</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4666</ID>
<type>AA_LABEL</type>
<position>278.5,-469</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5394</ID>
<type>AE_DFF_LOW</type>
<position>127,-820</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3949 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5395</ID>
<type>BA_TRI_STATE</type>
<position>160,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4036 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5396</ID>
<type>BA_TRI_STATE</type>
<position>137,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3949 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5397</ID>
<type>AE_DFF_LOW</type>
<position>173,-880</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4037 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5398</ID>
<type>AE_DFF_LOW</type>
<position>150,-820</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3950 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5399</ID>
<type>BA_TRI_STATE</type>
<position>183,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4037 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5400</ID>
<type>BA_TRI_STATE</type>
<position>160,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3950 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5401</ID>
<type>AE_DFF_LOW</type>
<position>198,-880</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4038 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5402</ID>
<type>AE_DFF_LOW</type>
<position>173,-820</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3951 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5403</ID>
<type>BA_TRI_STATE</type>
<position>208,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4038 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5404</ID>
<type>BA_TRI_STATE</type>
<position>183,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3951 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5405</ID>
<type>AE_DFF_LOW</type>
<position>221,-880</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4039 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5406</ID>
<type>AE_DFF_LOW</type>
<position>198,-820</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3952 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5407</ID>
<type>BA_TRI_STATE</type>
<position>231,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4039 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5408</ID>
<type>BA_TRI_STATE</type>
<position>208,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3952 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5409</ID>
<type>AA_AND2</type>
<position>28.5,-862.5</position>
<input>
<ID>IN_0</ID>4108 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4050 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5410</ID>
<type>AE_DFF_LOW</type>
<position>221,-820</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3953 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5411</ID>
<type>AA_AND2</type>
<position>40,-872</position>
<input>
<ID>IN_0</ID>4108 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4051 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5412</ID>
<type>BA_TRI_STATE</type>
<position>231,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3953 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5413</ID>
<type>AE_DFF_LOW</type>
<position>56,-861.5</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4042 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5414</ID>
<type>AA_AND2</type>
<position>28.5,-802.5</position>
<input>
<ID>IN_0</ID>4008 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3964 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5415</ID>
<type>BA_TRI_STATE</type>
<position>66,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4042 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5416</ID>
<type>AA_AND2</type>
<position>39.5,-812</position>
<input>
<ID>IN_0</ID>4008 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3965 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5417</ID>
<type>AE_DFF_LOW</type>
<position>79,-861.5</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4043 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5418</ID>
<type>AE_DFF_LOW</type>
<position>56,-801.5</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3956 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5419</ID>
<type>BA_TRI_STATE</type>
<position>89,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4043 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5420</ID>
<type>BA_TRI_STATE</type>
<position>66,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3956 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5421</ID>
<type>AE_DFF_LOW</type>
<position>104,-861.5</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4044 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5422</ID>
<type>AE_DFF_LOW</type>
<position>79,-801.5</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3957 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5423</ID>
<type>BA_TRI_STATE</type>
<position>114,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4044 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5424</ID>
<type>BA_TRI_STATE</type>
<position>89,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3957 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5425</ID>
<type>AE_DFF_LOW</type>
<position>127,-861.5</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4045 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5426</ID>
<type>AE_DFF_LOW</type>
<position>104,-801.5</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3958 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5427</ID>
<type>BA_TRI_STATE</type>
<position>137,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4045 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5428</ID>
<type>BA_TRI_STATE</type>
<position>114,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3958 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5429</ID>
<type>AE_DFF_LOW</type>
<position>150,-861.5</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4046 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5430</ID>
<type>AE_DFF_LOW</type>
<position>127,-801.5</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3959 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5431</ID>
<type>BA_TRI_STATE</type>
<position>160,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4046 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5432</ID>
<type>BA_TRI_STATE</type>
<position>137,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3959 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5433</ID>
<type>AE_DFF_LOW</type>
<position>173,-861.5</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4047 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5434</ID>
<type>AE_DFF_LOW</type>
<position>150,-801.5</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3960 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5435</ID>
<type>BA_TRI_STATE</type>
<position>183,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4047 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5436</ID>
<type>BA_TRI_STATE</type>
<position>160,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3960 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5437</ID>
<type>AE_DFF_LOW</type>
<position>198,-861.5</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4048 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5438</ID>
<type>AE_DFF_LOW</type>
<position>173,-801.5</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3961 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5439</ID>
<type>BA_TRI_STATE</type>
<position>208,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4048 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5440</ID>
<type>BA_TRI_STATE</type>
<position>183,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3961 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5441</ID>
<type>AE_DFF_LOW</type>
<position>221,-861.5</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4049 </output>
<input>
<ID>clock</ID>4050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5442</ID>
<type>AE_DFF_LOW</type>
<position>198,-801.5</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3962 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5443</ID>
<type>BA_TRI_STATE</type>
<position>231,-872</position>
<input>
<ID>ENABLE_0</ID>4051 </input>
<input>
<ID>IN_0</ID>4049 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5444</ID>
<type>BA_TRI_STATE</type>
<position>208,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3962 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5445</ID>
<type>AA_AND2</type>
<position>28.5,-996.5</position>
<input>
<ID>IN_0</ID>4115 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5446</ID>
<type>AE_DFF_LOW</type>
<position>221,-801.5</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3963 </output>
<input>
<ID>clock</ID>3964 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5447</ID>
<type>AA_AND2</type>
<position>39.5,-1006</position>
<input>
<ID>IN_0</ID>4115 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4061 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5448</ID>
<type>BA_TRI_STATE</type>
<position>231,-812</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3963 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5449</ID>
<type>AE_DFF_LOW</type>
<position>56,-995.5</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4052 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5450</ID>
<type>AA_AND2</type>
<position>39.5,-968.5</position>
<input>
<ID>IN_0</ID>4113 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4081 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5451</ID>
<type>AA_AND2</type>
<position>28.5,-783.5</position>
<input>
<ID>IN_0</ID>4007 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3974 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5452</ID>
<type>BA_TRI_STATE</type>
<position>66,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4052 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5453</ID>
<type>AA_AND2</type>
<position>39.5,-793</position>
<input>
<ID>IN_0</ID>4007 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3975 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5454</ID>
<type>AE_DFF_LOW</type>
<position>79,-995.5</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4053 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5455</ID>
<type>AE_DFF_LOW</type>
<position>56,-958</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4072 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5456</ID>
<type>AE_DFF_LOW</type>
<position>56,-782.5</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3966 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5457</ID>
<type>BA_TRI_STATE</type>
<position>89,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4053 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5458</ID>
<type>BA_TRI_STATE</type>
<position>66,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3966 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5459</ID>
<type>AE_DFF_LOW</type>
<position>104,-995.5</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4054 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5460</ID>
<type>BA_TRI_STATE</type>
<position>66,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4072 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5461</ID>
<type>AE_DFF_LOW</type>
<position>79,-782.5</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3967 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5462</ID>
<type>BA_TRI_STATE</type>
<position>114,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4054 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5463</ID>
<type>BA_TRI_STATE</type>
<position>89,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3967 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5464</ID>
<type>AE_DFF_LOW</type>
<position>127,-995.5</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4055 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5465</ID>
<type>AE_DFF_LOW</type>
<position>79,-958</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4073 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5466</ID>
<type>AE_DFF_LOW</type>
<position>104,-782.5</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3968 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5467</ID>
<type>BA_TRI_STATE</type>
<position>137,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4055 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5468</ID>
<type>BA_TRI_STATE</type>
<position>114,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3968 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5469</ID>
<type>AE_DFF_LOW</type>
<position>150,-995.5</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4056 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5470</ID>
<type>BA_TRI_STATE</type>
<position>89,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4073 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5471</ID>
<type>AE_DFF_LOW</type>
<position>127,-782.5</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3969 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5472</ID>
<type>BA_TRI_STATE</type>
<position>160,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4056 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5473</ID>
<type>BA_TRI_STATE</type>
<position>137,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3969 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5474</ID>
<type>AE_DFF_LOW</type>
<position>173,-995.5</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4057 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5475</ID>
<type>AE_DFF_LOW</type>
<position>104,-958</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4074 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5476</ID>
<type>AE_DFF_LOW</type>
<position>150,-782.5</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3970 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5477</ID>
<type>BA_TRI_STATE</type>
<position>183,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4057 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5478</ID>
<type>BA_TRI_STATE</type>
<position>160,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3970 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5479</ID>
<type>BA_TRI_STATE</type>
<position>114,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4074 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5480</ID>
<type>AE_DFF_LOW</type>
<position>173,-782.5</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3971 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5481</ID>
<type>BA_TRI_STATE</type>
<position>183,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3971 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5482</ID>
<type>AE_DFF_LOW</type>
<position>127,-958</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4075 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5483</ID>
<type>AE_DFF_LOW</type>
<position>198,-782.5</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3972 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5484</ID>
<type>BA_TRI_STATE</type>
<position>208,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3972 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5485</ID>
<type>AE_DFF_LOW</type>
<position>221,-782.5</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3973 </output>
<input>
<ID>clock</ID>3974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5486</ID>
<type>BA_TRI_STATE</type>
<position>231,-793</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3973 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5487</ID>
<type>AA_AND2</type>
<position>28.5,-765</position>
<input>
<ID>IN_0</ID>4006 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3984 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5488</ID>
<type>AA_AND2</type>
<position>39.5,-774.5</position>
<input>
<ID>IN_0</ID>4006 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3985 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5489</ID>
<type>AE_DFF_LOW</type>
<position>56,-764</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3976 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5490</ID>
<type>BA_TRI_STATE</type>
<position>66,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3976 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5491</ID>
<type>AE_DFF_LOW</type>
<position>79,-764</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3977 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5492</ID>
<type>BA_TRI_STATE</type>
<position>89,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3977 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5493</ID>
<type>AE_DFF_LOW</type>
<position>104,-764</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3978 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5494</ID>
<type>BA_TRI_STATE</type>
<position>114,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3978 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5495</ID>
<type>AE_DFF_LOW</type>
<position>127,-764</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3979 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5496</ID>
<type>BA_TRI_STATE</type>
<position>137,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3979 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5497</ID>
<type>AE_DFF_LOW</type>
<position>150,-764</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3980 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5498</ID>
<type>BA_TRI_STATE</type>
<position>160,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3980 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5499</ID>
<type>AE_DFF_LOW</type>
<position>173,-764</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3981 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5500</ID>
<type>BA_TRI_STATE</type>
<position>183,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3981 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5501</ID>
<type>AE_DFF_LOW</type>
<position>198,-764</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3982 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5502</ID>
<type>BA_TRI_STATE</type>
<position>208,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3982 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5503</ID>
<type>AE_DFF_LOW</type>
<position>221,-764</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3983 </output>
<input>
<ID>clock</ID>3984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5504</ID>
<type>BA_TRI_STATE</type>
<position>231,-774.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3983 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5505</ID>
<type>HA_JUNC_2</type>
<position>47.5,-677.5</position>
<input>
<ID>N_in0</ID>3986 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5506</ID>
<type>HA_JUNC_2</type>
<position>70.5,-677</position>
<input>
<ID>N_in0</ID>3987 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5507</ID>
<type>HA_JUNC_2</type>
<position>73.5,-677.5</position>
<input>
<ID>N_in0</ID>3988 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5508</ID>
<type>HA_JUNC_2</type>
<position>93,-677</position>
<input>
<ID>N_in0</ID>3989 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5509</ID>
<type>HA_JUNC_2</type>
<position>96.5,-677</position>
<input>
<ID>N_in0</ID>3990 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5510</ID>
<type>HA_JUNC_2</type>
<position>117.5,-677.5</position>
<input>
<ID>N_in0</ID>3991 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5511</ID>
<type>HA_JUNC_2</type>
<position>121.5,-677</position>
<input>
<ID>N_in0</ID>3992 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5512</ID>
<type>HA_JUNC_2</type>
<position>140,-677</position>
<input>
<ID>N_in0</ID>3993 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5513</ID>
<type>HA_JUNC_2</type>
<position>144,-677</position>
<input>
<ID>N_in0</ID>3994 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5514</ID>
<type>HA_JUNC_2</type>
<position>163,-677</position>
<input>
<ID>N_in0</ID>3995 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5515</ID>
<type>HA_JUNC_2</type>
<position>168,-677</position>
<input>
<ID>N_in0</ID>3996 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5516</ID>
<type>HA_JUNC_2</type>
<position>190.5,-677</position>
<input>
<ID>N_in0</ID>3998 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5517</ID>
<type>HA_JUNC_2</type>
<position>186,-677</position>
<input>
<ID>N_in0</ID>3997 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5518</ID>
<type>HA_JUNC_2</type>
<position>211.5,-677.5</position>
<input>
<ID>N_in0</ID>3999 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5519</ID>
<type>HA_JUNC_2</type>
<position>236,-678.5</position>
<input>
<ID>N_in0</ID>4001 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5520</ID>
<type>HA_JUNC_2</type>
<position>47.5,-844.5</position>
<input>
<ID>N_in0</ID>4120 </input>
<input>
<ID>N_in1</ID>3986 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5521</ID>
<type>HA_JUNC_2</type>
<position>70.5,-844</position>
<input>
<ID>N_in0</ID>4121 </input>
<input>
<ID>N_in1</ID>3987 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5522</ID>
<type>HA_JUNC_2</type>
<position>73.5,-844</position>
<input>
<ID>N_in0</ID>4122 </input>
<input>
<ID>N_in1</ID>3988 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5523</ID>
<type>HA_JUNC_2</type>
<position>93,-844</position>
<input>
<ID>N_in0</ID>4123 </input>
<input>
<ID>N_in1</ID>3989 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5524</ID>
<type>HA_JUNC_2</type>
<position>96.5,-844</position>
<input>
<ID>N_in0</ID>4124 </input>
<input>
<ID>N_in1</ID>3990 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5525</ID>
<type>HA_JUNC_2</type>
<position>117.5,-844</position>
<input>
<ID>N_in0</ID>4125 </input>
<input>
<ID>N_in1</ID>3991 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5526</ID>
<type>HA_JUNC_2</type>
<position>121.5,-844</position>
<input>
<ID>N_in0</ID>4126 </input>
<input>
<ID>N_in1</ID>3992 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5527</ID>
<type>HA_JUNC_2</type>
<position>140,-844</position>
<input>
<ID>N_in0</ID>4127 </input>
<input>
<ID>N_in1</ID>3993 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5528</ID>
<type>HA_JUNC_2</type>
<position>144,-844</position>
<input>
<ID>N_in0</ID>4128 </input>
<input>
<ID>N_in1</ID>3994 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5529</ID>
<type>HA_JUNC_2</type>
<position>163,-843.5</position>
<input>
<ID>N_in0</ID>4129 </input>
<input>
<ID>N_in1</ID>3995 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5530</ID>
<type>HA_JUNC_2</type>
<position>168,-843.5</position>
<input>
<ID>N_in0</ID>4130 </input>
<input>
<ID>N_in1</ID>3996 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5531</ID>
<type>HA_JUNC_2</type>
<position>186,-843</position>
<input>
<ID>N_in0</ID>4131 </input>
<input>
<ID>N_in1</ID>3997 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5532</ID>
<type>HA_JUNC_2</type>
<position>190.5,-843</position>
<input>
<ID>N_in0</ID>4132 </input>
<input>
<ID>N_in1</ID>3998 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5533</ID>
<type>HA_JUNC_2</type>
<position>211.5,-842.5</position>
<input>
<ID>N_in0</ID>4133 </input>
<input>
<ID>N_in1</ID>3999 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5534</ID>
<type>HA_JUNC_2</type>
<position>215,-842.5</position>
<input>
<ID>N_in0</ID>4134 </input>
<input>
<ID>N_in1</ID>4000 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5535</ID>
<type>HA_JUNC_2</type>
<position>215,-677.5</position>
<input>
<ID>N_in0</ID>4000 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5536</ID>
<type>HA_JUNC_2</type>
<position>236,-842.5</position>
<input>
<ID>N_in0</ID>4135 </input>
<input>
<ID>N_in1</ID>4001 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5537</ID>
<type>HA_JUNC_2</type>
<position>34.5,-677.5</position>
<input>
<ID>N_in0</ID>4011 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5538</ID>
<type>HA_JUNC_2</type>
<position>24.5,-677.5</position>
<input>
<ID>N_in0</ID>4010 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5539</ID>
<type>HA_JUNC_2</type>
<position>34.5,-844.5</position>
<input>
<ID>N_in0</ID>4119 </input>
<input>
<ID>N_in1</ID>4011 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5540</ID>
<type>HA_JUNC_2</type>
<position>24.5,-844.5</position>
<input>
<ID>N_in0</ID>4118 </input>
<input>
<ID>N_in1</ID>4010 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5541</ID>
<type>AA_LABEL</type>
<position>15.5,-678</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5542</ID>
<type>BI_DECODER_4x16</type>
<position>-124,-845</position>
<output>
<ID>OUT_0</ID>4115 </output>
<output>
<ID>OUT_1</ID>4114 </output>
<output>
<ID>OUT_10</ID>4007 </output>
<output>
<ID>OUT_11</ID>4006 </output>
<output>
<ID>OUT_12</ID>4005 </output>
<output>
<ID>OUT_13</ID>4004 </output>
<output>
<ID>OUT_14</ID>4003 </output>
<output>
<ID>OUT_15</ID>4002 </output>
<output>
<ID>OUT_2</ID>4113 </output>
<output>
<ID>OUT_3</ID>4112 </output>
<output>
<ID>OUT_4</ID>4111 </output>
<output>
<ID>OUT_5</ID>4110 </output>
<output>
<ID>OUT_6</ID>4109 </output>
<output>
<ID>OUT_7</ID>4108 </output>
<output>
<ID>OUT_8</ID>4009 </output>
<output>
<ID>OUT_9</ID>4008 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>5543</ID>
<type>AE_DFF_LOW</type>
<position>198,-995.5</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4058 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5544</ID>
<type>BA_TRI_STATE</type>
<position>208,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4058 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5545</ID>
<type>AE_DFF_LOW</type>
<position>221,-995.5</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4059 </output>
<input>
<ID>clock</ID>4060 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5546</ID>
<type>BA_TRI_STATE</type>
<position>231,-1006</position>
<input>
<ID>ENABLE_0</ID>4061 </input>
<input>
<ID>IN_0</ID>4059 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5547</ID>
<type>AA_AND2</type>
<position>28.5,-978</position>
<input>
<ID>IN_0</ID>4114 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5548</ID>
<type>AA_AND2</type>
<position>39.5,-987.5</position>
<input>
<ID>IN_0</ID>4114 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4071 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5549</ID>
<type>AE_DFF_LOW</type>
<position>56,-977</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4062 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5550</ID>
<type>BA_TRI_STATE</type>
<position>66,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4062 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5551</ID>
<type>AE_DFF_LOW</type>
<position>79,-977</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4063 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5552</ID>
<type>BA_TRI_STATE</type>
<position>89,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4063 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5553</ID>
<type>AE_DFF_LOW</type>
<position>104,-977</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4064 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5554</ID>
<type>BA_TRI_STATE</type>
<position>114,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4064 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5555</ID>
<type>AE_DFF_LOW</type>
<position>127,-977</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4065 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5556</ID>
<type>BA_TRI_STATE</type>
<position>137,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4065 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5557</ID>
<type>AE_DFF_LOW</type>
<position>150,-977</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4066 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5558</ID>
<type>BA_TRI_STATE</type>
<position>160,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4066 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5559</ID>
<type>AE_DFF_LOW</type>
<position>173,-977</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4067 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5560</ID>
<type>BA_TRI_STATE</type>
<position>183,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4067 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5561</ID>
<type>AE_DFF_LOW</type>
<position>198,-977</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4068 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5562</ID>
<type>BA_TRI_STATE</type>
<position>208,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4068 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5563</ID>
<type>AE_DFF_LOW</type>
<position>221,-977</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4069 </output>
<input>
<ID>clock</ID>4070 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5564</ID>
<type>BA_TRI_STATE</type>
<position>231,-987.5</position>
<input>
<ID>ENABLE_0</ID>4071 </input>
<input>
<ID>IN_0</ID>4069 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5565</ID>
<type>AA_AND2</type>
<position>28.5,-959</position>
<input>
<ID>IN_0</ID>4113 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5566</ID>
<type>BA_TRI_STATE</type>
<position>137,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4075 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5567</ID>
<type>AE_DFF_LOW</type>
<position>150,-958</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4076 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5568</ID>
<type>BA_TRI_STATE</type>
<position>160,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4076 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5569</ID>
<type>AE_DFF_LOW</type>
<position>173,-958</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4077 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5570</ID>
<type>BA_TRI_STATE</type>
<position>183,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4077 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5571</ID>
<type>AE_DFF_LOW</type>
<position>198,-958</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4078 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5572</ID>
<type>BA_TRI_STATE</type>
<position>208,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4078 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5573</ID>
<type>AA_AND2</type>
<position>28.5,-743</position>
<input>
<ID>IN_0</ID>4005 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3914 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5574</ID>
<type>AE_DFF_LOW</type>
<position>221,-958</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4079 </output>
<input>
<ID>clock</ID>4080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5575</ID>
<type>BA_TRI_STATE</type>
<position>231,-968.5</position>
<input>
<ID>ENABLE_0</ID>4081 </input>
<input>
<ID>IN_0</ID>4079 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5576</ID>
<type>AA_AND2</type>
<position>28.5,-940.5</position>
<input>
<ID>IN_0</ID>4112 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4090 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5577</ID>
<type>AA_AND2</type>
<position>39.5,-950</position>
<input>
<ID>IN_0</ID>4112 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4091 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5578</ID>
<type>AA_AND2</type>
<position>40,-752.5</position>
<input>
<ID>IN_0</ID>4005 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3915 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5579</ID>
<type>AE_DFF_LOW</type>
<position>56,-939.5</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4082 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5580</ID>
<type>BA_TRI_STATE</type>
<position>66,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4082 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5581</ID>
<type>AE_DFF_LOW</type>
<position>79,-939.5</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4083 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5582</ID>
<type>BA_TRI_STATE</type>
<position>89,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4083 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5583</ID>
<type>AE_DFF_LOW</type>
<position>56,-742</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3906 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5584</ID>
<type>AE_DFF_LOW</type>
<position>104,-939.5</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4084 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5585</ID>
<type>BA_TRI_STATE</type>
<position>114,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4084 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5586</ID>
<type>AE_DFF_LOW</type>
<position>127,-939.5</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4085 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5587</ID>
<type>BA_TRI_STATE</type>
<position>137,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4085 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5588</ID>
<type>AE_DFF_LOW</type>
<position>150,-939.5</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4086 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5589</ID>
<type>BA_TRI_STATE</type>
<position>66,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3906 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5590</ID>
<type>BA_TRI_STATE</type>
<position>160,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4086 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5591</ID>
<type>AE_DFF_LOW</type>
<position>173,-939.5</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4087 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5592</ID>
<type>BA_TRI_STATE</type>
<position>183,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4087 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5593</ID>
<type>AE_DFF_LOW</type>
<position>198,-939.5</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4088 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5594</ID>
<type>BA_TRI_STATE</type>
<position>208,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4088 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5595</ID>
<type>AE_DFF_LOW</type>
<position>221,-939.5</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4089 </output>
<input>
<ID>clock</ID>4090 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5596</ID>
<type>BA_TRI_STATE</type>
<position>231,-950</position>
<input>
<ID>ENABLE_0</ID>4091 </input>
<input>
<ID>IN_0</ID>4089 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5597</ID>
<type>HA_JUNC_2</type>
<position>47.5,-853</position>
<input>
<ID>N_in0</ID>4092 </input>
<input>
<ID>N_in1</ID>4120 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5598</ID>
<type>HA_JUNC_2</type>
<position>70.5,-852.5</position>
<input>
<ID>N_in0</ID>4093 </input>
<input>
<ID>N_in1</ID>4121 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5599</ID>
<type>HA_JUNC_2</type>
<position>73.5,-853</position>
<input>
<ID>N_in0</ID>4094 </input>
<input>
<ID>N_in1</ID>4122 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5600</ID>
<type>HA_JUNC_2</type>
<position>93,-852.5</position>
<input>
<ID>N_in0</ID>4095 </input>
<input>
<ID>N_in1</ID>4123 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5601</ID>
<type>HA_JUNC_2</type>
<position>96.5,-852.5</position>
<input>
<ID>N_in0</ID>4096 </input>
<input>
<ID>N_in1</ID>4124 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5602</ID>
<type>HA_JUNC_2</type>
<position>117.5,-853</position>
<input>
<ID>N_in0</ID>4097 </input>
<input>
<ID>N_in1</ID>4125 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5603</ID>
<type>HA_JUNC_2</type>
<position>121.5,-852.5</position>
<input>
<ID>N_in0</ID>4098 </input>
<input>
<ID>N_in1</ID>4126 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5604</ID>
<type>HA_JUNC_2</type>
<position>140,-852.5</position>
<input>
<ID>N_in0</ID>4099 </input>
<input>
<ID>N_in1</ID>4127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5605</ID>
<type>AE_DFF_LOW</type>
<position>79,-742</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3907 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5606</ID>
<type>HA_JUNC_2</type>
<position>144,-852.5</position>
<input>
<ID>N_in0</ID>4100 </input>
<input>
<ID>N_in1</ID>4128 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5607</ID>
<type>BA_TRI_STATE</type>
<position>89,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3907 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5608</ID>
<type>HA_JUNC_2</type>
<position>163,-852.5</position>
<input>
<ID>N_in0</ID>4101 </input>
<input>
<ID>N_in1</ID>4129 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5609</ID>
<type>AE_DFF_LOW</type>
<position>104,-742</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3908 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5610</ID>
<type>HA_JUNC_2</type>
<position>168,-852.5</position>
<input>
<ID>N_in0</ID>4102 </input>
<input>
<ID>N_in1</ID>4130 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5611</ID>
<type>BA_TRI_STATE</type>
<position>114,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3908 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5612</ID>
<type>HA_JUNC_2</type>
<position>190.5,-852.5</position>
<input>
<ID>N_in0</ID>4104 </input>
<input>
<ID>N_in1</ID>4132 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5613</ID>
<type>AE_DFF_LOW</type>
<position>127,-742</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3909 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5614</ID>
<type>HA_JUNC_2</type>
<position>186,-852.5</position>
<input>
<ID>N_in0</ID>4103 </input>
<input>
<ID>N_in1</ID>4131 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5615</ID>
<type>BA_TRI_STATE</type>
<position>137,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3909 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5616</ID>
<type>HA_JUNC_2</type>
<position>211.5,-853</position>
<input>
<ID>N_in0</ID>4105 </input>
<input>
<ID>N_in1</ID>4133 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5617</ID>
<type>AE_DFF_LOW</type>
<position>150,-742</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3910 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5618</ID>
<type>HA_JUNC_2</type>
<position>236,-854</position>
<input>
<ID>N_in0</ID>4107 </input>
<input>
<ID>N_in1</ID>4135 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5619</ID>
<type>BA_TRI_STATE</type>
<position>160,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3910 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5620</ID>
<type>AA_AND2</type>
<position>28.5,-918.5</position>
<input>
<ID>IN_0</ID>4111 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4020 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5621</ID>
<type>AE_DFF_LOW</type>
<position>173,-742</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3911 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5622</ID>
<type>AA_AND2</type>
<position>40,-928</position>
<input>
<ID>IN_0</ID>4111 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4021 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5623</ID>
<type>BA_TRI_STATE</type>
<position>183,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3911 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5624</ID>
<type>HA_JUNC_2</type>
<position>47.5,-1020</position>
<input>
<ID>N_in1</ID>4092 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5625</ID>
<type>AE_DFF_LOW</type>
<position>198,-742</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3912 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5626</ID>
<type>AE_DFF_LOW</type>
<position>56,-917.5</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4012 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5627</ID>
<type>BA_TRI_STATE</type>
<position>208,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3912 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5628</ID>
<type>HA_JUNC_2</type>
<position>70.5,-1019.5</position>
<input>
<ID>N_in1</ID>4093 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5629</ID>
<type>AE_DFF_LOW</type>
<position>221,-742</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3913 </output>
<input>
<ID>clock</ID>3914 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5630</ID>
<type>HA_JUNC_2</type>
<position>73.5,-1019.5</position>
<input>
<ID>N_in1</ID>4094 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5631</ID>
<type>BA_TRI_STATE</type>
<position>231,-752.5</position>
<input>
<ID>ENABLE_0</ID>3915 </input>
<input>
<ID>IN_0</ID>3913 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5632</ID>
<type>HA_JUNC_2</type>
<position>93,-1019.5</position>
<input>
<ID>N_in1</ID>4095 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5633</ID>
<type>AA_AND2</type>
<position>28.5,-724.5</position>
<input>
<ID>IN_0</ID>4004 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3924 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5634</ID>
<type>HA_JUNC_2</type>
<position>96.5,-1019.5</position>
<input>
<ID>N_in1</ID>4096 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5635</ID>
<type>AA_AND2</type>
<position>40,-734</position>
<input>
<ID>IN_0</ID>4004 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3925 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5636</ID>
<type>HA_JUNC_2</type>
<position>117.5,-1019.5</position>
<input>
<ID>N_in1</ID>4097 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5637</ID>
<type>AE_DFF_LOW</type>
<position>56,-723.5</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3916 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5638</ID>
<type>BA_TRI_STATE</type>
<position>66,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5639</ID>
<type>BA_TRI_STATE</type>
<position>66,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3916 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5640</ID>
<type>HA_JUNC_2</type>
<position>121.5,-1019.5</position>
<input>
<ID>N_in1</ID>4098 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5641</ID>
<type>AE_DFF_LOW</type>
<position>79,-723.5</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3917 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5642</ID>
<type>HA_JUNC_2</type>
<position>140,-1019.5</position>
<input>
<ID>N_in1</ID>4099 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5643</ID>
<type>BA_TRI_STATE</type>
<position>89,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3917 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5644</ID>
<type>HA_JUNC_2</type>
<position>144,-1019.5</position>
<input>
<ID>N_in1</ID>4100 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5645</ID>
<type>AE_DFF_LOW</type>
<position>104,-723.5</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3918 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5646</ID>
<type>HA_JUNC_2</type>
<position>163,-1019</position>
<input>
<ID>N_in1</ID>4101 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5647</ID>
<type>BA_TRI_STATE</type>
<position>114,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3918 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5648</ID>
<type>HA_JUNC_2</type>
<position>168,-1019</position>
<input>
<ID>N_in1</ID>4102 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5649</ID>
<type>AE_DFF_LOW</type>
<position>127,-723.5</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3919 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5650</ID>
<type>HA_JUNC_2</type>
<position>186,-1018.5</position>
<input>
<ID>N_in1</ID>4103 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5651</ID>
<type>BA_TRI_STATE</type>
<position>137,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3919 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5652</ID>
<type>HA_JUNC_2</type>
<position>190.5,-1018.5</position>
<input>
<ID>N_in1</ID>4104 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5653</ID>
<type>AE_DFF_LOW</type>
<position>150,-723.5</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3920 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5654</ID>
<type>HA_JUNC_2</type>
<position>211.5,-1018</position>
<input>
<ID>N_in1</ID>4105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5655</ID>
<type>BA_TRI_STATE</type>
<position>160,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3920 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5656</ID>
<type>HA_JUNC_2</type>
<position>215,-1018</position>
<input>
<ID>N_in1</ID>4106 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5657</ID>
<type>AE_DFF_LOW</type>
<position>173,-723.5</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3921 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5658</ID>
<type>HA_JUNC_2</type>
<position>215,-853</position>
<input>
<ID>N_in0</ID>4106 </input>
<input>
<ID>N_in1</ID>4134 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5659</ID>
<type>BA_TRI_STATE</type>
<position>183,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3921 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5660</ID>
<type>HA_JUNC_2</type>
<position>236,-1018</position>
<input>
<ID>N_in1</ID>4107 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5661</ID>
<type>AE_DFF_LOW</type>
<position>198,-723.5</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3922 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5662</ID>
<type>AE_DFF_LOW</type>
<position>79,-917.5</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4013 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5663</ID>
<type>BA_TRI_STATE</type>
<position>208,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3922 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5664</ID>
<type>BA_TRI_STATE</type>
<position>89,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5665</ID>
<type>AE_DFF_LOW</type>
<position>221,-723.5</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3923 </output>
<input>
<ID>clock</ID>3924 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5666</ID>
<type>HA_JUNC_2</type>
<position>34.5,-853</position>
<input>
<ID>N_in0</ID>4117 </input>
<input>
<ID>N_in1</ID>4119 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5667</ID>
<type>BA_TRI_STATE</type>
<position>231,-734</position>
<input>
<ID>ENABLE_0</ID>3925 </input>
<input>
<ID>IN_0</ID>3923 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5668</ID>
<type>AE_DFF_LOW</type>
<position>104,-917.5</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5669</ID>
<type>AA_AND2</type>
<position>28.5,-705.5</position>
<input>
<ID>IN_0</ID>4003 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3934 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5670</ID>
<type>HA_JUNC_2</type>
<position>24.5,-853</position>
<input>
<ID>N_in0</ID>4116 </input>
<input>
<ID>N_in1</ID>4118 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5671</ID>
<type>AA_AND2</type>
<position>40,-715</position>
<input>
<ID>IN_0</ID>4003 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3935 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5672</ID>
<type>BA_TRI_STATE</type>
<position>114,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4014 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5673</ID>
<type>AE_DFF_LOW</type>
<position>56,-704.5</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3926 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5674</ID>
<type>HA_JUNC_2</type>
<position>34.5,-1020</position>
<input>
<ID>N_in1</ID>4117 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5675</ID>
<type>BA_TRI_STATE</type>
<position>66,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5676</ID>
<type>AE_DFF_LOW</type>
<position>127,-917.5</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5677</ID>
<type>AE_DFF_LOW</type>
<position>79,-704.5</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3927 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5678</ID>
<type>HA_JUNC_2</type>
<position>24.5,-1020</position>
<input>
<ID>N_in1</ID>4116 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5679</ID>
<type>BA_TRI_STATE</type>
<position>89,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3927 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5680</ID>
<type>BA_TRI_STATE</type>
<position>137,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4015 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5681</ID>
<type>AE_DFF_LOW</type>
<position>104,-704.5</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3928 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5682</ID>
<type>AE_DFF_LOW</type>
<position>150,-917.5</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5683</ID>
<type>BA_TRI_STATE</type>
<position>114,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3928 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5684</ID>
<type>AA_LABEL</type>
<position>15.5,-853.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5685</ID>
<type>AE_DFF_LOW</type>
<position>127,-704.5</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3929 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5686</ID>
<type>BA_TRI_STATE</type>
<position>160,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4016 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5687</ID>
<type>BA_TRI_STATE</type>
<position>137,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3929 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5688</ID>
<type>AE_DFF_LOW</type>
<position>173,-917.5</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5689</ID>
<type>AE_DFF_LOW</type>
<position>150,-704.5</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3930 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5690</ID>
<type>BA_TRI_STATE</type>
<position>183,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4017 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5691</ID>
<type>BA_TRI_STATE</type>
<position>160,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3930 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5692</ID>
<type>AE_DFF_LOW</type>
<position>198,-917.5</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5693</ID>
<type>AE_DFF_LOW</type>
<position>173,-704.5</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3931 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5694</ID>
<type>BA_TRI_STATE</type>
<position>208,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4018 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5695</ID>
<type>BA_TRI_STATE</type>
<position>183,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3931 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5696</ID>
<type>AE_DFF_LOW</type>
<position>221,-917.5</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<input>
<ID>clock</ID>4020 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5697</ID>
<type>AE_DFF_LOW</type>
<position>198,-704.5</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3932 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5698</ID>
<type>BA_TRI_STATE</type>
<position>231,-928</position>
<input>
<ID>ENABLE_0</ID>4021 </input>
<input>
<ID>IN_0</ID>4019 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5699</ID>
<type>BA_TRI_STATE</type>
<position>208,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3932 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5700</ID>
<type>AA_AND2</type>
<position>28.5,-900</position>
<input>
<ID>IN_0</ID>4110 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5701</ID>
<type>AE_DFF_LOW</type>
<position>221,-704.5</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3933 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5702</ID>
<type>AA_AND2</type>
<position>40,-909.5</position>
<input>
<ID>IN_0</ID>4110 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4031 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5703</ID>
<type>BA_TRI_STATE</type>
<position>231,-715</position>
<input>
<ID>ENABLE_0</ID>3935 </input>
<input>
<ID>IN_0</ID>3933 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5704</ID>
<type>AE_DFF_LOW</type>
<position>56,-899</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4022 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5705</ID>
<type>AA_AND2</type>
<position>28.5,-687</position>
<input>
<ID>IN_0</ID>4002 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3944 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5706</ID>
<type>BA_TRI_STATE</type>
<position>66,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4022 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5707</ID>
<type>AA_AND2</type>
<position>40,-696.5</position>
<input>
<ID>IN_0</ID>4002 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5708</ID>
<type>AE_DFF_LOW</type>
<position>79,-899</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4023 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5709</ID>
<type>AE_DFF_LOW</type>
<position>56,-686</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3936 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5710</ID>
<type>BA_TRI_STATE</type>
<position>89,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4023 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5711</ID>
<type>BA_TRI_STATE</type>
<position>66,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3936 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5712</ID>
<type>AE_DFF_LOW</type>
<position>104,-899</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4024 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5713</ID>
<type>AE_DFF_LOW</type>
<position>79,-686</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3937 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5714</ID>
<type>BA_TRI_STATE</type>
<position>114,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4024 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5715</ID>
<type>BA_TRI_STATE</type>
<position>89,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3937 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5716</ID>
<type>AE_DFF_LOW</type>
<position>127,-899</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4025 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5717</ID>
<type>AE_DFF_LOW</type>
<position>104,-686</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3938 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5718</ID>
<type>BA_TRI_STATE</type>
<position>137,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4025 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5719</ID>
<type>BA_TRI_STATE</type>
<position>114,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3938 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5720</ID>
<type>AE_DFF_LOW</type>
<position>150,-899</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4026 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5721</ID>
<type>AE_DFF_LOW</type>
<position>127,-686</position>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>3939 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5722</ID>
<type>BA_TRI_STATE</type>
<position>160,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4026 </input>
<output>
<ID>OUT_0</ID>4101 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5723</ID>
<type>BA_TRI_STATE</type>
<position>137,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3939 </input>
<output>
<ID>OUT_0</ID>3993 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5724</ID>
<type>AE_DFF_LOW</type>
<position>173,-899</position>
<input>
<ID>IN_0</ID>4102 </input>
<output>
<ID>OUT_0</ID>4027 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5725</ID>
<type>AE_DFF_LOW</type>
<position>150,-686</position>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>3940 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5726</ID>
<type>BA_TRI_STATE</type>
<position>183,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4027 </input>
<output>
<ID>OUT_0</ID>4103 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5727</ID>
<type>BA_TRI_STATE</type>
<position>160,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3940 </input>
<output>
<ID>OUT_0</ID>3995 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5728</ID>
<type>AE_DFF_LOW</type>
<position>198,-899</position>
<input>
<ID>IN_0</ID>4104 </input>
<output>
<ID>OUT_0</ID>4028 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5729</ID>
<type>AE_DFF_LOW</type>
<position>173,-686</position>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>3941 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5730</ID>
<type>BA_TRI_STATE</type>
<position>208,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4028 </input>
<output>
<ID>OUT_0</ID>4105 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5731</ID>
<type>BA_TRI_STATE</type>
<position>183,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3941 </input>
<output>
<ID>OUT_0</ID>3997 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5732</ID>
<type>AE_DFF_LOW</type>
<position>221,-899</position>
<input>
<ID>IN_0</ID>4106 </input>
<output>
<ID>OUT_0</ID>4029 </output>
<input>
<ID>clock</ID>4030 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5733</ID>
<type>AE_DFF_LOW</type>
<position>198,-686</position>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>3942 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5734</ID>
<type>BA_TRI_STATE</type>
<position>231,-909.5</position>
<input>
<ID>ENABLE_0</ID>4031 </input>
<input>
<ID>IN_0</ID>4029 </input>
<output>
<ID>OUT_0</ID>4107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5735</ID>
<type>BA_TRI_STATE</type>
<position>208,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3942 </input>
<output>
<ID>OUT_0</ID>3999 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5736</ID>
<type>AA_AND2</type>
<position>28.5,-881</position>
<input>
<ID>IN_0</ID>4109 </input>
<input>
<ID>IN_1</ID>4116 </input>
<output>
<ID>OUT</ID>4040 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5737</ID>
<type>AE_DFF_LOW</type>
<position>221,-686</position>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>3943 </output>
<input>
<ID>clock</ID>3944 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5738</ID>
<type>AA_AND2</type>
<position>40,-890.5</position>
<input>
<ID>IN_0</ID>4109 </input>
<input>
<ID>IN_1</ID>4117 </input>
<output>
<ID>OUT</ID>4041 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5739</ID>
<type>BA_TRI_STATE</type>
<position>231,-696.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3943 </input>
<output>
<ID>OUT_0</ID>4001 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5740</ID>
<type>AE_DFF_LOW</type>
<position>56,-880</position>
<input>
<ID>IN_0</ID>4092 </input>
<output>
<ID>OUT_0</ID>4032 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5741</ID>
<type>AA_AND2</type>
<position>28.5,-821</position>
<input>
<ID>IN_0</ID>4009 </input>
<input>
<ID>IN_1</ID>4010 </input>
<output>
<ID>OUT</ID>3954 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5742</ID>
<type>BA_TRI_STATE</type>
<position>66,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4032 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5743</ID>
<type>AA_AND2</type>
<position>39.5,-830.5</position>
<input>
<ID>IN_0</ID>4009 </input>
<input>
<ID>IN_1</ID>4011 </input>
<output>
<ID>OUT</ID>3955 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5744</ID>
<type>AE_DFF_LOW</type>
<position>79,-880</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4033 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5745</ID>
<type>AE_DFF_LOW</type>
<position>56,-820</position>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>3946 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5746</ID>
<type>BA_TRI_STATE</type>
<position>89,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4033 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5747</ID>
<type>BA_TRI_STATE</type>
<position>66,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3946 </input>
<output>
<ID>OUT_0</ID>3987 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5748</ID>
<type>AE_DFF_LOW</type>
<position>104,-880</position>
<input>
<ID>IN_0</ID>4096 </input>
<output>
<ID>OUT_0</ID>4034 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5749</ID>
<type>AE_DFF_LOW</type>
<position>79,-820</position>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>3947 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5750</ID>
<type>BA_TRI_STATE</type>
<position>114,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4034 </input>
<output>
<ID>OUT_0</ID>4097 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5751</ID>
<type>BA_TRI_STATE</type>
<position>89,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3947 </input>
<output>
<ID>OUT_0</ID>3989 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5752</ID>
<type>AE_DFF_LOW</type>
<position>127,-880</position>
<input>
<ID>IN_0</ID>4098 </input>
<output>
<ID>OUT_0</ID>4035 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5753</ID>
<type>AE_DFF_LOW</type>
<position>104,-820</position>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>3948 </output>
<input>
<ID>clock</ID>3954 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5754</ID>
<type>BA_TRI_STATE</type>
<position>137,-890.5</position>
<input>
<ID>ENABLE_0</ID>4041 </input>
<input>
<ID>IN_0</ID>4035 </input>
<output>
<ID>OUT_0</ID>4099 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5755</ID>
<type>BA_TRI_STATE</type>
<position>114,-830.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3948 </input>
<output>
<ID>OUT_0</ID>3991 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5756</ID>
<type>AE_DFF_LOW</type>
<position>150,-880</position>
<input>
<ID>IN_0</ID>4100 </input>
<output>
<ID>OUT_0</ID>4036 </output>
<input>
<ID>clock</ID>4040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5758</ID>
<type>AA_LABEL</type>
<position>275,-837</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5759</ID>
<type>AE_DFF_LOW</type>
<position>124,-1202.5</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4179 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5760</ID>
<type>BA_TRI_STATE</type>
<position>157,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4266 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5761</ID>
<type>BA_TRI_STATE</type>
<position>134,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4179 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5762</ID>
<type>AE_DFF_LOW</type>
<position>170,-1262.5</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4267 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5763</ID>
<type>AE_DFF_LOW</type>
<position>147,-1202.5</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4180 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5764</ID>
<type>BA_TRI_STATE</type>
<position>180,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4267 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5765</ID>
<type>BA_TRI_STATE</type>
<position>157,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4180 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5766</ID>
<type>AE_DFF_LOW</type>
<position>195,-1262.5</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4268 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5767</ID>
<type>AE_DFF_LOW</type>
<position>170,-1202.5</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4181 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5768</ID>
<type>BA_TRI_STATE</type>
<position>205,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4268 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5769</ID>
<type>BA_TRI_STATE</type>
<position>180,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4181 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5770</ID>
<type>AE_DFF_LOW</type>
<position>218,-1262.5</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4269 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5771</ID>
<type>AE_DFF_LOW</type>
<position>195,-1202.5</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4182 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5772</ID>
<type>BA_TRI_STATE</type>
<position>228,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4269 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5773</ID>
<type>BA_TRI_STATE</type>
<position>205,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4182 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5774</ID>
<type>AA_AND2</type>
<position>25.5,-1245</position>
<input>
<ID>IN_0</ID>4338 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4280 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5775</ID>
<type>AE_DFF_LOW</type>
<position>218,-1202.5</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4183 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5776</ID>
<type>AA_AND2</type>
<position>37,-1254.5</position>
<input>
<ID>IN_0</ID>4338 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5777</ID>
<type>BA_TRI_STATE</type>
<position>228,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4183 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5778</ID>
<type>AE_DFF_LOW</type>
<position>53,-1244</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4272 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5779</ID>
<type>AA_AND2</type>
<position>25.5,-1185</position>
<input>
<ID>IN_0</ID>4238 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5780</ID>
<type>BA_TRI_STATE</type>
<position>63,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4272 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5781</ID>
<type>AA_AND2</type>
<position>36.5,-1194.5</position>
<input>
<ID>IN_0</ID>4238 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5782</ID>
<type>AE_DFF_LOW</type>
<position>76,-1244</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4273 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5783</ID>
<type>AE_DFF_LOW</type>
<position>53,-1184</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4186 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5784</ID>
<type>BA_TRI_STATE</type>
<position>86,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4273 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5785</ID>
<type>BA_TRI_STATE</type>
<position>63,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4186 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5786</ID>
<type>AE_DFF_LOW</type>
<position>101,-1244</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4274 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5787</ID>
<type>AE_DFF_LOW</type>
<position>76,-1184</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4187 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5788</ID>
<type>BA_TRI_STATE</type>
<position>111,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4274 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5789</ID>
<type>BA_TRI_STATE</type>
<position>86,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4187 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5790</ID>
<type>AE_DFF_LOW</type>
<position>124,-1244</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4275 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5791</ID>
<type>AE_DFF_LOW</type>
<position>101,-1184</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4188 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5792</ID>
<type>BA_TRI_STATE</type>
<position>134,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4275 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5793</ID>
<type>BA_TRI_STATE</type>
<position>111,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4188 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5794</ID>
<type>AE_DFF_LOW</type>
<position>147,-1244</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4276 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5795</ID>
<type>AE_DFF_LOW</type>
<position>124,-1184</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4189 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5796</ID>
<type>BA_TRI_STATE</type>
<position>157,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4276 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5797</ID>
<type>BA_TRI_STATE</type>
<position>134,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4189 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5798</ID>
<type>AE_DFF_LOW</type>
<position>170,-1244</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4277 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5799</ID>
<type>AE_DFF_LOW</type>
<position>147,-1184</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4190 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5800</ID>
<type>BA_TRI_STATE</type>
<position>180,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4277 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5801</ID>
<type>BA_TRI_STATE</type>
<position>157,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4190 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5802</ID>
<type>AE_DFF_LOW</type>
<position>195,-1244</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4278 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5803</ID>
<type>AE_DFF_LOW</type>
<position>170,-1184</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4191 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5804</ID>
<type>BA_TRI_STATE</type>
<position>205,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4278 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5805</ID>
<type>BA_TRI_STATE</type>
<position>180,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4191 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5806</ID>
<type>AE_DFF_LOW</type>
<position>218,-1244</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4279 </output>
<input>
<ID>clock</ID>4280 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5807</ID>
<type>AE_DFF_LOW</type>
<position>195,-1184</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4192 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5808</ID>
<type>BA_TRI_STATE</type>
<position>228,-1254.5</position>
<input>
<ID>ENABLE_0</ID>4281 </input>
<input>
<ID>IN_0</ID>4279 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5809</ID>
<type>BA_TRI_STATE</type>
<position>205,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4192 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5810</ID>
<type>AA_AND2</type>
<position>25.5,-1379</position>
<input>
<ID>IN_0</ID>4345 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4290 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5811</ID>
<type>AE_DFF_LOW</type>
<position>218,-1184</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4193 </output>
<input>
<ID>clock</ID>4194 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5812</ID>
<type>AA_AND2</type>
<position>36.5,-1388.5</position>
<input>
<ID>IN_0</ID>4345 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4291 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5813</ID>
<type>BA_TRI_STATE</type>
<position>228,-1194.5</position>
<input>
<ID>ENABLE_0</ID>4195 </input>
<input>
<ID>IN_0</ID>4193 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5814</ID>
<type>AE_DFF_LOW</type>
<position>53,-1378</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4282 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5815</ID>
<type>AA_AND2</type>
<position>36.5,-1351</position>
<input>
<ID>IN_0</ID>4343 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4311 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5816</ID>
<type>AA_AND2</type>
<position>25.5,-1166</position>
<input>
<ID>IN_0</ID>4237 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5817</ID>
<type>BA_TRI_STATE</type>
<position>63,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4282 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5818</ID>
<type>AA_AND2</type>
<position>36.5,-1175.5</position>
<input>
<ID>IN_0</ID>4237 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5819</ID>
<type>AE_DFF_LOW</type>
<position>76,-1378</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4283 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5820</ID>
<type>AE_DFF_LOW</type>
<position>53,-1340.5</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4302 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5821</ID>
<type>AE_DFF_LOW</type>
<position>53,-1165</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4196 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5822</ID>
<type>BA_TRI_STATE</type>
<position>86,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4283 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5823</ID>
<type>BA_TRI_STATE</type>
<position>63,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4196 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5824</ID>
<type>AE_DFF_LOW</type>
<position>101,-1378</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4284 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5825</ID>
<type>BA_TRI_STATE</type>
<position>63,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4302 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5826</ID>
<type>AE_DFF_LOW</type>
<position>76,-1165</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4197 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5827</ID>
<type>BA_TRI_STATE</type>
<position>111,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4284 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5828</ID>
<type>BA_TRI_STATE</type>
<position>86,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4197 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5829</ID>
<type>AE_DFF_LOW</type>
<position>124,-1378</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4285 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5830</ID>
<type>AE_DFF_LOW</type>
<position>76,-1340.5</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4303 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5831</ID>
<type>AE_DFF_LOW</type>
<position>101,-1165</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4198 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5832</ID>
<type>BA_TRI_STATE</type>
<position>134,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4285 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5833</ID>
<type>BA_TRI_STATE</type>
<position>111,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4198 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5834</ID>
<type>AE_DFF_LOW</type>
<position>147,-1378</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4286 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5835</ID>
<type>BA_TRI_STATE</type>
<position>86,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4303 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5836</ID>
<type>AE_DFF_LOW</type>
<position>124,-1165</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4199 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5837</ID>
<type>BA_TRI_STATE</type>
<position>157,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4286 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5838</ID>
<type>BA_TRI_STATE</type>
<position>134,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4199 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5839</ID>
<type>AE_DFF_LOW</type>
<position>170,-1378</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4287 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5840</ID>
<type>AE_DFF_LOW</type>
<position>101,-1340.5</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4304 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5841</ID>
<type>AE_DFF_LOW</type>
<position>147,-1165</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4200 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5842</ID>
<type>BA_TRI_STATE</type>
<position>180,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4287 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5843</ID>
<type>BA_TRI_STATE</type>
<position>157,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4200 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5844</ID>
<type>BA_TRI_STATE</type>
<position>111,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4304 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5845</ID>
<type>AE_DFF_LOW</type>
<position>170,-1165</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4201 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5846</ID>
<type>BA_TRI_STATE</type>
<position>180,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4201 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5847</ID>
<type>AE_DFF_LOW</type>
<position>124,-1340.5</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4305 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5848</ID>
<type>AE_DFF_LOW</type>
<position>195,-1165</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4202 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5849</ID>
<type>BA_TRI_STATE</type>
<position>205,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4202 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5850</ID>
<type>AE_DFF_LOW</type>
<position>218,-1165</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4203 </output>
<input>
<ID>clock</ID>4204 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5851</ID>
<type>BA_TRI_STATE</type>
<position>228,-1175.5</position>
<input>
<ID>ENABLE_0</ID>4205 </input>
<input>
<ID>IN_0</ID>4203 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5852</ID>
<type>AA_AND2</type>
<position>25.5,-1147.5</position>
<input>
<ID>IN_0</ID>4236 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5853</ID>
<type>AA_AND2</type>
<position>36.5,-1157</position>
<input>
<ID>IN_0</ID>4236 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5854</ID>
<type>AE_DFF_LOW</type>
<position>53,-1146.5</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4206 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5855</ID>
<type>BA_TRI_STATE</type>
<position>63,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4206 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5856</ID>
<type>AE_DFF_LOW</type>
<position>76,-1146.5</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4207 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5857</ID>
<type>BA_TRI_STATE</type>
<position>86,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4207 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5858</ID>
<type>AE_DFF_LOW</type>
<position>101,-1146.5</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4208 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5859</ID>
<type>BA_TRI_STATE</type>
<position>111,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4208 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5860</ID>
<type>AE_DFF_LOW</type>
<position>124,-1146.5</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4209 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5861</ID>
<type>BA_TRI_STATE</type>
<position>134,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4209 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5862</ID>
<type>AE_DFF_LOW</type>
<position>147,-1146.5</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4210 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5863</ID>
<type>BA_TRI_STATE</type>
<position>157,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4210 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5864</ID>
<type>AE_DFF_LOW</type>
<position>170,-1146.5</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4211 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5865</ID>
<type>BA_TRI_STATE</type>
<position>180,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4211 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5866</ID>
<type>AE_DFF_LOW</type>
<position>195,-1146.5</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4212 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5867</ID>
<type>BA_TRI_STATE</type>
<position>205,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4212 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5868</ID>
<type>AE_DFF_LOW</type>
<position>218,-1146.5</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4213 </output>
<input>
<ID>clock</ID>4214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5869</ID>
<type>BA_TRI_STATE</type>
<position>228,-1157</position>
<input>
<ID>ENABLE_0</ID>4215 </input>
<input>
<ID>IN_0</ID>4213 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5870</ID>
<type>HA_JUNC_2</type>
<position>44.5,-1060</position>
<input>
<ID>N_in0</ID>4216 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5871</ID>
<type>HA_JUNC_2</type>
<position>67.5,-1059.5</position>
<input>
<ID>N_in0</ID>4217 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5872</ID>
<type>HA_JUNC_2</type>
<position>70.5,-1060</position>
<input>
<ID>N_in0</ID>4218 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5873</ID>
<type>HA_JUNC_2</type>
<position>90,-1059.5</position>
<input>
<ID>N_in0</ID>4219 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5874</ID>
<type>HA_JUNC_2</type>
<position>93.5,-1059.5</position>
<input>
<ID>N_in0</ID>4220 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5875</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1060</position>
<input>
<ID>N_in0</ID>4221 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5876</ID>
<type>HA_JUNC_2</type>
<position>118.5,-1059.5</position>
<input>
<ID>N_in0</ID>4222 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5877</ID>
<type>HA_JUNC_2</type>
<position>137,-1059.5</position>
<input>
<ID>N_in0</ID>4223 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5878</ID>
<type>HA_JUNC_2</type>
<position>141,-1059.5</position>
<input>
<ID>N_in0</ID>4224 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5879</ID>
<type>HA_JUNC_2</type>
<position>160,-1059.5</position>
<input>
<ID>N_in0</ID>4225 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5880</ID>
<type>HA_JUNC_2</type>
<position>165,-1059.5</position>
<input>
<ID>N_in0</ID>4226 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5881</ID>
<type>HA_JUNC_2</type>
<position>187.5,-1059.5</position>
<input>
<ID>N_in0</ID>4228 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5882</ID>
<type>HA_JUNC_2</type>
<position>183,-1059.5</position>
<input>
<ID>N_in0</ID>4227 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5883</ID>
<type>HA_JUNC_2</type>
<position>208.5,-1060</position>
<input>
<ID>N_in0</ID>4229 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5884</ID>
<type>HA_JUNC_2</type>
<position>233,-1061</position>
<input>
<ID>N_in0</ID>4231 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5885</ID>
<type>HA_JUNC_2</type>
<position>44.5,-1227</position>
<input>
<ID>N_in0</ID>4350 </input>
<input>
<ID>N_in1</ID>4216 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5886</ID>
<type>HA_JUNC_2</type>
<position>67.5,-1226.5</position>
<input>
<ID>N_in0</ID>4351 </input>
<input>
<ID>N_in1</ID>4217 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5887</ID>
<type>HA_JUNC_2</type>
<position>70.5,-1226.5</position>
<input>
<ID>N_in0</ID>4352 </input>
<input>
<ID>N_in1</ID>4218 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5888</ID>
<type>HA_JUNC_2</type>
<position>90,-1226.5</position>
<input>
<ID>N_in0</ID>4353 </input>
<input>
<ID>N_in1</ID>4219 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5889</ID>
<type>HA_JUNC_2</type>
<position>93.5,-1226.5</position>
<input>
<ID>N_in0</ID>4354 </input>
<input>
<ID>N_in1</ID>4220 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5890</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1226.5</position>
<input>
<ID>N_in0</ID>4355 </input>
<input>
<ID>N_in1</ID>4221 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5891</ID>
<type>HA_JUNC_2</type>
<position>118.5,-1226.5</position>
<input>
<ID>N_in0</ID>4356 </input>
<input>
<ID>N_in1</ID>4222 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5892</ID>
<type>HA_JUNC_2</type>
<position>137,-1226.5</position>
<input>
<ID>N_in0</ID>4357 </input>
<input>
<ID>N_in1</ID>4223 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5893</ID>
<type>HA_JUNC_2</type>
<position>141,-1226.5</position>
<input>
<ID>N_in0</ID>4358 </input>
<input>
<ID>N_in1</ID>4224 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5894</ID>
<type>HA_JUNC_2</type>
<position>160,-1226</position>
<input>
<ID>N_in0</ID>4359 </input>
<input>
<ID>N_in1</ID>4225 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5895</ID>
<type>HA_JUNC_2</type>
<position>165,-1226</position>
<input>
<ID>N_in0</ID>4360 </input>
<input>
<ID>N_in1</ID>4226 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5896</ID>
<type>HA_JUNC_2</type>
<position>183,-1225.5</position>
<input>
<ID>N_in0</ID>4361 </input>
<input>
<ID>N_in1</ID>4227 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5897</ID>
<type>HA_JUNC_2</type>
<position>187.5,-1225.5</position>
<input>
<ID>N_in0</ID>4362 </input>
<input>
<ID>N_in1</ID>4228 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5898</ID>
<type>HA_JUNC_2</type>
<position>208.5,-1225</position>
<input>
<ID>N_in0</ID>4363 </input>
<input>
<ID>N_in1</ID>4229 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5899</ID>
<type>HA_JUNC_2</type>
<position>212,-1225</position>
<input>
<ID>N_in0</ID>4364 </input>
<input>
<ID>N_in1</ID>4230 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5900</ID>
<type>HA_JUNC_2</type>
<position>212,-1060</position>
<input>
<ID>N_in0</ID>4230 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5901</ID>
<type>HA_JUNC_2</type>
<position>233,-1225</position>
<input>
<ID>N_in0</ID>4365 </input>
<input>
<ID>N_in1</ID>4231 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5902</ID>
<type>HA_JUNC_2</type>
<position>31.5,-1060</position>
<input>
<ID>N_in0</ID>4241 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5903</ID>
<type>HA_JUNC_2</type>
<position>21.5,-1060</position>
<input>
<ID>N_in0</ID>4240 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5904</ID>
<type>HA_JUNC_2</type>
<position>31.5,-1227</position>
<input>
<ID>N_in0</ID>4349 </input>
<input>
<ID>N_in1</ID>4241 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5905</ID>
<type>HA_JUNC_2</type>
<position>21.5,-1227</position>
<input>
<ID>N_in0</ID>4348 </input>
<input>
<ID>N_in1</ID>4240 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5906</ID>
<type>AA_LABEL</type>
<position>12.5,-1060.5</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5907</ID>
<type>BI_DECODER_4x16</type>
<position>-127,-1227.5</position>
<output>
<ID>OUT_0</ID>4345 </output>
<output>
<ID>OUT_1</ID>4344 </output>
<output>
<ID>OUT_10</ID>4237 </output>
<output>
<ID>OUT_11</ID>4236 </output>
<output>
<ID>OUT_12</ID>4235 </output>
<output>
<ID>OUT_13</ID>4234 </output>
<output>
<ID>OUT_14</ID>4233 </output>
<output>
<ID>OUT_15</ID>4232 </output>
<output>
<ID>OUT_2</ID>4343 </output>
<output>
<ID>OUT_3</ID>4342 </output>
<output>
<ID>OUT_4</ID>4341 </output>
<output>
<ID>OUT_5</ID>4340 </output>
<output>
<ID>OUT_6</ID>4339 </output>
<output>
<ID>OUT_7</ID>4338 </output>
<output>
<ID>OUT_8</ID>4239 </output>
<output>
<ID>OUT_9</ID>4238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>5908</ID>
<type>AE_DFF_LOW</type>
<position>195,-1378</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4288 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5909</ID>
<type>BA_TRI_STATE</type>
<position>205,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4288 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5910</ID>
<type>AE_DFF_LOW</type>
<position>218,-1378</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4289 </output>
<input>
<ID>clock</ID>4290 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5911</ID>
<type>BA_TRI_STATE</type>
<position>228,-1388.5</position>
<input>
<ID>ENABLE_0</ID>4291 </input>
<input>
<ID>IN_0</ID>4289 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5912</ID>
<type>AA_AND2</type>
<position>25.5,-1360.5</position>
<input>
<ID>IN_0</ID>4344 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4300 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5913</ID>
<type>AA_AND2</type>
<position>36.5,-1370</position>
<input>
<ID>IN_0</ID>4344 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4301 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5914</ID>
<type>AE_DFF_LOW</type>
<position>53,-1359.5</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4292 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5915</ID>
<type>BA_TRI_STATE</type>
<position>63,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4292 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5916</ID>
<type>AE_DFF_LOW</type>
<position>76,-1359.5</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4293 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5917</ID>
<type>BA_TRI_STATE</type>
<position>86,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4293 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5918</ID>
<type>AE_DFF_LOW</type>
<position>101,-1359.5</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4294 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5919</ID>
<type>BA_TRI_STATE</type>
<position>111,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4294 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5920</ID>
<type>AE_DFF_LOW</type>
<position>124,-1359.5</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4295 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5921</ID>
<type>BA_TRI_STATE</type>
<position>134,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4295 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5922</ID>
<type>AE_DFF_LOW</type>
<position>147,-1359.5</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4296 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5923</ID>
<type>BA_TRI_STATE</type>
<position>157,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4296 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5924</ID>
<type>AE_DFF_LOW</type>
<position>170,-1359.5</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4297 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5925</ID>
<type>BA_TRI_STATE</type>
<position>180,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4297 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5926</ID>
<type>AE_DFF_LOW</type>
<position>195,-1359.5</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4298 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5927</ID>
<type>BA_TRI_STATE</type>
<position>205,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4298 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5928</ID>
<type>AE_DFF_LOW</type>
<position>218,-1359.5</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4299 </output>
<input>
<ID>clock</ID>4300 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5929</ID>
<type>BA_TRI_STATE</type>
<position>228,-1370</position>
<input>
<ID>ENABLE_0</ID>4301 </input>
<input>
<ID>IN_0</ID>4299 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5930</ID>
<type>AA_AND2</type>
<position>25.5,-1341.5</position>
<input>
<ID>IN_0</ID>4343 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4310 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5931</ID>
<type>BA_TRI_STATE</type>
<position>134,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4305 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5932</ID>
<type>AE_DFF_LOW</type>
<position>147,-1340.5</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4306 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5933</ID>
<type>BA_TRI_STATE</type>
<position>157,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4306 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5934</ID>
<type>AE_DFF_LOW</type>
<position>170,-1340.5</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4307 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5935</ID>
<type>BA_TRI_STATE</type>
<position>180,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4307 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5936</ID>
<type>AE_DFF_LOW</type>
<position>195,-1340.5</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4308 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5937</ID>
<type>BA_TRI_STATE</type>
<position>205,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4308 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5938</ID>
<type>AA_AND2</type>
<position>25.5,-1125.5</position>
<input>
<ID>IN_0</ID>4235 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5939</ID>
<type>AE_DFF_LOW</type>
<position>218,-1340.5</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4309 </output>
<input>
<ID>clock</ID>4310 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5940</ID>
<type>BA_TRI_STATE</type>
<position>228,-1351</position>
<input>
<ID>ENABLE_0</ID>4311 </input>
<input>
<ID>IN_0</ID>4309 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5941</ID>
<type>AA_AND2</type>
<position>25.5,-1323</position>
<input>
<ID>IN_0</ID>4342 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5942</ID>
<type>AA_AND2</type>
<position>36.5,-1332.5</position>
<input>
<ID>IN_0</ID>4342 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4321 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5943</ID>
<type>AA_AND2</type>
<position>37,-1135</position>
<input>
<ID>IN_0</ID>4235 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5944</ID>
<type>AE_DFF_LOW</type>
<position>53,-1322</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4312 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5945</ID>
<type>BA_TRI_STATE</type>
<position>63,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4312 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5946</ID>
<type>AE_DFF_LOW</type>
<position>76,-1322</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4313 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5947</ID>
<type>BA_TRI_STATE</type>
<position>86,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4313 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5948</ID>
<type>AE_DFF_LOW</type>
<position>53,-1124.5</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4136 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5949</ID>
<type>AE_DFF_LOW</type>
<position>101,-1322</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4314 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5950</ID>
<type>BA_TRI_STATE</type>
<position>111,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4314 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5951</ID>
<type>AE_DFF_LOW</type>
<position>124,-1322</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4315 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5952</ID>
<type>BA_TRI_STATE</type>
<position>134,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4315 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5953</ID>
<type>AE_DFF_LOW</type>
<position>147,-1322</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4316 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5954</ID>
<type>BA_TRI_STATE</type>
<position>63,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4136 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5955</ID>
<type>BA_TRI_STATE</type>
<position>157,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4316 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5956</ID>
<type>AE_DFF_LOW</type>
<position>170,-1322</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4317 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5957</ID>
<type>BA_TRI_STATE</type>
<position>180,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4317 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5958</ID>
<type>AE_DFF_LOW</type>
<position>195,-1322</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4318 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5959</ID>
<type>BA_TRI_STATE</type>
<position>205,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4318 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5960</ID>
<type>AE_DFF_LOW</type>
<position>218,-1322</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4319 </output>
<input>
<ID>clock</ID>4320 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5961</ID>
<type>BA_TRI_STATE</type>
<position>228,-1332.5</position>
<input>
<ID>ENABLE_0</ID>4321 </input>
<input>
<ID>IN_0</ID>4319 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5962</ID>
<type>HA_JUNC_2</type>
<position>44.5,-1235.5</position>
<input>
<ID>N_in0</ID>4322 </input>
<input>
<ID>N_in1</ID>4350 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5963</ID>
<type>HA_JUNC_2</type>
<position>67.5,-1235</position>
<input>
<ID>N_in0</ID>4323 </input>
<input>
<ID>N_in1</ID>4351 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5964</ID>
<type>HA_JUNC_2</type>
<position>70.5,-1235.5</position>
<input>
<ID>N_in0</ID>4324 </input>
<input>
<ID>N_in1</ID>4352 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5965</ID>
<type>HA_JUNC_2</type>
<position>90,-1235</position>
<input>
<ID>N_in0</ID>4325 </input>
<input>
<ID>N_in1</ID>4353 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5966</ID>
<type>HA_JUNC_2</type>
<position>93.5,-1235</position>
<input>
<ID>N_in0</ID>4326 </input>
<input>
<ID>N_in1</ID>4354 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5967</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1235.5</position>
<input>
<ID>N_in0</ID>4327 </input>
<input>
<ID>N_in1</ID>4355 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5968</ID>
<type>HA_JUNC_2</type>
<position>118.5,-1235</position>
<input>
<ID>N_in0</ID>4328 </input>
<input>
<ID>N_in1</ID>4356 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5969</ID>
<type>HA_JUNC_2</type>
<position>137,-1235</position>
<input>
<ID>N_in0</ID>4329 </input>
<input>
<ID>N_in1</ID>4357 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5970</ID>
<type>AE_DFF_LOW</type>
<position>76,-1124.5</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4137 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5971</ID>
<type>HA_JUNC_2</type>
<position>141,-1235</position>
<input>
<ID>N_in0</ID>4330 </input>
<input>
<ID>N_in1</ID>4358 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5972</ID>
<type>BA_TRI_STATE</type>
<position>86,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4137 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5973</ID>
<type>HA_JUNC_2</type>
<position>160,-1235</position>
<input>
<ID>N_in0</ID>4331 </input>
<input>
<ID>N_in1</ID>4359 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5974</ID>
<type>AE_DFF_LOW</type>
<position>101,-1124.5</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4138 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5975</ID>
<type>HA_JUNC_2</type>
<position>165,-1235</position>
<input>
<ID>N_in0</ID>4332 </input>
<input>
<ID>N_in1</ID>4360 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5976</ID>
<type>BA_TRI_STATE</type>
<position>111,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4138 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5977</ID>
<type>HA_JUNC_2</type>
<position>187.5,-1235</position>
<input>
<ID>N_in0</ID>4334 </input>
<input>
<ID>N_in1</ID>4362 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5978</ID>
<type>AE_DFF_LOW</type>
<position>124,-1124.5</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4139 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5979</ID>
<type>HA_JUNC_2</type>
<position>183,-1235</position>
<input>
<ID>N_in0</ID>4333 </input>
<input>
<ID>N_in1</ID>4361 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5980</ID>
<type>BA_TRI_STATE</type>
<position>134,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4139 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5981</ID>
<type>HA_JUNC_2</type>
<position>208.5,-1235.5</position>
<input>
<ID>N_in0</ID>4335 </input>
<input>
<ID>N_in1</ID>4363 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5982</ID>
<type>AE_DFF_LOW</type>
<position>147,-1124.5</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4140 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5983</ID>
<type>HA_JUNC_2</type>
<position>233,-1236.5</position>
<input>
<ID>N_in0</ID>4337 </input>
<input>
<ID>N_in1</ID>4365 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5984</ID>
<type>BA_TRI_STATE</type>
<position>157,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4140 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5985</ID>
<type>AA_AND2</type>
<position>25.5,-1301</position>
<input>
<ID>IN_0</ID>4341 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5986</ID>
<type>AE_DFF_LOW</type>
<position>170,-1124.5</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4141 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5987</ID>
<type>AA_AND2</type>
<position>37,-1310.5</position>
<input>
<ID>IN_0</ID>4341 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5988</ID>
<type>BA_TRI_STATE</type>
<position>180,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4141 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5989</ID>
<type>HA_JUNC_2</type>
<position>44.5,-1402.5</position>
<input>
<ID>N_in1</ID>4322 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5990</ID>
<type>AE_DFF_LOW</type>
<position>195,-1124.5</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4142 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5991</ID>
<type>AE_DFF_LOW</type>
<position>53,-1300</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4242 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5992</ID>
<type>BA_TRI_STATE</type>
<position>205,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4142 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5993</ID>
<type>HA_JUNC_2</type>
<position>67.5,-1402</position>
<input>
<ID>N_in1</ID>4323 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5994</ID>
<type>AE_DFF_LOW</type>
<position>218,-1124.5</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4143 </output>
<input>
<ID>clock</ID>4144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5995</ID>
<type>HA_JUNC_2</type>
<position>70.5,-1402</position>
<input>
<ID>N_in1</ID>4324 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5996</ID>
<type>BA_TRI_STATE</type>
<position>228,-1135</position>
<input>
<ID>ENABLE_0</ID>4145 </input>
<input>
<ID>IN_0</ID>4143 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5997</ID>
<type>HA_JUNC_2</type>
<position>90,-1402</position>
<input>
<ID>N_in1</ID>4325 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5998</ID>
<type>AA_AND2</type>
<position>25.5,-1107</position>
<input>
<ID>IN_0</ID>4234 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5999</ID>
<type>HA_JUNC_2</type>
<position>93.5,-1402</position>
<input>
<ID>N_in1</ID>4326 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6000</ID>
<type>AA_AND2</type>
<position>37,-1116.5</position>
<input>
<ID>IN_0</ID>4234 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6001</ID>
<type>HA_JUNC_2</type>
<position>114.5,-1402</position>
<input>
<ID>N_in1</ID>4327 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6002</ID>
<type>AE_DFF_LOW</type>
<position>53,-1106</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4146 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6003</ID>
<type>BA_TRI_STATE</type>
<position>63,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4242 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6004</ID>
<type>BA_TRI_STATE</type>
<position>63,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4146 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6005</ID>
<type>HA_JUNC_2</type>
<position>118.5,-1402</position>
<input>
<ID>N_in1</ID>4328 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6006</ID>
<type>AE_DFF_LOW</type>
<position>76,-1106</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4147 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6007</ID>
<type>HA_JUNC_2</type>
<position>137,-1402</position>
<input>
<ID>N_in1</ID>4329 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6008</ID>
<type>BA_TRI_STATE</type>
<position>86,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4147 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6009</ID>
<type>HA_JUNC_2</type>
<position>141,-1402</position>
<input>
<ID>N_in1</ID>4330 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6010</ID>
<type>AE_DFF_LOW</type>
<position>101,-1106</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4148 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6011</ID>
<type>HA_JUNC_2</type>
<position>160,-1401.5</position>
<input>
<ID>N_in1</ID>4331 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6012</ID>
<type>BA_TRI_STATE</type>
<position>111,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4148 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6013</ID>
<type>HA_JUNC_2</type>
<position>165,-1401.5</position>
<input>
<ID>N_in1</ID>4332 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6014</ID>
<type>AE_DFF_LOW</type>
<position>124,-1106</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4149 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6015</ID>
<type>HA_JUNC_2</type>
<position>183,-1401</position>
<input>
<ID>N_in1</ID>4333 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6016</ID>
<type>BA_TRI_STATE</type>
<position>134,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4149 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6017</ID>
<type>HA_JUNC_2</type>
<position>187.5,-1401</position>
<input>
<ID>N_in1</ID>4334 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6018</ID>
<type>AE_DFF_LOW</type>
<position>147,-1106</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4150 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6019</ID>
<type>HA_JUNC_2</type>
<position>208.5,-1400.5</position>
<input>
<ID>N_in1</ID>4335 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6020</ID>
<type>BA_TRI_STATE</type>
<position>157,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4150 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6021</ID>
<type>HA_JUNC_2</type>
<position>212,-1400.5</position>
<input>
<ID>N_in1</ID>4336 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6022</ID>
<type>AE_DFF_LOW</type>
<position>170,-1106</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4151 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6023</ID>
<type>HA_JUNC_2</type>
<position>212,-1235.5</position>
<input>
<ID>N_in0</ID>4336 </input>
<input>
<ID>N_in1</ID>4364 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6024</ID>
<type>BA_TRI_STATE</type>
<position>180,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4151 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6025</ID>
<type>HA_JUNC_2</type>
<position>233,-1400.5</position>
<input>
<ID>N_in1</ID>4337 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6026</ID>
<type>AE_DFF_LOW</type>
<position>195,-1106</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4152 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6027</ID>
<type>AE_DFF_LOW</type>
<position>76,-1300</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4243 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6028</ID>
<type>BA_TRI_STATE</type>
<position>205,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4152 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6029</ID>
<type>BA_TRI_STATE</type>
<position>86,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4243 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6030</ID>
<type>AE_DFF_LOW</type>
<position>218,-1106</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4153 </output>
<input>
<ID>clock</ID>4154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6031</ID>
<type>HA_JUNC_2</type>
<position>31.5,-1235.5</position>
<input>
<ID>N_in0</ID>4347 </input>
<input>
<ID>N_in1</ID>4349 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6032</ID>
<type>BA_TRI_STATE</type>
<position>228,-1116.5</position>
<input>
<ID>ENABLE_0</ID>4155 </input>
<input>
<ID>IN_0</ID>4153 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6033</ID>
<type>AE_DFF_LOW</type>
<position>101,-1300</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4244 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6034</ID>
<type>AA_AND2</type>
<position>25.5,-1088</position>
<input>
<ID>IN_0</ID>4233 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6035</ID>
<type>HA_JUNC_2</type>
<position>21.5,-1235.5</position>
<input>
<ID>N_in0</ID>4346 </input>
<input>
<ID>N_in1</ID>4348 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6036</ID>
<type>AA_AND2</type>
<position>37,-1097.5</position>
<input>
<ID>IN_0</ID>4233 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6037</ID>
<type>BA_TRI_STATE</type>
<position>111,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4244 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6038</ID>
<type>AE_DFF_LOW</type>
<position>53,-1087</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4156 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6039</ID>
<type>HA_JUNC_2</type>
<position>31.5,-1402.5</position>
<input>
<ID>N_in1</ID>4347 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6040</ID>
<type>BA_TRI_STATE</type>
<position>63,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4156 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6041</ID>
<type>AE_DFF_LOW</type>
<position>124,-1300</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4245 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6042</ID>
<type>AE_DFF_LOW</type>
<position>76,-1087</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4157 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6043</ID>
<type>HA_JUNC_2</type>
<position>21.5,-1402.5</position>
<input>
<ID>N_in1</ID>4346 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6044</ID>
<type>BA_TRI_STATE</type>
<position>86,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4157 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6045</ID>
<type>BA_TRI_STATE</type>
<position>134,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4245 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6046</ID>
<type>AE_DFF_LOW</type>
<position>101,-1087</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4158 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6047</ID>
<type>AE_DFF_LOW</type>
<position>147,-1300</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4246 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6048</ID>
<type>BA_TRI_STATE</type>
<position>111,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4158 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6049</ID>
<type>AA_LABEL</type>
<position>12.5,-1236</position>
<gparam>LABEL_TEXT CLOCK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6050</ID>
<type>AE_DFF_LOW</type>
<position>124,-1087</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4159 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6051</ID>
<type>BA_TRI_STATE</type>
<position>157,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4246 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6052</ID>
<type>BA_TRI_STATE</type>
<position>134,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4159 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6053</ID>
<type>AE_DFF_LOW</type>
<position>170,-1300</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4247 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6054</ID>
<type>AE_DFF_LOW</type>
<position>147,-1087</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4160 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6055</ID>
<type>BA_TRI_STATE</type>
<position>180,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4247 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6056</ID>
<type>BA_TRI_STATE</type>
<position>157,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4160 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6057</ID>
<type>AE_DFF_LOW</type>
<position>195,-1300</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4248 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6058</ID>
<type>AE_DFF_LOW</type>
<position>170,-1087</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4161 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6059</ID>
<type>BA_TRI_STATE</type>
<position>205,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4248 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6060</ID>
<type>BA_TRI_STATE</type>
<position>180,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4161 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6061</ID>
<type>AE_DFF_LOW</type>
<position>218,-1300</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4249 </output>
<input>
<ID>clock</ID>4250 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6062</ID>
<type>AE_DFF_LOW</type>
<position>195,-1087</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4162 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6063</ID>
<type>BA_TRI_STATE</type>
<position>228,-1310.5</position>
<input>
<ID>ENABLE_0</ID>4251 </input>
<input>
<ID>IN_0</ID>4249 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6064</ID>
<type>BA_TRI_STATE</type>
<position>205,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4162 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6065</ID>
<type>AA_AND2</type>
<position>25.5,-1282.5</position>
<input>
<ID>IN_0</ID>4340 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6066</ID>
<type>AE_DFF_LOW</type>
<position>218,-1087</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4163 </output>
<input>
<ID>clock</ID>4164 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6067</ID>
<type>AA_AND2</type>
<position>37,-1292</position>
<input>
<ID>IN_0</ID>4340 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6068</ID>
<type>BA_TRI_STATE</type>
<position>228,-1097.5</position>
<input>
<ID>ENABLE_0</ID>4165 </input>
<input>
<ID>IN_0</ID>4163 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6069</ID>
<type>AE_DFF_LOW</type>
<position>53,-1281.5</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4252 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6070</ID>
<type>AA_AND2</type>
<position>25.5,-1069.5</position>
<input>
<ID>IN_0</ID>4232 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6071</ID>
<type>BA_TRI_STATE</type>
<position>63,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4252 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6072</ID>
<type>AA_AND2</type>
<position>37,-1079</position>
<input>
<ID>IN_0</ID>4232 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6073</ID>
<type>AE_DFF_LOW</type>
<position>76,-1281.5</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4253 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6074</ID>
<type>AE_DFF_LOW</type>
<position>53,-1068.5</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4166 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6075</ID>
<type>BA_TRI_STATE</type>
<position>86,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4253 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6076</ID>
<type>BA_TRI_STATE</type>
<position>63,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4166 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6077</ID>
<type>AE_DFF_LOW</type>
<position>101,-1281.5</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4254 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6078</ID>
<type>AE_DFF_LOW</type>
<position>76,-1068.5</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4167 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6079</ID>
<type>BA_TRI_STATE</type>
<position>111,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4254 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6080</ID>
<type>BA_TRI_STATE</type>
<position>86,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4167 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6081</ID>
<type>AE_DFF_LOW</type>
<position>124,-1281.5</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4255 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6082</ID>
<type>AE_DFF_LOW</type>
<position>101,-1068.5</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4168 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6083</ID>
<type>BA_TRI_STATE</type>
<position>134,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4255 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6084</ID>
<type>BA_TRI_STATE</type>
<position>111,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4168 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6085</ID>
<type>AE_DFF_LOW</type>
<position>147,-1281.5</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4256 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6086</ID>
<type>AE_DFF_LOW</type>
<position>124,-1068.5</position>
<input>
<ID>IN_0</ID>4222 </input>
<output>
<ID>OUT_0</ID>4169 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6087</ID>
<type>BA_TRI_STATE</type>
<position>157,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4256 </input>
<output>
<ID>OUT_0</ID>4331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6088</ID>
<type>BA_TRI_STATE</type>
<position>134,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4169 </input>
<output>
<ID>OUT_0</ID>4223 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6089</ID>
<type>AE_DFF_LOW</type>
<position>170,-1281.5</position>
<input>
<ID>IN_0</ID>4332 </input>
<output>
<ID>OUT_0</ID>4257 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6090</ID>
<type>AE_DFF_LOW</type>
<position>147,-1068.5</position>
<input>
<ID>IN_0</ID>4224 </input>
<output>
<ID>OUT_0</ID>4170 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6091</ID>
<type>BA_TRI_STATE</type>
<position>180,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4257 </input>
<output>
<ID>OUT_0</ID>4333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6092</ID>
<type>BA_TRI_STATE</type>
<position>157,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4170 </input>
<output>
<ID>OUT_0</ID>4225 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6093</ID>
<type>AE_DFF_LOW</type>
<position>195,-1281.5</position>
<input>
<ID>IN_0</ID>4334 </input>
<output>
<ID>OUT_0</ID>4258 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6094</ID>
<type>AE_DFF_LOW</type>
<position>170,-1068.5</position>
<input>
<ID>IN_0</ID>4226 </input>
<output>
<ID>OUT_0</ID>4171 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6095</ID>
<type>BA_TRI_STATE</type>
<position>205,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4258 </input>
<output>
<ID>OUT_0</ID>4335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6096</ID>
<type>BA_TRI_STATE</type>
<position>180,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4171 </input>
<output>
<ID>OUT_0</ID>4227 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6097</ID>
<type>AE_DFF_LOW</type>
<position>218,-1281.5</position>
<input>
<ID>IN_0</ID>4336 </input>
<output>
<ID>OUT_0</ID>4259 </output>
<input>
<ID>clock</ID>4260 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6098</ID>
<type>AE_DFF_LOW</type>
<position>195,-1068.5</position>
<input>
<ID>IN_0</ID>4228 </input>
<output>
<ID>OUT_0</ID>4172 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6099</ID>
<type>BA_TRI_STATE</type>
<position>228,-1292</position>
<input>
<ID>ENABLE_0</ID>4261 </input>
<input>
<ID>IN_0</ID>4259 </input>
<output>
<ID>OUT_0</ID>4337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6100</ID>
<type>BA_TRI_STATE</type>
<position>205,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4172 </input>
<output>
<ID>OUT_0</ID>4229 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6101</ID>
<type>AA_AND2</type>
<position>25.5,-1263.5</position>
<input>
<ID>IN_0</ID>4339 </input>
<input>
<ID>IN_1</ID>4346 </input>
<output>
<ID>OUT</ID>4270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6102</ID>
<type>AE_DFF_LOW</type>
<position>218,-1068.5</position>
<input>
<ID>IN_0</ID>4230 </input>
<output>
<ID>OUT_0</ID>4173 </output>
<input>
<ID>clock</ID>4174 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6103</ID>
<type>AA_AND2</type>
<position>37,-1273</position>
<input>
<ID>IN_0</ID>4339 </input>
<input>
<ID>IN_1</ID>4347 </input>
<output>
<ID>OUT</ID>4271 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6104</ID>
<type>BA_TRI_STATE</type>
<position>228,-1079</position>
<input>
<ID>ENABLE_0</ID>4175 </input>
<input>
<ID>IN_0</ID>4173 </input>
<output>
<ID>OUT_0</ID>4231 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6105</ID>
<type>AE_DFF_LOW</type>
<position>53,-1262.5</position>
<input>
<ID>IN_0</ID>4322 </input>
<output>
<ID>OUT_0</ID>4262 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6106</ID>
<type>AA_AND2</type>
<position>25.5,-1203.5</position>
<input>
<ID>IN_0</ID>4239 </input>
<input>
<ID>IN_1</ID>4240 </input>
<output>
<ID>OUT</ID>4184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6107</ID>
<type>BA_TRI_STATE</type>
<position>63,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4262 </input>
<output>
<ID>OUT_0</ID>4323 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6108</ID>
<type>AA_AND2</type>
<position>36.5,-1213</position>
<input>
<ID>IN_0</ID>4239 </input>
<input>
<ID>IN_1</ID>4241 </input>
<output>
<ID>OUT</ID>4185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6109</ID>
<type>AE_DFF_LOW</type>
<position>76,-1262.5</position>
<input>
<ID>IN_0</ID>4324 </input>
<output>
<ID>OUT_0</ID>4263 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6110</ID>
<type>AE_DFF_LOW</type>
<position>53,-1202.5</position>
<input>
<ID>IN_0</ID>4216 </input>
<output>
<ID>OUT_0</ID>4176 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6111</ID>
<type>BA_TRI_STATE</type>
<position>86,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4263 </input>
<output>
<ID>OUT_0</ID>4325 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6112</ID>
<type>BA_TRI_STATE</type>
<position>63,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4176 </input>
<output>
<ID>OUT_0</ID>4217 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6113</ID>
<type>AE_DFF_LOW</type>
<position>101,-1262.5</position>
<input>
<ID>IN_0</ID>4326 </input>
<output>
<ID>OUT_0</ID>4264 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6114</ID>
<type>AE_DFF_LOW</type>
<position>76,-1202.5</position>
<input>
<ID>IN_0</ID>4218 </input>
<output>
<ID>OUT_0</ID>4177 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6115</ID>
<type>BA_TRI_STATE</type>
<position>111,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4264 </input>
<output>
<ID>OUT_0</ID>4327 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6116</ID>
<type>BA_TRI_STATE</type>
<position>86,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4177 </input>
<output>
<ID>OUT_0</ID>4219 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6117</ID>
<type>AE_DFF_LOW</type>
<position>124,-1262.5</position>
<input>
<ID>IN_0</ID>4328 </input>
<output>
<ID>OUT_0</ID>4265 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6118</ID>
<type>AE_DFF_LOW</type>
<position>101,-1202.5</position>
<input>
<ID>IN_0</ID>4220 </input>
<output>
<ID>OUT_0</ID>4178 </output>
<input>
<ID>clock</ID>4184 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6119</ID>
<type>BA_TRI_STATE</type>
<position>134,-1273</position>
<input>
<ID>ENABLE_0</ID>4271 </input>
<input>
<ID>IN_0</ID>4265 </input>
<output>
<ID>OUT_0</ID>4329 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6120</ID>
<type>BA_TRI_STATE</type>
<position>111,-1213</position>
<input>
<ID>ENABLE_0</ID>4185 </input>
<input>
<ID>IN_0</ID>4178 </input>
<output>
<ID>OUT_0</ID>4221 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6121</ID>
<type>AE_DFF_LOW</type>
<position>147,-1262.5</position>
<input>
<ID>IN_0</ID>4330 </input>
<output>
<ID>OUT_0</ID>4266 </output>
<input>
<ID>clock</ID>4270 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6123</ID>
<type>AA_LABEL</type>
<position>272,-1225.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 32</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6124</ID>
<type>AE_DFF_LOW</type>
<position>122,-1589.5</position>
<input>
<ID>IN_0</ID>4452 </input>
<output>
<ID>OUT_0</ID>4409 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6125</ID>
<type>BA_TRI_STATE</type>
<position>155,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4496 </input>
<output>
<ID>OUT_0</ID>4561 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6126</ID>
<type>BA_TRI_STATE</type>
<position>132,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4409 </input>
<output>
<ID>OUT_0</ID>4453 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6127</ID>
<type>AE_DFF_LOW</type>
<position>168,-1649.5</position>
<input>
<ID>IN_0</ID>4562 </input>
<output>
<ID>OUT_0</ID>4497 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6128</ID>
<type>AE_DFF_LOW</type>
<position>145,-1589.5</position>
<input>
<ID>IN_0</ID>4454 </input>
<output>
<ID>OUT_0</ID>4410 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6129</ID>
<type>BA_TRI_STATE</type>
<position>178,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4497 </input>
<output>
<ID>OUT_0</ID>4563 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6130</ID>
<type>BA_TRI_STATE</type>
<position>155,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4410 </input>
<output>
<ID>OUT_0</ID>4455 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6131</ID>
<type>AE_DFF_LOW</type>
<position>193,-1649.5</position>
<input>
<ID>IN_0</ID>4564 </input>
<output>
<ID>OUT_0</ID>4498 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6132</ID>
<type>AE_DFF_LOW</type>
<position>168,-1589.5</position>
<input>
<ID>IN_0</ID>4456 </input>
<output>
<ID>OUT_0</ID>4411 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6133</ID>
<type>BA_TRI_STATE</type>
<position>203,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4498 </input>
<output>
<ID>OUT_0</ID>4565 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6134</ID>
<type>BA_TRI_STATE</type>
<position>178,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4411 </input>
<output>
<ID>OUT_0</ID>4457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6135</ID>
<type>AE_DFF_LOW</type>
<position>216,-1649.5</position>
<input>
<ID>IN_0</ID>4566 </input>
<output>
<ID>OUT_0</ID>4499 </output>
<input>
<ID>clock</ID>4500 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6136</ID>
<type>AE_DFF_LOW</type>
<position>193,-1589.5</position>
<input>
<ID>IN_0</ID>4458 </input>
<output>
<ID>OUT_0</ID>4412 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6137</ID>
<type>BA_TRI_STATE</type>
<position>226,-1660</position>
<input>
<ID>ENABLE_0</ID>4501 </input>
<input>
<ID>IN_0</ID>4499 </input>
<output>
<ID>OUT_0</ID>4567 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6138</ID>
<type>BA_TRI_STATE</type>
<position>203,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4412 </input>
<output>
<ID>OUT_0</ID>4459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6139</ID>
<type>AA_AND2</type>
<position>23.5,-1632</position>
<input>
<ID>IN_0</ID>4568 </input>
<input>
<ID>IN_1</ID>4576 </input>
<output>
<ID>OUT</ID>4510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6140</ID>
<type>AE_DFF_LOW</type>
<position>216,-1589.5</position>
<input>
<ID>IN_0</ID>4460 </input>
<output>
<ID>OUT_0</ID>4413 </output>
<input>
<ID>clock</ID>4414 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6141</ID>
<type>AA_AND2</type>
<position>35,-1641.5</position>
<input>
<ID>IN_0</ID>4568 </input>
<input>
<ID>IN_1</ID>4577 </input>
<output>
<ID>OUT</ID>4511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6142</ID>
<type>BA_TRI_STATE</type>
<position>226,-1600</position>
<input>
<ID>ENABLE_0</ID>4415 </input>
<input>
<ID>IN_0</ID>4413 </input>
<output>
<ID>OUT_0</ID>4461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6143</ID>
<type>AE_DFF_LOW</type>
<position>51,-1631</position>
<input>
<ID>IN_0</ID>4552 </input>
<output>
<ID>OUT_0</ID>4502 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6144</ID>
<type>AA_AND2</type>
<position>23.5,-1572</position>
<input>
<ID>IN_0</ID>4468 </input>
<input>
<ID>IN_1</ID>4470 </input>
<output>
<ID>OUT</ID>4424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6145</ID>
<type>BA_TRI_STATE</type>
<position>61,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4502 </input>
<output>
<ID>OUT_0</ID>4553 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6146</ID>
<type>AA_AND2</type>
<position>34.5,-1581.5</position>
<input>
<ID>IN_0</ID>4468 </input>
<input>
<ID>IN_1</ID>4471 </input>
<output>
<ID>OUT</ID>4425 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6147</ID>
<type>AE_DFF_LOW</type>
<position>74,-1631</position>
<input>
<ID>IN_0</ID>4554 </input>
<output>
<ID>OUT_0</ID>4503 </output>
<input>
<ID>clock</ID>4510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6148</ID>
<type>AE_DFF_LOW</type>
<position>51,-1571</position>
<input>
<ID>IN_0</ID>4446 </input>
<output>
<ID>OUT_0</ID>4416 </output>
<input>
<ID>clock</ID>4424 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6149</ID>
<type>BA_TRI_STATE</type>
<position>84,-1641.5</position>
<input>
<ID>ENABLE_0</ID>4511 </input>
<input>
<ID>IN_0</ID>4503 </input>
<output>
<ID>OUT_0</ID>4555 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6150</ID>
<type>BA_TRI_STATE</type>
<position>61,-1581.5</position>
<input>
<ID>ENABLE_0</ID>4425 </input>
<input>
<ID>IN_0</ID>4416 </input>
<output>
<ID>OUT_0</ID>4447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3761.5,81,-3761.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3761.5,75,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3746,75,-3746</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3761.5,104,-3761.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3761.5,98,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3746,98,-3746</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3761.5,129,-3761.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3761.5,123,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3746,123,-3746</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3761.5,152,-3761.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3761.5,146,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3746,146,-3746</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3761.5,175,-3761.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3761.5,169,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3746,169,-3746</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3761.5,198,-3761.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3761.5,192,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3746,192,-3746</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3761.5,223,-3761.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3761.5,217,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3746,217,-3746</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3761.5,246,-3761.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3761.5,240,-3746</points>
<intersection>-3761.5 1</intersection>
<intersection>-3746 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3746,240,-3746</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3749,233,-3749</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>190</GID>
<name>clock</name></connection>
<connection>
<GID>212</GID>
<name>clock</name></connection>
<connection>
<GID>216</GID>
<name>clock</name></connection>
<connection>
<GID>220</GID>
<name>clock</name></connection>
<connection>
<GID>224</GID>
<name>clock</name></connection>
<connection>
<GID>228</GID>
<name>clock</name></connection>
<connection>
<GID>232</GID>
<name>clock</name></connection>
<connection>
<GID>236</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3758.5,244,-3758.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<connection>
<GID>196</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>214</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>218</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>222</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>226</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>230</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>234</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>238</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3743,81,-3743</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3743,75,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3727.5,75,-3727.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3743,104,-3743</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3743,98,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3727.5,98,-3727.5</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3743,129,-3743</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3743,123,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3727.5,123,-3727.5</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3743,152,-3743</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3743,146,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3727.5,146,-3727.5</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3743,175,-3743</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3743,169,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3727.5,169,-3727.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3743,198,-3743</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3743,192,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3727.5,192,-3727.5</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3743,223,-3743</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3743,217,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3727.5,217,-3727.5</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3743,246,-3743</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3743,240,-3727.5</points>
<intersection>-3743 1</intersection>
<intersection>-3727.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3727.5,240,-3727.5</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3730.5,233,-3730.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<connection>
<GID>244</GID>
<name>clock</name></connection>
<connection>
<GID>248</GID>
<name>clock</name></connection>
<connection>
<GID>252</GID>
<name>clock</name></connection>
<connection>
<GID>256</GID>
<name>clock</name></connection>
<connection>
<GID>260</GID>
<name>clock</name></connection>
<connection>
<GID>264</GID>
<name>clock</name></connection>
<connection>
<GID>268</GID>
<name>clock</name></connection>
<connection>
<GID>272</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3740,244,-3740</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<connection>
<GID>246</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>250</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>254</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>258</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>262</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>266</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>270</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>274</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3724,81,-3724</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3724,75,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3708.5,75,-3708.5</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3724,104,-3724</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3724,98,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3708.5,98,-3708.5</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3724,129,-3724</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3724,123,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3708.5,123,-3708.5</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3724,152,-3724</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3724,146,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3708.5,146,-3708.5</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3724,175,-3724</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3724,169,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3708.5,169,-3708.5</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3724,198,-3724</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3724,192,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3708.5,192,-3708.5</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3724,223,-3724</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3724,217,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3708.5,217,-3708.5</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3724,246,-3724</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3724,240,-3708.5</points>
<intersection>-3724 1</intersection>
<intersection>-3708.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3708.5,240,-3708.5</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3711.5,233,-3711.5</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<connection>
<GID>280</GID>
<name>clock</name></connection>
<connection>
<GID>284</GID>
<name>clock</name></connection>
<connection>
<GID>288</GID>
<name>clock</name></connection>
<connection>
<GID>292</GID>
<name>clock</name></connection>
<connection>
<GID>296</GID>
<name>clock</name></connection>
<connection>
<GID>300</GID>
<name>clock</name></connection>
<connection>
<GID>304</GID>
<name>clock</name></connection>
<connection>
<GID>308</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3721,244,-3721</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<connection>
<GID>282</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>286</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>290</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>294</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>298</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>302</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>306</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>310</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3705.5,81,-3705.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3705.5,75,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3690,75,-3690</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3705.5,104,-3705.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3705.5,98,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3690,98,-3690</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3705.5,129,-3705.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3705.5,123,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3690,123,-3690</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3705.5,152,-3705.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3705.5,146,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3690,146,-3690</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3705.5,175,-3705.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3705.5,169,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3690,169,-3690</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3705.5,198,-3705.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3705.5,192,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3690,192,-3690</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3705.5,223,-3705.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3705.5,217,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3690,217,-3690</points>
<connection>
<GID>340</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3705.5,246,-3705.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3705.5,240,-3690</points>
<intersection>-3705.5 1</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3690,240,-3690</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3693,233,-3693</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<connection>
<GID>316</GID>
<name>clock</name></connection>
<connection>
<GID>320</GID>
<name>clock</name></connection>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<connection>
<GID>328</GID>
<name>clock</name></connection>
<connection>
<GID>332</GID>
<name>clock</name></connection>
<connection>
<GID>336</GID>
<name>clock</name></connection>
<connection>
<GID>340</GID>
<name>clock</name></connection>
<connection>
<GID>344</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3702.5,244,-3702.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<connection>
<GID>318</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>322</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>326</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>330</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>334</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>338</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>342</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>346</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3839.5,81,-3839.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3839.5,75,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3824,75,-3824</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3839.5,104,-3839.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3839.5,98,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3824,98,-3824</points>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3839.5,129,-3839.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3839.5,123,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3824,123,-3824</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3839.5,152,-3839.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3839.5,146,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3824,146,-3824</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3839.5,175,-3839.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3839.5,169,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3824,169,-3824</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3839.5,198,-3839.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3839.5,192,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3824,192,-3824</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3839.5,223,-3839.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3839.5,217,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3824,217,-3824</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3839.5,246,-3839.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3839.5,240,-3824</points>
<intersection>-3839.5 1</intersection>
<intersection>-3824 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3824,240,-3824</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3827,233,-3827</points>
<connection>
<GID>360</GID>
<name>clock</name></connection>
<connection>
<GID>356</GID>
<name>clock</name></connection>
<connection>
<GID>352</GID>
<name>clock</name></connection>
<connection>
<GID>348</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>clock</name></connection>
<connection>
<GID>13</GID>
<name>clock</name></connection>
<connection>
<GID>9</GID>
<name>clock</name></connection>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<connection>
<GID>1</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3836.5,244,-3836.5</points>
<connection>
<GID>362</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>358</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>354</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<connection>
<GID>19</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>15</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>11</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3821,81,-3821</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3821,75,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3805.5,75,-3805.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3821,104,-3821</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3821,98,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3805.5,98,-3805.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3821,129,-3821</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3821,123,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3805.5,123,-3805.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3821,152,-3821</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3821,146,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3805.5,146,-3805.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3821,175,-3821</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3821,169,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3805.5,169,-3805.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3821,198,-3821</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3821,192,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3805.5,192,-3805.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3821,223,-3821</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3821,217,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3805.5,217,-3805.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3821,246,-3821</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3821,240,-3805.5</points>
<intersection>-3821 1</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3805.5,240,-3805.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3808.5,233,-3808.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<connection>
<GID>41</GID>
<name>clock</name></connection>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<connection>
<GID>49</GID>
<name>clock</name></connection>
<connection>
<GID>53</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3818,244,-3818</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>31</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>35</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>39</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>43</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>47</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>51</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>55</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3802,81,-3802</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3802,75,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3786.5,75,-3786.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3802,104,-3802</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3802,98,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3786.5,98,-3786.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3802,129,-3802</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3802,123,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3786.5,123,-3786.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3802,152,-3802</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3802,146,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3786.5,146,-3786.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3802,175,-3802</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3802,169,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3786.5,169,-3786.5</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3802,198,-3802</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3802,192,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3786.5,192,-3786.5</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3802,223,-3802</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3802,217,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3786.5,217,-3786.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3802,246,-3802</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3802,240,-3786.5</points>
<intersection>-3802 1</intersection>
<intersection>-3786.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3786.5,240,-3786.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3789.5,233,-3789.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<connection>
<GID>73</GID>
<name>clock</name></connection>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<connection>
<GID>83</GID>
<name>clock</name></connection>
<connection>
<GID>87</GID>
<name>clock</name></connection>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<connection>
<GID>92</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3799,244,-3799</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<connection>
<GID>65</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>70</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>75</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>80</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>85</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>88</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>91</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>93</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3783.5,81,-3783.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3783.5,75,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3768,75,-3768</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3783.5,104,-3783.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3783.5,98,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3768,98,-3768</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3783.5,129,-3783.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3783.5,123,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3768,123,-3768</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3783.5,152,-3783.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3783.5,146,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3768,146,-3768</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3783.5,175,-3783.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3783.5,169,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3768,169,-3768</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3783.5,198,-3783.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3783.5,192,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3768,192,-3768</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3783.5,223,-3783.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3783.5,217,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3768,217,-3768</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3783.5,246,-3783.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3783.5,240,-3768</points>
<intersection>-3783.5 1</intersection>
<intersection>-3768 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3768,240,-3768</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-241,185,-241</points>
<connection>
<GID>2208</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-241,179,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-225.5,179,-225.5</points>
<connection>
<GID>2207</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3771,233,-3771</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<connection>
<GID>98</GID>
<name>clock</name></connection>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<connection>
<GID>102</GID>
<name>clock</name></connection>
<connection>
<GID>104</GID>
<name>clock</name></connection>
<connection>
<GID>106</GID>
<name>clock</name></connection>
<connection>
<GID>108</GID>
<name>clock</name></connection>
<connection>
<GID>110</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-241,210,-241</points>
<connection>
<GID>2210</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-241,204,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-225.5,204,-225.5</points>
<connection>
<GID>2209</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3780.5,244,-3780.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<connection>
<GID>97</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>99</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>101</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>103</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>105</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>107</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>109</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>111</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-241,233,-241</points>
<connection>
<GID>4159</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-241,227,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-225.5,227,-225.5</points>
<connection>
<GID>4158</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-3849.5,62.5,-3684.5</points>
<connection>
<GID>127</GID>
<name>N_in1</name></connection>
<connection>
<GID>112</GID>
<name>N_in0</name></connection>
<intersection>-3824 12</intersection>
<intersection>-3805.5 11</intersection>
<intersection>-3786.5 10</intersection>
<intersection>-3768 9</intersection>
<intersection>-3746 8</intersection>
<intersection>-3727.5 7</intersection>
<intersection>-3708.5 6</intersection>
<intersection>-3690 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-3690,68,-3690</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>62.5,-3708.5,68,-3708.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>62.5,-3727.5,68,-3727.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>62.5,-3746,68,-3746</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>62.5,-3768,68,-3768</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>62.5,-3786.5,68,-3786.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>62.5,-3805.5,68,-3805.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>62.5,-3824,68,-3824</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-228.5,220,-228.5</points>
<connection>
<GID>4158</GID>
<name>clock</name></connection>
<connection>
<GID>2209</GID>
<name>clock</name></connection>
<connection>
<GID>2207</GID>
<name>clock</name></connection>
<connection>
<GID>2205</GID>
<name>clock</name></connection>
<connection>
<GID>1687</GID>
<name>OUT</name></connection>
<connection>
<GID>1969</GID>
<name>clock</name></connection>
<connection>
<GID>1965</GID>
<name>clock</name></connection>
<connection>
<GID>1961</GID>
<name>clock</name></connection>
<connection>
<GID>1957</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-3849,85.5,-3684</points>
<connection>
<GID>128</GID>
<name>N_in1</name></connection>
<connection>
<GID>113</GID>
<name>N_in0</name></connection>
<intersection>-3833 4</intersection>
<intersection>-3814.5 5</intersection>
<intersection>-3795.5 6</intersection>
<intersection>-3777 7</intersection>
<intersection>-3755 8</intersection>
<intersection>-3736.5 9</intersection>
<intersection>-3717.5 10</intersection>
<intersection>-3699 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>81,-3833,85.5,-3833</points>
<intersection>81 12</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>81,-3814.5,85.5,-3814.5</points>
<intersection>81 13</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>81,-3795.5,85.5,-3795.5</points>
<intersection>81 14</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>81,-3777,85.5,-3777</points>
<intersection>81 15</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>81,-3755,85.5,-3755</points>
<intersection>81 18</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>81,-3736.5,85.5,-3736.5</points>
<intersection>81 19</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>81,-3717.5,85.5,-3717.5</points>
<intersection>81 20</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>81,-3699,85.5,-3699</points>
<intersection>81 21</intersection>
<intersection>85.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>81,-3834,81,-3833</points>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<intersection>-3833 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>81,-3815.5,81,-3814.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>81,-3796.5,81,-3795.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>81,-3778,81,-3777</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-3777 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>81,-3756,81,-3755</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-3755 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>81,-3737.5,81,-3736.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>81,-3718.5,81,-3717.5</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>81,-3700,81,-3699</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>-3699 11</intersection></vsegment></shape></wire>
<wire>
<ID>3161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-238,231,-238</points>
<connection>
<GID>4159</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>2210</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>2208</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>2206</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>2204</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1967</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1963</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1959</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1955</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-3849,88.5,-3684.5</points>
<connection>
<GID>129</GID>
<name>N_in1</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection>
<intersection>-3824 10</intersection>
<intersection>-3805.5 9</intersection>
<intersection>-3786.5 8</intersection>
<intersection>-3768 7</intersection>
<intersection>-3746 6</intersection>
<intersection>-3727.5 5</intersection>
<intersection>-3708.5 4</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-3690,91,-3690</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>88.5,-3708.5,91,-3708.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>88.5,-3727.5,91,-3727.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>88.5,-3746,91,-3746</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>88.5,-3768,91,-3768</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>88.5,-3786.5,91,-3786.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>88.5,-3805.5,91,-3805.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>88.5,-3824,91,-3824</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-222.5,68,-222.5</points>
<connection>
<GID>4163</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-222.5,62,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-207,62,-207</points>
<connection>
<GID>4162</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-3849,108,-3684</points>
<connection>
<GID>130</GID>
<name>N_in1</name></connection>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>-3833 6</intersection>
<intersection>-3814.5 7</intersection>
<intersection>-3795.5 8</intersection>
<intersection>-3777 9</intersection>
<intersection>-3755 10</intersection>
<intersection>-3736.5 11</intersection>
<intersection>-3717.5 12</intersection>
<intersection>-3699 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>104,-3833,108,-3833</points>
<intersection>104 14</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>104,-3814.5,108,-3814.5</points>
<intersection>104 15</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>104,-3795.5,108,-3795.5</points>
<intersection>104 16</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>104,-3777,108,-3777</points>
<intersection>104 17</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>104,-3755,108,-3755</points>
<intersection>104 20</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>104,-3736.5,108,-3736.5</points>
<intersection>104 21</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>104,-3717.5,108,-3717.5</points>
<intersection>104 22</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>104,-3699,108,-3699</points>
<intersection>104 23</intersection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>104,-3834,104,-3833</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-3833 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>104,-3815.5,104,-3814.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>104,-3796.5,104,-3795.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>104,-3778,104,-3777</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>-3777 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>104,-3756,104,-3755</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>-3755 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>104,-3737.5,104,-3736.5</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>104,-3718.5,104,-3717.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>104,-3700,104,-3699</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>-3699 13</intersection></vsegment></shape></wire>
<wire>
<ID>3163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-222.5,91,-222.5</points>
<connection>
<GID>4165</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-222.5,85,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-207,85,-207</points>
<connection>
<GID>4164</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-3849,111.5,-3684</points>
<connection>
<GID>131</GID>
<name>N_in1</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<intersection>-3824 13</intersection>
<intersection>-3805.5 12</intersection>
<intersection>-3786.5 11</intersection>
<intersection>-3768 10</intersection>
<intersection>-3746 9</intersection>
<intersection>-3727.5 8</intersection>
<intersection>-3708.5 7</intersection>
<intersection>-3690 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>111.5,-3690,116,-3690</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111.5,-3708.5,116,-3708.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111.5,-3727.5,116,-3727.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111.5,-3746,116,-3746</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111.5,-3768,116,-3768</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>111.5,-3786.5,116,-3786.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>111.5,-3805.5,116,-3805.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111.5,-3824,116,-3824</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-222.5,116,-222.5</points>
<connection>
<GID>4167</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-222.5,110,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-207,110,-207</points>
<connection>
<GID>4166</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-3849,132.5,-3684.5</points>
<connection>
<GID>132</GID>
<name>N_in1</name></connection>
<connection>
<GID>117</GID>
<name>N_in0</name></connection>
<intersection>-3833 6</intersection>
<intersection>-3814.5 7</intersection>
<intersection>-3795.5 8</intersection>
<intersection>-3777 9</intersection>
<intersection>-3755 10</intersection>
<intersection>-3736.5 11</intersection>
<intersection>-3717.5 12</intersection>
<intersection>-3699 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>129,-3833,132.5,-3833</points>
<intersection>129 14</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>129,-3814.5,132.5,-3814.5</points>
<intersection>129 15</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>129,-3795.5,132.5,-3795.5</points>
<intersection>129 16</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>129,-3777,132.5,-3777</points>
<intersection>129 17</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>129,-3755,132.5,-3755</points>
<intersection>129 20</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>129,-3736.5,132.5,-3736.5</points>
<intersection>129 21</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>129,-3717.5,132.5,-3717.5</points>
<intersection>129 22</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>129,-3699,132.5,-3699</points>
<intersection>129 23</intersection>
<intersection>132.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>129,-3834,129,-3833</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<intersection>-3833 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>129,-3815.5,129,-3814.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>129,-3796.5,129,-3795.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>129,-3778,129,-3777</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>-3777 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>129,-3756,129,-3755</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>-3755 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>129,-3737.5,129,-3736.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>129,-3718.5,129,-3717.5</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>129,-3700,129,-3699</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>-3699 13</intersection></vsegment></shape></wire>
<wire>
<ID>3165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-222.5,139,-222.5</points>
<connection>
<GID>4169</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-222.5,133,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-207,133,-207</points>
<connection>
<GID>4168</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-3849,136.5,-3684</points>
<connection>
<GID>133</GID>
<name>N_in1</name></connection>
<connection>
<GID>118</GID>
<name>N_in0</name></connection>
<intersection>-3824 13</intersection>
<intersection>-3805.5 12</intersection>
<intersection>-3786.5 11</intersection>
<intersection>-3768 10</intersection>
<intersection>-3746 9</intersection>
<intersection>-3727.5 8</intersection>
<intersection>-3708.5 7</intersection>
<intersection>-3690 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>136.5,-3690,139,-3690</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>136.5,-3708.5,139,-3708.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>136.5,-3727.5,139,-3727.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>136.5,-3746,139,-3746</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>136.5,-3768,139,-3768</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>136.5,-3786.5,139,-3786.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>136.5,-3805.5,139,-3805.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>136.5,-3824,139,-3824</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-222.5,162,-222.5</points>
<connection>
<GID>4171</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-222.5,156,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-207,156,-207</points>
<connection>
<GID>4170</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-3849,155,-3684</points>
<connection>
<GID>134</GID>
<name>N_in1</name></connection>
<connection>
<GID>119</GID>
<name>N_in0</name></connection>
<intersection>-3833 6</intersection>
<intersection>-3814.5 7</intersection>
<intersection>-3795.5 8</intersection>
<intersection>-3777 9</intersection>
<intersection>-3755 10</intersection>
<intersection>-3736.5 11</intersection>
<intersection>-3717.5 12</intersection>
<intersection>-3699 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>152,-3833,155,-3833</points>
<intersection>152 14</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>152,-3814.5,155,-3814.5</points>
<intersection>152 15</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>152,-3795.5,155,-3795.5</points>
<intersection>152 16</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-3777,155,-3777</points>
<intersection>152 17</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>152,-3755,155,-3755</points>
<intersection>152 20</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>152,-3736.5,155,-3736.5</points>
<intersection>152 21</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>152,-3717.5,155,-3717.5</points>
<intersection>152 22</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>152,-3699,155,-3699</points>
<intersection>152 23</intersection>
<intersection>155 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>152,-3834,152,-3833</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-3833 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>152,-3815.5,152,-3814.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>152,-3796.5,152,-3795.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>152,-3778,152,-3777</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-3777 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>152,-3756,152,-3755</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>-3755 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>152,-3737.5,152,-3736.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>152,-3718.5,152,-3717.5</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>152,-3700,152,-3699</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>-3699 13</intersection></vsegment></shape></wire>
<wire>
<ID>3167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-222.5,185,-222.5</points>
<connection>
<GID>4173</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-222.5,179,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-207,179,-207</points>
<connection>
<GID>4172</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-3849,159,-3684</points>
<connection>
<GID>135</GID>
<name>N_in1</name></connection>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<intersection>-3824 13</intersection>
<intersection>-3805.5 12</intersection>
<intersection>-3786.5 11</intersection>
<intersection>-3768 10</intersection>
<intersection>-3746 9</intersection>
<intersection>-3727.5 8</intersection>
<intersection>-3708.5 7</intersection>
<intersection>-3690 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>159,-3690,162,-3690</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>159,-3708.5,162,-3708.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>159,-3727.5,162,-3727.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>159,-3746,162,-3746</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>159,-3768,162,-3768</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>159,-3786.5,162,-3786.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>159,-3805.5,162,-3805.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>159,-3824,162,-3824</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>3168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-222.5,210,-222.5</points>
<connection>
<GID>4175</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-222.5,204,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-207,204,-207</points>
<connection>
<GID>4174</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-3848.5,178,-3684</points>
<connection>
<GID>136</GID>
<name>N_in1</name></connection>
<connection>
<GID>121</GID>
<name>N_in0</name></connection>
<intersection>-3833 6</intersection>
<intersection>-3814.5 7</intersection>
<intersection>-3795.5 8</intersection>
<intersection>-3777 9</intersection>
<intersection>-3755 10</intersection>
<intersection>-3736.5 11</intersection>
<intersection>-3717.5 12</intersection>
<intersection>-3699 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>175,-3833,178,-3833</points>
<intersection>175 14</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>175,-3814.5,178,-3814.5</points>
<intersection>175 15</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>175,-3795.5,178,-3795.5</points>
<intersection>175 16</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>175,-3777,178,-3777</points>
<intersection>175 17</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>175,-3755,178,-3755</points>
<intersection>175 20</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>175,-3736.5,178,-3736.5</points>
<intersection>175 21</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>175,-3717.5,178,-3717.5</points>
<intersection>175 22</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>175,-3699,178,-3699</points>
<intersection>175 23</intersection>
<intersection>178 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>175,-3834,175,-3833</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-3833 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>175,-3815.5,175,-3814.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>175,-3796.5,175,-3795.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>175,-3778,175,-3777</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>-3777 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>175,-3756,175,-3755</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>-3755 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>175,-3737.5,175,-3736.5</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>175,-3718.5,175,-3717.5</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>175,-3700,175,-3699</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>-3699 13</intersection></vsegment></shape></wire>
<wire>
<ID>3169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-222.5,233,-222.5</points>
<connection>
<GID>4177</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-222.5,227,-207</points>
<intersection>-222.5 1</intersection>
<intersection>-207 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-207,227,-207</points>
<connection>
<GID>4176</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-3848.5,183,-3684</points>
<connection>
<GID>137</GID>
<name>N_in1</name></connection>
<connection>
<GID>122</GID>
<name>N_in0</name></connection>
<intersection>-3824 13</intersection>
<intersection>-3805.5 12</intersection>
<intersection>-3786.5 11</intersection>
<intersection>-3768 10</intersection>
<intersection>-3746 9</intersection>
<intersection>-3727.5 8</intersection>
<intersection>-3708.5 7</intersection>
<intersection>-3690 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>183,-3690,185,-3690</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>183,-3708.5,185,-3708.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>183,-3727.5,185,-3727.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>183,-3746,185,-3746</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183,-3768,185,-3768</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183,-3786.5,185,-3786.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183,-3805.5,185,-3805.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183,-3824,185,-3824</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>3170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-210,220,-210</points>
<connection>
<GID>4176</GID>
<name>clock</name></connection>
<connection>
<GID>4174</GID>
<name>clock</name></connection>
<connection>
<GID>4172</GID>
<name>clock</name></connection>
<connection>
<GID>4170</GID>
<name>clock</name></connection>
<connection>
<GID>4168</GID>
<name>clock</name></connection>
<connection>
<GID>4166</GID>
<name>clock</name></connection>
<connection>
<GID>4164</GID>
<name>clock</name></connection>
<connection>
<GID>4162</GID>
<name>clock</name></connection>
<connection>
<GID>4160</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-3848,201,-3684</points>
<connection>
<GID>138</GID>
<name>N_in1</name></connection>
<connection>
<GID>124</GID>
<name>N_in0</name></connection>
<intersection>-3833 16</intersection>
<intersection>-3814.5 15</intersection>
<intersection>-3795.5 14</intersection>
<intersection>-3777 13</intersection>
<intersection>-3755 12</intersection>
<intersection>-3736.5 11</intersection>
<intersection>-3717.5 10</intersection>
<intersection>-3699 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>198,-3699,201,-3699</points>
<intersection>198 26</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>198,-3717.5,201,-3717.5</points>
<intersection>198 25</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>198,-3736.5,201,-3736.5</points>
<intersection>198 24</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>198,-3755,201,-3755</points>
<intersection>198 23</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>198,-3777,201,-3777</points>
<intersection>198 20</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>198,-3795.5,201,-3795.5</points>
<intersection>198 19</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>198,-3814.5,201,-3814.5</points>
<intersection>198 18</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>198,-3833,201,-3833</points>
<intersection>198 17</intersection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>198,-3834,198,-3833</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-3833 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>198,-3815.5,198,-3814.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>198,-3796.5,198,-3795.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>198,-3778,198,-3777</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>-3777 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>198,-3756,198,-3755</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>-3755 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>198,-3737.5,198,-3736.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>198,-3718.5,198,-3717.5</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>198,-3700,198,-3699</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>-3699 9</intersection></vsegment></shape></wire>
<wire>
<ID>3171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-219.5,231,-219.5</points>
<connection>
<GID>4177</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4175</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4173</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4171</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4169</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4167</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4165</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4163</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4161</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-3848,205.5,-3684</points>
<connection>
<GID>139</GID>
<name>N_in1</name></connection>
<connection>
<GID>123</GID>
<name>N_in0</name></connection>
<intersection>-3824 13</intersection>
<intersection>-3805.5 12</intersection>
<intersection>-3786.5 11</intersection>
<intersection>-3768 10</intersection>
<intersection>-3746 9</intersection>
<intersection>-3727.5 8</intersection>
<intersection>-3708.5 7</intersection>
<intersection>-3690 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>205.5,-3690,210,-3690</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205.5,-3708.5,210,-3708.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>205.5,-3727.5,210,-3727.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>205.5,-3746,210,-3746</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>205.5,-3768,210,-3768</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205.5,-3786.5,210,-3786.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>205.5,-3805.5,210,-3805.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>205.5,-3824,210,-3824</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-288.5,49.5,-123.5</points>
<connection>
<GID>4195</GID>
<name>N_in1</name></connection>
<connection>
<GID>4178</GID>
<name>N_in0</name></connection>
<intersection>-263 12</intersection>
<intersection>-244.5 11</intersection>
<intersection>-225.5 10</intersection>
<intersection>-207 9</intersection>
<intersection>-185 8</intersection>
<intersection>-166.5 7</intersection>
<intersection>-147.5 6</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-129,55,-129</points>
<connection>
<GID>4271</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>49.5,-147.5,55,-147.5</points>
<connection>
<GID>4253</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>49.5,-166.5,55,-166.5</points>
<connection>
<GID>4235</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>49.5,-185,55,-185</points>
<connection>
<GID>4196</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>49.5,-207,55,-207</points>
<connection>
<GID>4162</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>49.5,-225.5,55,-225.5</points>
<connection>
<GID>1957</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>49.5,-244.5,55,-244.5</points>
<connection>
<GID>1671</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>49.5,-263,55,-263</points>
<connection>
<GID>4289</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-3847.5,226.5,-3684.5</points>
<connection>
<GID>140</GID>
<name>N_in1</name></connection>
<connection>
<GID>125</GID>
<name>N_in0</name></connection>
<intersection>-3833 6</intersection>
<intersection>-3814.5 7</intersection>
<intersection>-3795.5 8</intersection>
<intersection>-3777 9</intersection>
<intersection>-3755 10</intersection>
<intersection>-3736.5 11</intersection>
<intersection>-3717.5 12</intersection>
<intersection>-3699 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>223,-3833,226.5,-3833</points>
<intersection>223 14</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>223,-3814.5,226.5,-3814.5</points>
<intersection>223 15</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>223,-3795.5,226.5,-3795.5</points>
<intersection>223 16</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>223,-3777,226.5,-3777</points>
<intersection>223 17</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>223,-3755,226.5,-3755</points>
<intersection>223 20</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>223,-3736.5,226.5,-3736.5</points>
<intersection>223 21</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>223,-3717.5,226.5,-3717.5</points>
<intersection>223 22</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>223,-3699,226.5,-3699</points>
<intersection>223 23</intersection>
<intersection>226.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>223,-3834,223,-3833</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-3833 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>223,-3815.5,223,-3814.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>223,-3796.5,223,-3795.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>223,-3778,223,-3777</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>-3777 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>223,-3756,223,-3755</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>-3755 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>223,-3737.5,223,-3736.5</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>223,-3718.5,223,-3717.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>223,-3700,223,-3699</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-3699 13</intersection></vsegment></shape></wire>
<wire>
<ID>3173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-288,72.5,-123</points>
<connection>
<GID>4197</GID>
<name>N_in1</name></connection>
<connection>
<GID>4179</GID>
<name>N_in0</name></connection>
<intersection>-272.5 4</intersection>
<intersection>-254 5</intersection>
<intersection>-235 6</intersection>
<intersection>-216.5 7</intersection>
<intersection>-194.5 8</intersection>
<intersection>-176 9</intersection>
<intersection>-157 10</intersection>
<intersection>-138.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68,-272.5,72.5,-272.5</points>
<intersection>68 12</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68,-254,72.5,-254</points>
<intersection>68 14</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68,-235,72.5,-235</points>
<intersection>68 13</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68,-216.5,72.5,-216.5</points>
<intersection>68 15</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68,-194.5,72.5,-194.5</points>
<intersection>68 18</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68,-176,72.5,-176</points>
<intersection>68 19</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68,-157,72.5,-157</points>
<intersection>68 20</intersection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>68,-138.5,72.5,-138.5</points>
<intersection>68 21</intersection>
<intersection>72.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>68,-273,68,-272.5</points>
<connection>
<GID>4290</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>68,-235.5,68,-235</points>
<connection>
<GID>1959</GID>
<name>OUT_0</name></connection>
<intersection>-235 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>68,-254.5,68,-254</points>
<connection>
<GID>1672</GID>
<name>OUT_0</name></connection>
<intersection>-254 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>68,-217,68,-216.5</points>
<connection>
<GID>4163</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>68,-195,68,-194.5</points>
<connection>
<GID>4202</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>68,-176.5,68,-176</points>
<connection>
<GID>4236</GID>
<name>OUT_0</name></connection>
<intersection>-176 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>68,-157.5,68,-157</points>
<connection>
<GID>4254</GID>
<name>OUT_0</name></connection>
<intersection>-157 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>68,-139,68,-138.5</points>
<connection>
<GID>4272</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-3847.5,230,-3684.5</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<connection>
<GID>141</GID>
<name>N_in1</name></connection>
<intersection>-3824 11</intersection>
<intersection>-3805.5 10</intersection>
<intersection>-3786.5 9</intersection>
<intersection>-3768 7</intersection>
<intersection>-3746 6</intersection>
<intersection>-3727.5 5</intersection>
<intersection>-3708.5 4</intersection>
<intersection>-3690 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>230,-3690,233,-3690</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>230,-3708.5,233,-3708.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>230,-3727.5,233,-3727.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>230,-3746,233,-3746</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>230,-3768,233,-3768</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>230,-3786.5,233,-3786.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>230,-3805.5,233,-3805.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>230,-3824,233,-3824</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>3174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-288,75.5,-123.5</points>
<connection>
<GID>4198</GID>
<name>N_in1</name></connection>
<connection>
<GID>4180</GID>
<name>N_in0</name></connection>
<intersection>-263 10</intersection>
<intersection>-244.5 9</intersection>
<intersection>-225.5 8</intersection>
<intersection>-207 7</intersection>
<intersection>-185 6</intersection>
<intersection>-166.5 5</intersection>
<intersection>-147.5 4</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-129,78,-129</points>
<connection>
<GID>4273</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>75.5,-147.5,78,-147.5</points>
<connection>
<GID>4255</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>75.5,-166.5,78,-166.5</points>
<connection>
<GID>4237</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>75.5,-185,78,-185</points>
<connection>
<GID>4214</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>75.5,-207,78,-207</points>
<connection>
<GID>4164</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>75.5,-225.5,78,-225.5</points>
<connection>
<GID>1961</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>75.5,-244.5,78,-244.5</points>
<connection>
<GID>1673</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>75.5,-263,78,-263</points>
<connection>
<GID>4291</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-3847.5,251,-3685.5</points>
<connection>
<GID>126</GID>
<name>N_in0</name></connection>
<connection>
<GID>143</GID>
<name>N_in1</name></connection>
<intersection>-3833 11</intersection>
<intersection>-3814.5 10</intersection>
<intersection>-3795.5 9</intersection>
<intersection>-3777 8</intersection>
<intersection>-3755 7</intersection>
<intersection>-3736.5 6</intersection>
<intersection>-3717.5 5</intersection>
<intersection>-3699 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>246,-3699,251,-3699</points>
<intersection>246 21</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>246,-3717.5,251,-3717.5</points>
<intersection>246 20</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>246,-3736.5,251,-3736.5</points>
<intersection>246 19</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>246,-3755,251,-3755</points>
<intersection>246 18</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>246,-3777,251,-3777</points>
<intersection>246 15</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>246,-3795.5,251,-3795.5</points>
<intersection>246 14</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>246,-3814.5,251,-3814.5</points>
<intersection>246 13</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>246,-3833,251,-3833</points>
<intersection>246 12</intersection>
<intersection>251 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>246,-3834,246,-3833</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-3833 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>246,-3815.5,246,-3814.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>-3814.5 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>246,-3796.5,246,-3795.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>-3795.5 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>246,-3778,246,-3777</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>-3777 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>246,-3756,246,-3755</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-3755 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>246,-3737.5,246,-3736.5</points>
<connection>
<GID>274</GID>
<name>OUT_0</name></connection>
<intersection>-3736.5 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>246,-3718.5,246,-3717.5</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>-3717.5 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>246,-3700,246,-3699</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>-3699 4</intersection></vsegment></shape></wire>
<wire>
<ID>3175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-288,95,-123</points>
<connection>
<GID>4199</GID>
<name>N_in1</name></connection>
<connection>
<GID>4181</GID>
<name>N_in0</name></connection>
<intersection>-272.5 6</intersection>
<intersection>-254 7</intersection>
<intersection>-235 8</intersection>
<intersection>-216.5 9</intersection>
<intersection>-194.5 10</intersection>
<intersection>-176 11</intersection>
<intersection>-157 12</intersection>
<intersection>-138.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91,-272.5,95,-272.5</points>
<intersection>91 14</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>91,-254,95,-254</points>
<intersection>91 16</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>91,-235,95,-235</points>
<intersection>91 15</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>91,-216.5,95,-216.5</points>
<intersection>91 17</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>91,-194.5,95,-194.5</points>
<intersection>91 20</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>91,-176,95,-176</points>
<intersection>91 21</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>91,-157,95,-157</points>
<intersection>91 22</intersection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>91,-138.5,95,-138.5</points>
<intersection>91 23</intersection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>91,-273,91,-272.5</points>
<connection>
<GID>4292</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>91,-235.5,91,-235</points>
<connection>
<GID>1963</GID>
<name>OUT_0</name></connection>
<intersection>-235 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>91,-254.5,91,-254</points>
<connection>
<GID>1674</GID>
<name>OUT_0</name></connection>
<intersection>-254 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>91,-217,91,-216.5</points>
<connection>
<GID>4165</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>91,-195,91,-194.5</points>
<connection>
<GID>4215</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>91,-176.5,91,-176</points>
<connection>
<GID>4238</GID>
<name>OUT_0</name></connection>
<intersection>-176 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>91,-157.5,91,-157</points>
<connection>
<GID>4256</GID>
<name>OUT_0</name></connection>
<intersection>-157 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>91,-139,91,-138.5</points>
<connection>
<GID>4274</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-106,-3692,40.5,-3692</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>-106 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-106,-3843.5,-106,-3692</points>
<connection>
<GID>149</GID>
<name>OUT_15</name></connection>
<intersection>-3701.5 4</intersection>
<intersection>-3692 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-106,-3701.5,52,-3701.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>-106 3</intersection></hsegment></shape></wire>
<wire>
<ID>3176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-288,98.5,-123</points>
<connection>
<GID>4200</GID>
<name>N_in1</name></connection>
<connection>
<GID>4182</GID>
<name>N_in0</name></connection>
<intersection>-263 13</intersection>
<intersection>-244.5 12</intersection>
<intersection>-225.5 11</intersection>
<intersection>-207 10</intersection>
<intersection>-185 9</intersection>
<intersection>-166.5 8</intersection>
<intersection>-147.5 7</intersection>
<intersection>-129 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>98.5,-129,103,-129</points>
<connection>
<GID>4275</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>98.5,-147.5,103,-147.5</points>
<connection>
<GID>4257</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>98.5,-166.5,103,-166.5</points>
<connection>
<GID>4239</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>98.5,-185,103,-185</points>
<connection>
<GID>4217</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>98.5,-207,103,-207</points>
<connection>
<GID>4166</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>98.5,-225.5,103,-225.5</points>
<connection>
<GID>1965</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>98.5,-244.5,103,-244.5</points>
<connection>
<GID>1675</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>98.5,-263,103,-263</points>
<connection>
<GID>4293</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-105,-3710.5,40.5,-3710.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>-105 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-105,-3844.5,-105,-3710.5</points>
<intersection>-3844.5 6</intersection>
<intersection>-3720 5</intersection>
<intersection>-3710.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-105,-3720,52,-3720</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>-105 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-106,-3844.5,-105,-3844.5</points>
<connection>
<GID>149</GID>
<name>OUT_14</name></connection>
<intersection>-105 4</intersection></hsegment></shape></wire>
<wire>
<ID>3177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-288,119.5,-123.5</points>
<connection>
<GID>4201</GID>
<name>N_in1</name></connection>
<connection>
<GID>4183</GID>
<name>N_in0</name></connection>
<intersection>-272.5 6</intersection>
<intersection>-254 7</intersection>
<intersection>-235 8</intersection>
<intersection>-216.5 9</intersection>
<intersection>-194.5 10</intersection>
<intersection>-176 11</intersection>
<intersection>-157 12</intersection>
<intersection>-138.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116,-272.5,119.5,-272.5</points>
<intersection>116 14</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116,-254,119.5,-254</points>
<intersection>116 16</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>116,-235,119.5,-235</points>
<intersection>116 15</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116,-216.5,119.5,-216.5</points>
<intersection>116 17</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116,-194.5,119.5,-194.5</points>
<intersection>116 20</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>116,-176,119.5,-176</points>
<intersection>116 21</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>116,-157,119.5,-157</points>
<intersection>116 22</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>116,-138.5,119.5,-138.5</points>
<intersection>116 23</intersection>
<intersection>119.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>116,-273,116,-272.5</points>
<connection>
<GID>4294</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>116,-235.5,116,-235</points>
<connection>
<GID>1967</GID>
<name>OUT_0</name></connection>
<intersection>-235 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>116,-254.5,116,-254</points>
<connection>
<GID>1676</GID>
<name>OUT_0</name></connection>
<intersection>-254 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>116,-217,116,-216.5</points>
<connection>
<GID>4167</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>116,-195,116,-194.5</points>
<connection>
<GID>4219</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>116,-176.5,116,-176</points>
<connection>
<GID>4240</GID>
<name>OUT_0</name></connection>
<intersection>-176 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>116,-157.5,116,-157</points>
<connection>
<GID>4258</GID>
<name>OUT_0</name></connection>
<intersection>-157 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>116,-139,116,-138.5</points>
<connection>
<GID>4276</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-104,-3729.5,40.5,-3729.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-104 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-104,-3845.5,-104,-3729.5</points>
<intersection>-3845.5 6</intersection>
<intersection>-3739 4</intersection>
<intersection>-3729.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-104,-3739,52,-3739</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-104 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-106,-3845.5,-104,-3845.5</points>
<connection>
<GID>149</GID>
<name>OUT_13</name></connection>
<intersection>-104 3</intersection></hsegment></shape></wire>
<wire>
<ID>3178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-288,123.5,-123</points>
<connection>
<GID>4203</GID>
<name>N_in1</name></connection>
<connection>
<GID>4184</GID>
<name>N_in0</name></connection>
<intersection>-263 13</intersection>
<intersection>-244.5 12</intersection>
<intersection>-225.5 11</intersection>
<intersection>-207 10</intersection>
<intersection>-185 9</intersection>
<intersection>-166.5 8</intersection>
<intersection>-147.5 7</intersection>
<intersection>-129 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>123.5,-129,126,-129</points>
<connection>
<GID>4277</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>123.5,-147.5,126,-147.5</points>
<connection>
<GID>4259</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>123.5,-166.5,126,-166.5</points>
<connection>
<GID>4241</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>123.5,-185,126,-185</points>
<connection>
<GID>4221</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>123.5,-207,126,-207</points>
<connection>
<GID>4168</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>123.5,-225.5,126,-225.5</points>
<connection>
<GID>1969</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>123.5,-244.5,126,-244.5</points>
<connection>
<GID>1677</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>123.5,-263,126,-263</points>
<connection>
<GID>4295</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-103,-3748,40.5,-3748</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-103 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-103,-3846.5,-103,-3748</points>
<intersection>-3846.5 5</intersection>
<intersection>-3757.5 4</intersection>
<intersection>-3748 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-103,-3757.5,52,-3757.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-103 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3846.5,-103,-3846.5</points>
<connection>
<GID>149</GID>
<name>OUT_12</name></connection>
<intersection>-103 3</intersection></hsegment></shape></wire>
<wire>
<ID>3179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-288,142,-123</points>
<connection>
<GID>4204</GID>
<name>N_in1</name></connection>
<connection>
<GID>4185</GID>
<name>N_in0</name></connection>
<intersection>-272.5 6</intersection>
<intersection>-254 7</intersection>
<intersection>-235 8</intersection>
<intersection>-216.5 9</intersection>
<intersection>-194.5 10</intersection>
<intersection>-176 11</intersection>
<intersection>-157 12</intersection>
<intersection>-138.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-272.5,142,-272.5</points>
<intersection>139 14</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,-254,142,-254</points>
<intersection>139 15</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>139,-235,142,-235</points>
<intersection>139 16</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>139,-216.5,142,-216.5</points>
<intersection>139 17</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>139,-194.5,142,-194.5</points>
<intersection>139 20</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139,-176,142,-176</points>
<intersection>139 21</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>139,-157,142,-157</points>
<intersection>139 22</intersection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>139,-138.5,142,-138.5</points>
<intersection>139 23</intersection>
<intersection>142 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>139,-273,139,-272.5</points>
<connection>
<GID>4296</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>139,-254.5,139,-254</points>
<connection>
<GID>1678</GID>
<name>OUT_0</name></connection>
<intersection>-254 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>139,-235.5,139,-235</points>
<connection>
<GID>2204</GID>
<name>OUT_0</name></connection>
<intersection>-235 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>139,-217,139,-216.5</points>
<connection>
<GID>4169</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>139,-195,139,-194.5</points>
<connection>
<GID>4223</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>139,-176.5,139,-176</points>
<connection>
<GID>4242</GID>
<name>OUT_0</name></connection>
<intersection>-176 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>139,-157.5,139,-157</points>
<connection>
<GID>4260</GID>
<name>OUT_0</name></connection>
<intersection>-157 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>139,-139,139,-138.5</points>
<connection>
<GID>4278</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-102,-3770,40.5,-3770</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-102 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-102,-3847.5,-102,-3770</points>
<intersection>-3847.5 6</intersection>
<intersection>-3779.5 4</intersection>
<intersection>-3770 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-102,-3779.5,51.5,-3779.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-102 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-106,-3847.5,-102,-3847.5</points>
<connection>
<GID>149</GID>
<name>OUT_11</name></connection>
<intersection>-102 3</intersection></hsegment></shape></wire>
<wire>
<ID>3180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-288,146,-123</points>
<connection>
<GID>4205</GID>
<name>N_in1</name></connection>
<connection>
<GID>4186</GID>
<name>N_in0</name></connection>
<intersection>-263 13</intersection>
<intersection>-244.5 12</intersection>
<intersection>-225.5 11</intersection>
<intersection>-207 10</intersection>
<intersection>-185 9</intersection>
<intersection>-166.5 8</intersection>
<intersection>-147.5 7</intersection>
<intersection>-129 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>146,-129,149,-129</points>
<connection>
<GID>4279</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>146,-147.5,149,-147.5</points>
<connection>
<GID>4261</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>146,-166.5,149,-166.5</points>
<connection>
<GID>4243</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>146,-185,149,-185</points>
<connection>
<GID>4224</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>146,-207,149,-207</points>
<connection>
<GID>4170</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>146,-225.5,149,-225.5</points>
<connection>
<GID>2205</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>146,-244.5,149,-244.5</points>
<connection>
<GID>1679</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>146,-263,149,-263</points>
<connection>
<GID>4297</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101,-3788.5,40.5,-3788.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-101 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-101,-3848.5,-101,-3788.5</points>
<intersection>-3848.5 5</intersection>
<intersection>-3798 4</intersection>
<intersection>-3788.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-101,-3798,51.5,-3798</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-101 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3848.5,-101,-3848.5</points>
<connection>
<GID>149</GID>
<name>OUT_10</name></connection>
<intersection>-101 3</intersection></hsegment></shape></wire>
<wire>
<ID>3181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-287.5,165,-123</points>
<connection>
<GID>4206</GID>
<name>N_in1</name></connection>
<connection>
<GID>4187</GID>
<name>N_in0</name></connection>
<intersection>-272.5 6</intersection>
<intersection>-254 7</intersection>
<intersection>-235 8</intersection>
<intersection>-216.5 9</intersection>
<intersection>-194.5 10</intersection>
<intersection>-176 11</intersection>
<intersection>-157 12</intersection>
<intersection>-138.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>162,-272.5,165,-272.5</points>
<intersection>162 15</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162,-254,165,-254</points>
<intersection>162 16</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>162,-235,165,-235</points>
<intersection>162 17</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162,-216.5,165,-216.5</points>
<intersection>162 18</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>162,-194.5,165,-194.5</points>
<intersection>162 21</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>162,-176,165,-176</points>
<intersection>162 22</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>162,-157,165,-157</points>
<intersection>162 23</intersection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>162,-138.5,165,-138.5</points>
<intersection>162 14</intersection>
<intersection>165 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>162,-139,162,-138.5</points>
<connection>
<GID>4280</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>162,-273,162,-272.5</points>
<connection>
<GID>4298</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>162,-254.5,162,-254</points>
<connection>
<GID>1680</GID>
<name>OUT_0</name></connection>
<intersection>-254 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>162,-235.5,162,-235</points>
<connection>
<GID>2206</GID>
<name>OUT_0</name></connection>
<intersection>-235 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>162,-217,162,-216.5</points>
<connection>
<GID>4171</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>162,-195,162,-194.5</points>
<connection>
<GID>4226</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>162,-176.5,162,-176</points>
<connection>
<GID>4244</GID>
<name>OUT_0</name></connection>
<intersection>-176 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>162,-157.5,162,-157</points>
<connection>
<GID>4262</GID>
<name>OUT_0</name></connection>
<intersection>-157 12</intersection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100,-3807.5,40.5,-3807.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-100 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-100,-3849.5,-100,-3807.5</points>
<intersection>-3849.5 5</intersection>
<intersection>-3817 4</intersection>
<intersection>-3807.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-100,-3817,51.5,-3817</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-100 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3849.5,-100,-3849.5</points>
<connection>
<GID>149</GID>
<name>OUT_9</name></connection>
<intersection>-100 3</intersection></hsegment></shape></wire>
<wire>
<ID>3182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-287.5,170,-123</points>
<connection>
<GID>4207</GID>
<name>N_in1</name></connection>
<connection>
<GID>4188</GID>
<name>N_in0</name></connection>
<intersection>-263 13</intersection>
<intersection>-244.5 12</intersection>
<intersection>-225.5 11</intersection>
<intersection>-207 10</intersection>
<intersection>-185 9</intersection>
<intersection>-166.5 8</intersection>
<intersection>-147.5 7</intersection>
<intersection>-129 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>170,-129,172,-129</points>
<connection>
<GID>4281</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>170,-147.5,172,-147.5</points>
<connection>
<GID>4263</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>170,-166.5,172,-166.5</points>
<connection>
<GID>4245</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>170,-185,172,-185</points>
<connection>
<GID>4227</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>170,-207,172,-207</points>
<connection>
<GID>4172</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>170,-225.5,172,-225.5</points>
<connection>
<GID>2207</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>170,-244.5,172,-244.5</points>
<connection>
<GID>1681</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>170,-263,172,-263</points>
<connection>
<GID>4299</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-99,-3826,40.5,-3826</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-99 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-99,-3850.5,-99,-3826</points>
<intersection>-3850.5 5</intersection>
<intersection>-3835.5 4</intersection>
<intersection>-3826 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-99,-3835.5,51.5,-3835.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>-99 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3850.5,-99,-3850.5</points>
<connection>
<GID>149</GID>
<name>OUT_8</name></connection>
<intersection>-99 3</intersection></hsegment></shape></wire>
<wire>
<ID>3183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-287,188,-123</points>
<connection>
<GID>4208</GID>
<name>N_in1</name></connection>
<connection>
<GID>4190</GID>
<name>N_in0</name></connection>
<intersection>-272.5 16</intersection>
<intersection>-254 15</intersection>
<intersection>-235 14</intersection>
<intersection>-216.5 13</intersection>
<intersection>-194.5 12</intersection>
<intersection>-176 11</intersection>
<intersection>-157 10</intersection>
<intersection>-138.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>185,-138.5,188,-138.5</points>
<intersection>185 17</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>185,-157,188,-157</points>
<intersection>185 26</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>185,-176,188,-176</points>
<intersection>185 25</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185,-194.5,188,-194.5</points>
<intersection>185 24</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>185,-216.5,188,-216.5</points>
<intersection>185 21</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>185,-235,188,-235</points>
<intersection>185 20</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>185,-254,188,-254</points>
<intersection>185 19</intersection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>185,-272.5,188,-272.5</points>
<intersection>185 18</intersection>
<intersection>188 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>185,-139,185,-138.5</points>
<connection>
<GID>4282</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>185,-273,185,-272.5</points>
<connection>
<GID>4300</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>185,-254.5,185,-254</points>
<connection>
<GID>1682</GID>
<name>OUT_0</name></connection>
<intersection>-254 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>185,-235.5,185,-235</points>
<connection>
<GID>2208</GID>
<name>OUT_0</name></connection>
<intersection>-235 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>185,-217,185,-216.5</points>
<connection>
<GID>4173</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>185,-195,185,-194.5</points>
<connection>
<GID>4228</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>185,-176.5,185,-176</points>
<connection>
<GID>4246</GID>
<name>OUT_0</name></connection>
<intersection>-176 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>185,-157.5,185,-157</points>
<connection>
<GID>4264</GID>
<name>OUT_0</name></connection>
<intersection>-157 10</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-3849.5,39.5,-3684.5</points>
<connection>
<GID>147</GID>
<name>N_in1</name></connection>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<intersection>-3828 10</intersection>
<intersection>-3809.5 9</intersection>
<intersection>-3790.5 8</intersection>
<intersection>-3772 7</intersection>
<intersection>-3750 6</intersection>
<intersection>-3731.5 5</intersection>
<intersection>-3712.5 4</intersection>
<intersection>-3694 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>39.5,-3694,40.5,-3694</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39.5,-3712.5,40.5,-3712.5</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>39.5,-3731.5,40.5,-3731.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>39.5,-3750,40.5,-3750</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>39.5,-3772,40.5,-3772</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>39.5,-3790.5,40.5,-3790.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>39.5,-3809.5,40.5,-3809.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>39.5,-3828,40.5,-3828</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-287,192.5,-123</points>
<connection>
<GID>4209</GID>
<name>N_in1</name></connection>
<connection>
<GID>4189</GID>
<name>N_in0</name></connection>
<intersection>-263 13</intersection>
<intersection>-244.5 12</intersection>
<intersection>-225.5 11</intersection>
<intersection>-207 10</intersection>
<intersection>-185 9</intersection>
<intersection>-166.5 8</intersection>
<intersection>-147.5 7</intersection>
<intersection>-129 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>192.5,-129,197,-129</points>
<connection>
<GID>4283</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>192.5,-147.5,197,-147.5</points>
<connection>
<GID>4265</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>192.5,-166.5,197,-166.5</points>
<connection>
<GID>4247</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>192.5,-185,197,-185</points>
<connection>
<GID>4229</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>192.5,-207,197,-207</points>
<connection>
<GID>4174</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>192.5,-225.5,197,-225.5</points>
<connection>
<GID>2209</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>192.5,-244.5,197,-244.5</points>
<connection>
<GID>1683</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>192.5,-263,197,-263</points>
<connection>
<GID>1665</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-3849.5,49.5,-3684.5</points>
<connection>
<GID>146</GID>
<name>N_in1</name></connection>
<connection>
<GID>144</GID>
<name>N_in0</name></connection>
<intersection>-3837.5 3</intersection>
<intersection>-3819 5</intersection>
<intersection>-3800 7</intersection>
<intersection>-3781.5 9</intersection>
<intersection>-3759.5 11</intersection>
<intersection>-3741 13</intersection>
<intersection>-3722 15</intersection>
<intersection>-3703.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49.5,-3837.5,51.5,-3837.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>49.5,-3819,51.5,-3819</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>49.5,-3800,51.5,-3800</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>49.5,-3781.5,51.5,-3781.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>49.5,-3759.5,52,-3759.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>49.5,-3741,52,-3741</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>49.5,-3722,52,-3722</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>49.5,-3703.5,52,-3703.5</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-286.5,213.5,-123.5</points>
<connection>
<GID>4210</GID>
<name>N_in1</name></connection>
<connection>
<GID>4191</GID>
<name>N_in0</name></connection>
<intersection>-272.5 6</intersection>
<intersection>-254 7</intersection>
<intersection>-235 8</intersection>
<intersection>-216.5 9</intersection>
<intersection>-194.5 10</intersection>
<intersection>-176 11</intersection>
<intersection>-157 12</intersection>
<intersection>-138.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>210,-272.5,213.5,-272.5</points>
<intersection>210 15</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>210,-254,213.5,-254</points>
<intersection>210 16</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>210,-235,213.5,-235</points>
<intersection>210 17</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>210,-216.5,213.5,-216.5</points>
<intersection>210 18</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210,-194.5,213.5,-194.5</points>
<intersection>210 21</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>210,-176,213.5,-176</points>
<intersection>210 22</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>210,-157,213.5,-157</points>
<intersection>210 23</intersection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>210,-138.5,213.5,-138.5</points>
<intersection>210 14</intersection>
<intersection>213.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>210,-139,210,-138.5</points>
<connection>
<GID>4284</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>210,-273,210,-272.5</points>
<connection>
<GID>1666</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>210,-254.5,210,-254</points>
<connection>
<GID>1684</GID>
<name>OUT_0</name></connection>
<intersection>-254 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>210,-235.5,210,-235</points>
<connection>
<GID>2210</GID>
<name>OUT_0</name></connection>
<intersection>-235 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>210,-217,210,-216.5</points>
<connection>
<GID>4175</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>210,-195,210,-194.5</points>
<connection>
<GID>4230</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>210,-176.5,210,-176</points>
<connection>
<GID>4248</GID>
<name>OUT_0</name></connection>
<intersection>-176 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>210,-157.5,210,-157</points>
<connection>
<GID>4266</GID>
<name>OUT_0</name></connection>
<intersection>-157 12</intersection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3937,81,-3937</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3937,75,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3921.5,75,-3921.5</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-286.5,217,-123.5</points>
<connection>
<GID>4211</GID>
<name>N_in1</name></connection>
<connection>
<GID>4212</GID>
<name>N_in0</name></connection>
<intersection>-263 11</intersection>
<intersection>-244.5 10</intersection>
<intersection>-225.5 9</intersection>
<intersection>-207 7</intersection>
<intersection>-185 6</intersection>
<intersection>-166.5 5</intersection>
<intersection>-147.5 4</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-129,220,-129</points>
<connection>
<GID>4285</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>217,-147.5,220,-147.5</points>
<connection>
<GID>4267</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,-166.5,220,-166.5</points>
<connection>
<GID>4249</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>217,-185,220,-185</points>
<connection>
<GID>4231</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>217,-207,220,-207</points>
<connection>
<GID>4176</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>217,-225.5,220,-225.5</points>
<connection>
<GID>4158</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>217,-244.5,220,-244.5</points>
<connection>
<GID>1685</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>217,-263,220,-263</points>
<connection>
<GID>1667</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3937,104,-3937</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3937,98,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3921.5,98,-3921.5</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-286.5,238,-124.5</points>
<connection>
<GID>4213</GID>
<name>N_in1</name></connection>
<connection>
<GID>4192</GID>
<name>N_in0</name></connection>
<intersection>-272.5 11</intersection>
<intersection>-254 10</intersection>
<intersection>-235 9</intersection>
<intersection>-216.5 8</intersection>
<intersection>-194.5 7</intersection>
<intersection>-176 6</intersection>
<intersection>-157 5</intersection>
<intersection>-138.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>233,-138.5,238,-138.5</points>
<intersection>233 12</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>233,-157,238,-157</points>
<intersection>233 21</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>233,-176,238,-176</points>
<intersection>233 20</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>233,-194.5,238,-194.5</points>
<intersection>233 19</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>233,-216.5,238,-216.5</points>
<intersection>233 16</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>233,-235,238,-235</points>
<intersection>233 15</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>233,-254,238,-254</points>
<intersection>233 14</intersection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>233,-272.5,238,-272.5</points>
<intersection>233 13</intersection>
<intersection>238 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>233,-139,233,-138.5</points>
<connection>
<GID>4286</GID>
<name>OUT_0</name></connection>
<intersection>-138.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>233,-273,233,-272.5</points>
<connection>
<GID>1668</GID>
<name>OUT_0</name></connection>
<intersection>-272.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>233,-254.5,233,-254</points>
<connection>
<GID>1686</GID>
<name>OUT_0</name></connection>
<intersection>-254 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>233,-235.5,233,-235</points>
<connection>
<GID>4159</GID>
<name>OUT_0</name></connection>
<intersection>-235 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>233,-217,233,-216.5</points>
<connection>
<GID>4177</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>233,-195,233,-194.5</points>
<connection>
<GID>4232</GID>
<name>OUT_0</name></connection>
<intersection>-194.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>233,-176.5,233,-176</points>
<connection>
<GID>4250</GID>
<name>OUT_0</name></connection>
<intersection>-176 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>233,-157.5,233,-157</points>
<connection>
<GID>4268</GID>
<name>OUT_0</name></connection>
<intersection>-157 5</intersection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3937,129,-3937</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3937,123,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3921.5,123,-3921.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3188</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-112,-131,27.5,-131</points>
<connection>
<GID>4269</GID>
<name>IN_0</name></connection>
<intersection>-112 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-112,-140.5,-112,-115</points>
<intersection>-140.5 4</intersection>
<intersection>-131 2</intersection>
<intersection>-115 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-112,-140.5,39,-140.5</points>
<connection>
<GID>4270</GID>
<name>IN_0</name></connection>
<intersection>-112 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119,-115,-112,-115</points>
<connection>
<GID>1664</GID>
<name>OUT_7</name></connection>
<intersection>-112 3</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3937,152,-3937</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3937,146,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3921.5,146,-3921.5</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3189</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-113,-149.5,27.5,-149.5</points>
<connection>
<GID>4251</GID>
<name>IN_0</name></connection>
<intersection>-113 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-113,-159,-113,-116</points>
<intersection>-159 5</intersection>
<intersection>-149.5 2</intersection>
<intersection>-116 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-113,-159,39,-159</points>
<connection>
<GID>4252</GID>
<name>IN_0</name></connection>
<intersection>-113 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119,-116,-113,-116</points>
<connection>
<GID>1664</GID>
<name>OUT_6</name></connection>
<intersection>-113 4</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3937,175,-3937</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3937,169,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3921.5,169,-3921.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3190</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-114,-168.5,27.5,-168.5</points>
<connection>
<GID>4233</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114,-178,-114,-117</points>
<intersection>-178 4</intersection>
<intersection>-168.5 2</intersection>
<intersection>-117 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-114,-178,39,-178</points>
<connection>
<GID>4234</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119,-117,-114,-117</points>
<connection>
<GID>1664</GID>
<name>OUT_5</name></connection>
<intersection>-114 3</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3937,198,-3937</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3937,192,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3921.5,192,-3921.5</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3191</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-115,-187,27.5,-187</points>
<connection>
<GID>4193</GID>
<name>IN_0</name></connection>
<intersection>-115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-115,-196.5,-115,-118</points>
<intersection>-196.5 4</intersection>
<intersection>-187 2</intersection>
<intersection>-118 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-115,-196.5,39,-196.5</points>
<connection>
<GID>4194</GID>
<name>IN_0</name></connection>
<intersection>-115 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-118,-115,-118</points>
<connection>
<GID>1664</GID>
<name>OUT_4</name></connection>
<intersection>-115 3</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3937,223,-3937</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3937,217,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3921.5,217,-3921.5</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,-209,27.5,-209</points>
<connection>
<GID>4160</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-116,-218.5,-116,-119</points>
<intersection>-218.5 4</intersection>
<intersection>-209 1</intersection>
<intersection>-119 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-116,-218.5,38.5,-218.5</points>
<connection>
<GID>4161</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-119,-116,-119</points>
<connection>
<GID>1664</GID>
<name>OUT_3</name></connection>
<intersection>-116 3</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3937,246,-3937</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3937,240,-3921.5</points>
<intersection>-3937 1</intersection>
<intersection>-3921.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3921.5,240,-3921.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-117,-227.5,27.5,-227.5</points>
<connection>
<GID>1687</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-237,-117,-120</points>
<intersection>-237 4</intersection>
<intersection>-227.5 1</intersection>
<intersection>-120 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-237,38.5,-237</points>
<connection>
<GID>1955</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-120,-117,-120</points>
<connection>
<GID>1664</GID>
<name>OUT_2</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3924.5,233,-3924.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<connection>
<GID>233</GID>
<name>clock</name></connection>
<connection>
<GID>269</GID>
<name>clock</name></connection>
<connection>
<GID>275</GID>
<name>clock</name></connection>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<connection>
<GID>289</GID>
<name>clock</name></connection>
<connection>
<GID>295</GID>
<name>clock</name></connection>
<connection>
<GID>299</GID>
<name>clock</name></connection>
<connection>
<GID>303</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118,-246.5,27.5,-246.5</points>
<connection>
<GID>1669</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118,-256,-118,-121</points>
<intersection>-256 4</intersection>
<intersection>-246.5 1</intersection>
<intersection>-121 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118,-256,38.5,-256</points>
<connection>
<GID>1670</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-121,-118,-121</points>
<connection>
<GID>1664</GID>
<name>OUT_1</name></connection>
<intersection>-118 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3934,244,-3934</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<connection>
<GID>245</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>271</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>279</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>287</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>293</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>297</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>301</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>305</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,-265,27.5,-265</points>
<connection>
<GID>4287</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-274.5,-119,-122</points>
<connection>
<GID>1664</GID>
<name>OUT_0</name></connection>
<intersection>-274.5 4</intersection>
<intersection>-265 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-274.5,38.5,-274.5</points>
<connection>
<GID>4288</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3918.5,81,-3918.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3918.5,75,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3903,75,-3903</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-288.5,26.5,-123.5</points>
<connection>
<GID>4222</GID>
<name>N_in1</name></connection>
<connection>
<GID>4218</GID>
<name>N_in0</name></connection>
<intersection>-267 10</intersection>
<intersection>-248.5 9</intersection>
<intersection>-229.5 8</intersection>
<intersection>-211 7</intersection>
<intersection>-189 6</intersection>
<intersection>-170.5 5</intersection>
<intersection>-151.5 4</intersection>
<intersection>-133 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-133,27.5,-133</points>
<connection>
<GID>4269</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-151.5,27.5,-151.5</points>
<connection>
<GID>4251</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-170.5,27.5,-170.5</points>
<connection>
<GID>4233</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>26.5,-189,27.5,-189</points>
<connection>
<GID>4193</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>26.5,-211,27.5,-211</points>
<connection>
<GID>4160</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>26.5,-229.5,27.5,-229.5</points>
<connection>
<GID>1687</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>26.5,-248.5,27.5,-248.5</points>
<connection>
<GID>1669</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>26.5,-267,27.5,-267</points>
<connection>
<GID>4287</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3918.5,104,-3918.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3918.5,98,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3903,98,-3903</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-288.5,36.5,-123.5</points>
<connection>
<GID>4220</GID>
<name>N_in1</name></connection>
<connection>
<GID>4216</GID>
<name>N_in0</name></connection>
<intersection>-276.5 3</intersection>
<intersection>-258 5</intersection>
<intersection>-239 7</intersection>
<intersection>-220.5 9</intersection>
<intersection>-198.5 11</intersection>
<intersection>-180 13</intersection>
<intersection>-161 15</intersection>
<intersection>-142.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-276.5,38.5,-276.5</points>
<connection>
<GID>4288</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>36.5,-258,38.5,-258</points>
<connection>
<GID>1670</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>36.5,-239,38.5,-239</points>
<connection>
<GID>1955</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>36.5,-220.5,38.5,-220.5</points>
<connection>
<GID>4161</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>36.5,-198.5,39,-198.5</points>
<connection>
<GID>4194</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>36.5,-180,39,-180</points>
<connection>
<GID>4234</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>36.5,-161,39,-161</points>
<connection>
<GID>4252</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>36.5,-142.5,39,-142.5</points>
<connection>
<GID>4270</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3918.5,129,-3918.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3918.5,123,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3903,123,-3903</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-121.5,26.5,-115</points>
<connection>
<GID>1660</GID>
<name>N_in0</name></connection>
<connection>
<GID>4218</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3918.5,152,-3918.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3918.5,146,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3903,146,-3903</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-121.5,36.5,-115</points>
<connection>
<GID>1659</GID>
<name>N_in0</name></connection>
<connection>
<GID>4216</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3918.5,175,-3918.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3918.5,169,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3903,169,-3903</points>
<connection>
<GID>327</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-121.5,49.5,-115</points>
<connection>
<GID>1635</GID>
<name>N_in0</name></connection>
<connection>
<GID>4178</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3918.5,198,-3918.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3918.5,192,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3903,192,-3903</points>
<connection>
<GID>331</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-121,72.5,-114.5</points>
<connection>
<GID>1636</GID>
<name>N_in0</name></connection>
<connection>
<GID>4179</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3918.5,223,-3918.5</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3918.5,217,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3903,217,-3903</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-121.5,75.5,-114.5</points>
<connection>
<GID>1637</GID>
<name>N_in0</name></connection>
<connection>
<GID>4180</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3918.5,246,-3918.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3918.5,240,-3903</points>
<intersection>-3918.5 1</intersection>
<intersection>-3903 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3903,240,-3903</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-121,95,-114.5</points>
<connection>
<GID>1638</GID>
<name>N_in0</name></connection>
<connection>
<GID>4181</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3906,233,-3906</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<connection>
<GID>315</GID>
<name>clock</name></connection>
<connection>
<GID>319</GID>
<name>clock</name></connection>
<connection>
<GID>323</GID>
<name>clock</name></connection>
<connection>
<GID>327</GID>
<name>clock</name></connection>
<connection>
<GID>331</GID>
<name>clock</name></connection>
<connection>
<GID>335</GID>
<name>clock</name></connection>
<connection>
<GID>339</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-121,98.5,-114.5</points>
<connection>
<GID>1639</GID>
<name>N_in0</name></connection>
<connection>
<GID>4182</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3915.5,244,-3915.5</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<connection>
<GID>313</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>317</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>321</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>325</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>329</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>333</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>337</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>341</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-121.5,119.5,-114.5</points>
<connection>
<GID>1640</GID>
<name>N_in0</name></connection>
<connection>
<GID>4183</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3899.5,81,-3899.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3899.5,75,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3884,75,-3884</points>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-121,123.5,-114.5</points>
<connection>
<GID>1641</GID>
<name>N_in0</name></connection>
<connection>
<GID>4184</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3899.5,104,-3899.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3899.5,98,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3884,98,-3884</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-121,142,-114.5</points>
<connection>
<GID>1642</GID>
<name>N_in0</name></connection>
<connection>
<GID>4185</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3899.5,129,-3899.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3899.5,123,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3884,123,-3884</points>
<connection>
<GID>355</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-121,146,-114.5</points>
<connection>
<GID>1643</GID>
<name>N_in0</name></connection>
<connection>
<GID>4186</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3899.5,152,-3899.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3899.5,146,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3884,146,-3884</points>
<connection>
<GID>359</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-121,165,-114</points>
<connection>
<GID>1644</GID>
<name>N_in0</name></connection>
<connection>
<GID>4187</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3899.5,175,-3899.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3899.5,169,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3884,169,-3884</points>
<connection>
<GID>363</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-121,170,-114</points>
<connection>
<GID>1645</GID>
<name>N_in0</name></connection>
<connection>
<GID>4188</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3899.5,198,-3899.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3899.5,192,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3884,192,-3884</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-121,188,-113.5</points>
<connection>
<GID>1646</GID>
<name>N_in0</name></connection>
<connection>
<GID>4190</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3899.5,223,-3899.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3899.5,217,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3884,217,-3884</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-121,192.5,-113.5</points>
<connection>
<GID>1647</GID>
<name>N_in0</name></connection>
<connection>
<GID>4189</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3899.5,246,-3899.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3899.5,240,-3884</points>
<intersection>-3899.5 1</intersection>
<intersection>-3884 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3884,240,-3884</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-121.5,213.5,-113</points>
<connection>
<GID>1648</GID>
<name>N_in0</name></connection>
<connection>
<GID>4191</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3887,233,-3887</points>
<connection>
<GID>363</GID>
<name>clock</name></connection>
<connection>
<GID>359</GID>
<name>clock</name></connection>
<connection>
<GID>355</GID>
<name>clock</name></connection>
<connection>
<GID>351</GID>
<name>clock</name></connection>
<connection>
<GID>347</GID>
<name>clock</name></connection>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<connection>
<GID>4</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-121.5,217,-113</points>
<connection>
<GID>1649</GID>
<name>N_in0</name></connection>
<connection>
<GID>4212</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3896.5,244,-3896.5</points>
<connection>
<GID>361</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>357</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>353</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>349</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>10</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-122.5,238,-113</points>
<connection>
<GID>1653</GID>
<name>N_in0</name></connection>
<connection>
<GID>4192</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3881,81,-3881</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3881,75,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3865.5,75,-3865.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-385,68.5,-385</points>
<connection>
<GID>4461</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-385,62.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-369.5,62.5,-369.5</points>
<connection>
<GID>4455</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3881,104,-3881</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3881,98,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3865.5,98,-3865.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-385,91.5,-385</points>
<connection>
<GID>4479</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-385,85.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-369.5,85.5,-369.5</points>
<connection>
<GID>4477</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3881,129,-3881</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3881,123,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3865.5,123,-3865.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-385,116.5,-385</points>
<connection>
<GID>4483</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-385,110.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-369.5,110.5,-369.5</points>
<connection>
<GID>4481</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3881,152,-3881</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3881,146,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3865.5,146,-3865.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-385,139.5,-385</points>
<connection>
<GID>4487</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-385,133.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-369.5,133.5,-369.5</points>
<connection>
<GID>4485</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3881,175,-3881</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3881,169,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3865.5,169,-3865.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-385,162.5,-385</points>
<connection>
<GID>4491</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-385,156.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-369.5,156.5,-369.5</points>
<connection>
<GID>4489</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3881,198,-3881</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3881,192,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3865.5,192,-3865.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-385,185.5,-385</points>
<connection>
<GID>4495</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-385,179.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-369.5,179.5,-369.5</points>
<connection>
<GID>4493</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3881,223,-3881</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3881,217,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3865.5,217,-3865.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-385,210.5,-385</points>
<connection>
<GID>4499</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-385,204.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-369.5,204.5,-369.5</points>
<connection>
<GID>4497</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3881,246,-3881</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3881,240,-3865.5</points>
<intersection>-3881 1</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3865.5,240,-3865.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-385,233.5,-385</points>
<connection>
<GID>4503</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-385,227.5,-369.5</points>
<intersection>-385 1</intersection>
<intersection>-369.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-369.5,227.5,-369.5</points>
<connection>
<GID>4501</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3868.5,233,-3868.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<connection>
<GID>28</GID>
<name>clock</name></connection>
<connection>
<GID>32</GID>
<name>clock</name></connection>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<connection>
<GID>40</GID>
<name>clock</name></connection>
<connection>
<GID>44</GID>
<name>clock</name></connection>
<connection>
<GID>48</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-372.5,220.5,-372.5</points>
<connection>
<GID>4501</GID>
<name>clock</name></connection>
<connection>
<GID>4497</GID>
<name>clock</name></connection>
<connection>
<GID>4493</GID>
<name>clock</name></connection>
<connection>
<GID>4489</GID>
<name>clock</name></connection>
<connection>
<GID>4485</GID>
<name>clock</name></connection>
<connection>
<GID>4481</GID>
<name>clock</name></connection>
<connection>
<GID>4477</GID>
<name>clock</name></connection>
<connection>
<GID>4455</GID>
<name>clock</name></connection>
<connection>
<GID>4445</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-3878,244,-3878</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>22</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>26</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>30</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>34</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>38</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>42</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>46</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>50</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-382,231.5,-382</points>
<connection>
<GID>4503</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4499</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4495</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4491</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4487</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4483</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4479</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4461</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4450</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-4015,81,-4015</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-4015,75,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3999.5,75,-3999.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-366.5,68.5,-366.5</points>
<connection>
<GID>4511</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-366.5,62.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-351,62.5,-351</points>
<connection>
<GID>4509</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-4015,104,-4015</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-4015,98,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3999.5,98,-3999.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-366.5,91.5,-366.5</points>
<connection>
<GID>4515</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-366.5,85.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-351,85.5,-351</points>
<connection>
<GID>4513</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-4015,129,-4015</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-4015,123,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3999.5,123,-3999.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-366.5,116.5,-366.5</points>
<connection>
<GID>4519</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-366.5,110.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-351,110.5,-351</points>
<connection>
<GID>4517</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-4015,152,-4015</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-4015,146,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3999.5,146,-3999.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-366.5,139.5,-366.5</points>
<connection>
<GID>4523</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-366.5,133.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-351,133.5,-351</points>
<connection>
<GID>4521</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-4015,175,-4015</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-4015,169,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3999.5,169,-3999.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-366.5,162.5,-366.5</points>
<connection>
<GID>4527</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-366.5,156.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-351,156.5,-351</points>
<connection>
<GID>4525</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-4015,198,-4015</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-4015,192,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3999.5,192,-3999.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-366.5,185.5,-366.5</points>
<connection>
<GID>4531</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-366.5,179.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-351,179.5,-351</points>
<connection>
<GID>4529</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-4015,223,-4015</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-4015,217,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3999.5,217,-3999.5</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-366.5,210.5,-366.5</points>
<connection>
<GID>4535</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-366.5,204.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-351,204.5,-351</points>
<connection>
<GID>4533</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-4015,246,-4015</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-4015,240,-3999.5</points>
<intersection>-4015 1</intersection>
<intersection>-3999.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3999.5,240,-3999.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-366.5,233.5,-366.5</points>
<connection>
<GID>4539</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-366.5,227.5,-351</points>
<intersection>-366.5 1</intersection>
<intersection>-351 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-351,227.5,-351</points>
<connection>
<GID>4537</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-4002.5,233,-4002.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<connection>
<GID>61</GID>
<name>clock</name></connection>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<connection>
<GID>81</GID>
<name>clock</name></connection>
<connection>
<GID>150</GID>
<name>clock</name></connection>
<connection>
<GID>152</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-354,220.5,-354</points>
<connection>
<GID>4537</GID>
<name>clock</name></connection>
<connection>
<GID>4533</GID>
<name>clock</name></connection>
<connection>
<GID>4529</GID>
<name>clock</name></connection>
<connection>
<GID>4525</GID>
<name>clock</name></connection>
<connection>
<GID>4521</GID>
<name>clock</name></connection>
<connection>
<GID>4517</GID>
<name>clock</name></connection>
<connection>
<GID>4513</GID>
<name>clock</name></connection>
<connection>
<GID>4509</GID>
<name>clock</name></connection>
<connection>
<GID>4505</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-4012,244,-4012</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>64</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>69</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>74</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>79</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>84</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>151</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>153</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-363.5,231.5,-363.5</points>
<connection>
<GID>4539</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4535</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4531</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4527</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4523</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4519</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4515</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4511</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4507</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3996.5,81,-3996.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3996.5,75,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3981,75,-3981</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-347.5,68.5,-347.5</points>
<connection>
<GID>4547</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-347.5,62.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-332,62.5,-332</points>
<connection>
<GID>4545</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3996.5,104,-3996.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3996.5,98,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3981,98,-3981</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-347.5,91.5,-347.5</points>
<connection>
<GID>4551</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-347.5,85.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-332,85.5,-332</points>
<connection>
<GID>4549</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3996.5,129,-3996.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3996.5,123,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3981,123,-3981</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-347.5,116.5,-347.5</points>
<connection>
<GID>4555</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-347.5,110.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-332,110.5,-332</points>
<connection>
<GID>4553</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3996.5,152,-3996.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3996.5,146,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3981,146,-3981</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-347.5,139.5,-347.5</points>
<connection>
<GID>4559</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-347.5,133.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-332,133.5,-332</points>
<connection>
<GID>4557</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3996.5,175,-3996.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3996.5,169,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3981,169,-3981</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-347.5,162.5,-347.5</points>
<connection>
<GID>4563</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-347.5,156.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-332,156.5,-332</points>
<connection>
<GID>4561</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3996.5,198,-3996.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3996.5,192,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3981,192,-3981</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-347.5,185.5,-347.5</points>
<connection>
<GID>4567</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-347.5,179.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-332,179.5,-332</points>
<connection>
<GID>4565</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3996.5,223,-3996.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3996.5,217,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3981,217,-3981</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-347.5,210.5,-347.5</points>
<connection>
<GID>4571</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-347.5,204.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-332,204.5,-332</points>
<connection>
<GID>4569</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3996.5,246,-3996.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3996.5,240,-3981</points>
<intersection>-3996.5 1</intersection>
<intersection>-3981 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3981,240,-3981</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-347.5,233.5,-347.5</points>
<connection>
<GID>4575</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-347.5,227.5,-332</points>
<intersection>-347.5 1</intersection>
<intersection>-332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-332,227.5,-332</points>
<connection>
<GID>4573</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3984,233,-3984</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<connection>
<GID>156</GID>
<name>clock</name></connection>
<connection>
<GID>158</GID>
<name>clock</name></connection>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<connection>
<GID>162</GID>
<name>clock</name></connection>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<connection>
<GID>168</GID>
<name>clock</name></connection>
<connection>
<GID>170</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-335,220.5,-335</points>
<connection>
<GID>4573</GID>
<name>clock</name></connection>
<connection>
<GID>4569</GID>
<name>clock</name></connection>
<connection>
<GID>4565</GID>
<name>clock</name></connection>
<connection>
<GID>4561</GID>
<name>clock</name></connection>
<connection>
<GID>4557</GID>
<name>clock</name></connection>
<connection>
<GID>4553</GID>
<name>clock</name></connection>
<connection>
<GID>4549</GID>
<name>clock</name></connection>
<connection>
<GID>4545</GID>
<name>clock</name></connection>
<connection>
<GID>4541</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3993.5,244,-3993.5</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<connection>
<GID>157</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>159</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>161</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>163</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>165</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>167</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>169</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>171</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-344.5,231.5,-344.5</points>
<connection>
<GID>4575</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4571</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4567</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4563</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4559</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4555</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4551</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4547</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4543</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3977.5,81,-3977.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3977.5,75,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3962,75,-3962</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-329,68.5,-329</points>
<connection>
<GID>4583</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-329,62.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-313.5,62.5,-313.5</points>
<connection>
<GID>4581</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3977.5,104,-3977.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3977.5,98,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3962,98,-3962</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-329,91.5,-329</points>
<connection>
<GID>4587</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-329,85.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-313.5,85.5,-313.5</points>
<connection>
<GID>4585</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3977.5,129,-3977.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3977.5,123,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3962,123,-3962</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-329,116.5,-329</points>
<connection>
<GID>4591</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-329,110.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-313.5,110.5,-313.5</points>
<connection>
<GID>4589</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3977.5,152,-3977.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3977.5,146,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3962,146,-3962</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-329,139.5,-329</points>
<connection>
<GID>4595</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-329,133.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-313.5,133.5,-313.5</points>
<connection>
<GID>4593</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3977.5,175,-3977.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3977.5,169,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3962,169,-3962</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-329,162.5,-329</points>
<connection>
<GID>4599</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-329,156.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-313.5,156.5,-313.5</points>
<connection>
<GID>4597</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3977.5,198,-3977.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3977.5,192,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3962,192,-3962</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-329,185.5,-329</points>
<connection>
<GID>4603</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-329,179.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-313.5,179.5,-313.5</points>
<connection>
<GID>4601</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3977.5,223,-3977.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3977.5,217,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3962,217,-3962</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-329,210.5,-329</points>
<connection>
<GID>4607</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-329,204.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-313.5,204.5,-313.5</points>
<connection>
<GID>4605</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3977.5,246,-3977.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3977.5,240,-3962</points>
<intersection>-3977.5 1</intersection>
<intersection>-3962 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3962,240,-3962</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-329,233.5,-329</points>
<connection>
<GID>4611</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-329,227.5,-313.5</points>
<intersection>-329 1</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-313.5,227.5,-313.5</points>
<connection>
<GID>4609</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3965,233,-3965</points>
<connection>
<GID>181</GID>
<name>clock</name></connection>
<connection>
<GID>178</GID>
<name>clock</name></connection>
<connection>
<GID>176</GID>
<name>clock</name></connection>
<connection>
<GID>174</GID>
<name>clock</name></connection>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>clock</name></connection>
<connection>
<GID>82</GID>
<name>clock</name></connection>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<connection>
<GID>62</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-316.5,220.5,-316.5</points>
<connection>
<GID>4609</GID>
<name>clock</name></connection>
<connection>
<GID>4605</GID>
<name>clock</name></connection>
<connection>
<GID>4601</GID>
<name>clock</name></connection>
<connection>
<GID>4597</GID>
<name>clock</name></connection>
<connection>
<GID>4593</GID>
<name>clock</name></connection>
<connection>
<GID>4589</GID>
<name>clock</name></connection>
<connection>
<GID>4585</GID>
<name>clock</name></connection>
<connection>
<GID>4581</GID>
<name>clock</name></connection>
<connection>
<GID>4577</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3974.5,244,-3974.5</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>77</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>86</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>173</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>175</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>177</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>179</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>182</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-326,231.5,-326</points>
<connection>
<GID>4611</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4607</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4603</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4599</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4595</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4591</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4587</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4583</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4579</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-3959,81,-3959</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-3959,75,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-3943.5,75,-3943.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>3256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-463,68.5,-463</points>
<connection>
<GID>4619</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-463,62.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-447.5,62.5,-447.5</points>
<connection>
<GID>4617</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-3959,104,-3959</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-3959,98,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-3943.5,98,-3943.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>3257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-463,91.5,-463</points>
<connection>
<GID>4623</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-463,85.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-447.5,85.5,-447.5</points>
<connection>
<GID>4621</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-3959,129,-3959</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-3959,123,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-3943.5,123,-3943.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>3258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-463,116.5,-463</points>
<connection>
<GID>4627</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-463,110.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-447.5,110.5,-447.5</points>
<connection>
<GID>4625</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-3959,152,-3959</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>146,-3959,146,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-3943.5,146,-3943.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>146 2</intersection></hsegment></shape></wire>
<wire>
<ID>3259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-463,139.5,-463</points>
<connection>
<GID>4631</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-463,133.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-447.5,133.5,-447.5</points>
<connection>
<GID>4629</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-3959,175,-3959</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>169 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>169,-3959,169,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>168,-3943.5,169,-3943.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>169 2</intersection></hsegment></shape></wire>
<wire>
<ID>3260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-463,162.5,-463</points>
<connection>
<GID>4635</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-463,156.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-447.5,156.5,-447.5</points>
<connection>
<GID>4633</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-3959,198,-3959</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>192 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192,-3959,192,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-3943.5,192,-3943.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>192 2</intersection></hsegment></shape></wire>
<wire>
<ID>3261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-463,185.5,-463</points>
<connection>
<GID>4639</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-463,179.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-447.5,179.5,-447.5</points>
<connection>
<GID>4637</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-3959,223,-3959</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-3959,217,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-3943.5,217,-3943.5</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>3262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-463,210.5,-463</points>
<connection>
<GID>4643</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-463,204.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-447.5,204.5,-447.5</points>
<connection>
<GID>4641</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-3959,246,-3959</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>240 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>240,-3959,240,-3943.5</points>
<intersection>-3959 1</intersection>
<intersection>-3943.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>239,-3943.5,240,-3943.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>240 2</intersection></hsegment></shape></wire>
<wire>
<ID>3263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-463,233.5,-463</points>
<connection>
<GID>4647</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-463,227.5,-447.5</points>
<intersection>-463 1</intersection>
<intersection>-447.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-447.5,227.5,-447.5</points>
<connection>
<GID>4645</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-3946.5,233,-3946.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>clock</name></connection>
<connection>
<GID>188</GID>
<name>clock</name></connection>
<connection>
<GID>191</GID>
<name>clock</name></connection>
<connection>
<GID>193</GID>
<name>clock</name></connection>
<connection>
<GID>195</GID>
<name>clock</name></connection>
<connection>
<GID>198</GID>
<name>clock</name></connection>
<connection>
<GID>200</GID>
<name>clock</name></connection>
<connection>
<GID>202</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-450.5,220.5,-450.5</points>
<connection>
<GID>4613</GID>
<name>OUT</name></connection>
<connection>
<GID>4645</GID>
<name>clock</name></connection>
<connection>
<GID>4641</GID>
<name>clock</name></connection>
<connection>
<GID>4637</GID>
<name>clock</name></connection>
<connection>
<GID>4633</GID>
<name>clock</name></connection>
<connection>
<GID>4629</GID>
<name>clock</name></connection>
<connection>
<GID>4625</GID>
<name>clock</name></connection>
<connection>
<GID>4621</GID>
<name>clock</name></connection>
<connection>
<GID>4617</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-3956,244,-3956</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<connection>
<GID>187</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>189</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>192</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>194</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>197</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>199</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>201</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>203</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-460,231.5,-460</points>
<connection>
<GID>4647</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4643</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4639</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4635</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4631</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4627</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4623</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4619</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4615</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-4025,62.5,-3860</points>
<connection>
<GID>231</GID>
<name>N_in1</name></connection>
<connection>
<GID>204</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 12</intersection>
<intersection>-3981 11</intersection>
<intersection>-3962 10</intersection>
<intersection>-3943.5 9</intersection>
<intersection>-3921.5 8</intersection>
<intersection>-3903 7</intersection>
<intersection>-3884 6</intersection>
<intersection>-3865.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-3865.5,68,-3865.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>62.5,-3884,68,-3884</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>62.5,-3903,68,-3903</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>62.5,-3921.5,68,-3921.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>62.5,-3943.5,68,-3943.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>62.5,-3962,68,-3962</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>62.5,-3981,68,-3981</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>62.5,-3999.5,68,-3999.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-444.5,68.5,-444.5</points>
<connection>
<GID>4655</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-444.5,62.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-429,62.5,-429</points>
<connection>
<GID>4653</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-4024.5,85.5,-3859.5</points>
<connection>
<GID>235</GID>
<name>N_in1</name></connection>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<intersection>-4008 4</intersection>
<intersection>-3989.5 5</intersection>
<intersection>-3970.5 6</intersection>
<intersection>-3952 7</intersection>
<intersection>-3930 8</intersection>
<intersection>-3911.5 9</intersection>
<intersection>-3892.5 10</intersection>
<intersection>-3874 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>81,-4008,85.5,-4008</points>
<intersection>81 12</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>81,-3989.5,85.5,-3989.5</points>
<intersection>81 14</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>81,-3970.5,85.5,-3970.5</points>
<intersection>81 13</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>81,-3952,85.5,-3952</points>
<intersection>81 15</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>81,-3930,85.5,-3930</points>
<intersection>81 18</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>81,-3911.5,85.5,-3911.5</points>
<intersection>81 19</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>81,-3892.5,85.5,-3892.5</points>
<intersection>81 20</intersection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>81,-3874,85.5,-3874</points>
<intersection>81 21</intersection>
<intersection>85.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>81,-4009.5,81,-4008</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-4008 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>81,-3972,81,-3970.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>81,-3991,81,-3989.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>81,-3953.5,81,-3952</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>-3952 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>81,-3931.5,81,-3930</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>-3930 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>81,-3913,81,-3911.5</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>81,-3894,81,-3892.5</points>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>81,-3875.5,81,-3874</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-3874 11</intersection></vsegment></shape></wire>
<wire>
<ID>3267</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-444.5,91.5,-444.5</points>
<connection>
<GID>4659</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-444.5,85.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-429,85.5,-429</points>
<connection>
<GID>4657</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-4024.5,88.5,-3860</points>
<connection>
<GID>237</GID>
<name>N_in1</name></connection>
<connection>
<GID>206</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 10</intersection>
<intersection>-3981 9</intersection>
<intersection>-3962 8</intersection>
<intersection>-3943.5 7</intersection>
<intersection>-3921.5 6</intersection>
<intersection>-3903 5</intersection>
<intersection>-3884 4</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-3865.5,91,-3865.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>88.5,-3884,91,-3884</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>88.5,-3903,91,-3903</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>88.5,-3921.5,91,-3921.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>88.5,-3943.5,91,-3943.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>88.5,-3962,91,-3962</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>88.5,-3981,91,-3981</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>88.5,-3999.5,91,-3999.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-444.5,116.5,-444.5</points>
<connection>
<GID>4663</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-444.5,110.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-429,110.5,-429</points>
<connection>
<GID>4661</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-4024.5,108,-3859.5</points>
<connection>
<GID>239</GID>
<name>N_in1</name></connection>
<connection>
<GID>207</GID>
<name>N_in0</name></connection>
<intersection>-4008 6</intersection>
<intersection>-3989.5 7</intersection>
<intersection>-3970.5 8</intersection>
<intersection>-3952 9</intersection>
<intersection>-3930 10</intersection>
<intersection>-3911.5 11</intersection>
<intersection>-3892.5 12</intersection>
<intersection>-3874 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>104,-4008,108,-4008</points>
<intersection>104 14</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>104,-3989.5,108,-3989.5</points>
<intersection>104 16</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>104,-3970.5,108,-3970.5</points>
<intersection>104 15</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>104,-3952,108,-3952</points>
<intersection>104 17</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>104,-3930,108,-3930</points>
<intersection>104 20</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>104,-3911.5,108,-3911.5</points>
<intersection>104 21</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>104,-3892.5,108,-3892.5</points>
<intersection>104 22</intersection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>104,-3874,108,-3874</points>
<intersection>104 23</intersection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>104,-4009.5,104,-4008</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-4008 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>104,-3972,104,-3970.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>104,-3991,104,-3989.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>104,-3953.5,104,-3952</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>-3952 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>104,-3931.5,104,-3930</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-3930 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>104,-3913,104,-3911.5</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>104,-3894,104,-3892.5</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>104,-3875.5,104,-3874</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-3874 13</intersection></vsegment></shape></wire>
<wire>
<ID>3269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-444.5,139.5,-444.5</points>
<connection>
<GID>4304</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-444.5,133.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-429,133.5,-429</points>
<connection>
<GID>4302</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-4024.5,111.5,-3859.5</points>
<connection>
<GID>241</GID>
<name>N_in1</name></connection>
<connection>
<GID>208</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 13</intersection>
<intersection>-3981 12</intersection>
<intersection>-3962 11</intersection>
<intersection>-3943.5 10</intersection>
<intersection>-3921.5 9</intersection>
<intersection>-3903 8</intersection>
<intersection>-3884 7</intersection>
<intersection>-3865.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>111.5,-3865.5,116,-3865.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111.5,-3884,116,-3884</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111.5,-3903,116,-3903</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111.5,-3921.5,116,-3921.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111.5,-3943.5,116,-3943.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>111.5,-3962,116,-3962</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>111.5,-3981,116,-3981</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111.5,-3999.5,116,-3999.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-444.5,162.5,-444.5</points>
<connection>
<GID>4308</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-444.5,156.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-429,156.5,-429</points>
<connection>
<GID>4306</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-4024.5,132.5,-3860</points>
<connection>
<GID>243</GID>
<name>N_in1</name></connection>
<connection>
<GID>209</GID>
<name>N_in0</name></connection>
<intersection>-4008 6</intersection>
<intersection>-3989.5 7</intersection>
<intersection>-3970.5 8</intersection>
<intersection>-3952 9</intersection>
<intersection>-3930 10</intersection>
<intersection>-3911.5 11</intersection>
<intersection>-3892.5 12</intersection>
<intersection>-3874 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>129,-4008,132.5,-4008</points>
<intersection>129 14</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>129,-3989.5,132.5,-3989.5</points>
<intersection>129 16</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>129,-3970.5,132.5,-3970.5</points>
<intersection>129 15</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>129,-3952,132.5,-3952</points>
<intersection>129 17</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>129,-3930,132.5,-3930</points>
<intersection>129 20</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>129,-3911.5,132.5,-3911.5</points>
<intersection>129 21</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>129,-3892.5,132.5,-3892.5</points>
<intersection>129 22</intersection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>129,-3874,132.5,-3874</points>
<intersection>129 23</intersection>
<intersection>132.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>129,-4009.5,129,-4008</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-4008 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>129,-3972,129,-3970.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>129,-3991,129,-3989.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>129,-3953.5,129,-3952</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-3952 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>129,-3931.5,129,-3930</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>-3930 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>129,-3913,129,-3911.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>129,-3894,129,-3892.5</points>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>129,-3875.5,129,-3874</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-3874 13</intersection></vsegment></shape></wire>
<wire>
<ID>3271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-444.5,185.5,-444.5</points>
<connection>
<GID>4312</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-444.5,179.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-429,179.5,-429</points>
<connection>
<GID>4310</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-4024.5,136.5,-3859.5</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<connection>
<GID>210</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 13</intersection>
<intersection>-3981 12</intersection>
<intersection>-3962 11</intersection>
<intersection>-3943.5 10</intersection>
<intersection>-3921.5 9</intersection>
<intersection>-3903 8</intersection>
<intersection>-3884 7</intersection>
<intersection>-3865.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>136.5,-3865.5,139,-3865.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>136.5,-3884,139,-3884</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>136.5,-3903,139,-3903</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>136.5,-3921.5,139,-3921.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>136.5,-3943.5,139,-3943.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>136.5,-3962,139,-3962</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>136.5,-3981,139,-3981</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>136.5,-3999.5,139,-3999.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3272</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-444.5,210.5,-444.5</points>
<connection>
<GID>4316</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-444.5,204.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-429,204.5,-429</points>
<connection>
<GID>4314</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-4024.5,155,-3859.5</points>
<connection>
<GID>249</GID>
<name>N_in1</name></connection>
<connection>
<GID>211</GID>
<name>N_in0</name></connection>
<intersection>-4008 6</intersection>
<intersection>-3989.5 7</intersection>
<intersection>-3970.5 8</intersection>
<intersection>-3952 9</intersection>
<intersection>-3930 10</intersection>
<intersection>-3911.5 11</intersection>
<intersection>-3892.5 12</intersection>
<intersection>-3874 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>152,-4008,155,-4008</points>
<intersection>152 14</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>152,-3989.5,155,-3989.5</points>
<intersection>152 15</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>152,-3970.5,155,-3970.5</points>
<intersection>152 16</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-3952,155,-3952</points>
<intersection>152 17</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>152,-3930,155,-3930</points>
<intersection>152 20</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>152,-3911.5,155,-3911.5</points>
<intersection>152 21</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>152,-3892.5,155,-3892.5</points>
<intersection>152 22</intersection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>152,-3874,155,-3874</points>
<intersection>152 23</intersection>
<intersection>155 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>152,-4009.5,152,-4008</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>-4008 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>152,-3991,152,-3989.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>152,-3972,152,-3970.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>152,-3953.5,152,-3952</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>-3952 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>152,-3931.5,152,-3930</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>-3930 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>152,-3913,152,-3911.5</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>152,-3894,152,-3892.5</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>152,-3875.5,152,-3874</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-3874 13</intersection></vsegment></shape></wire>
<wire>
<ID>3273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-444.5,233.5,-444.5</points>
<connection>
<GID>4320</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-444.5,227.5,-429</points>
<intersection>-444.5 1</intersection>
<intersection>-429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-429,227.5,-429</points>
<connection>
<GID>4318</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-4024.5,159,-3859.5</points>
<connection>
<GID>251</GID>
<name>N_in1</name></connection>
<connection>
<GID>213</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 13</intersection>
<intersection>-3981 12</intersection>
<intersection>-3962 11</intersection>
<intersection>-3943.5 10</intersection>
<intersection>-3921.5 9</intersection>
<intersection>-3903 8</intersection>
<intersection>-3884 7</intersection>
<intersection>-3865.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>159,-3865.5,162,-3865.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>159,-3884,162,-3884</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>159,-3903,162,-3903</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>159,-3921.5,162,-3921.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>159,-3943.5,162,-3943.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>159,-3962,162,-3962</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>159,-3981,162,-3981</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>159,-3999.5,162,-3999.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>3274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-432,220.5,-432</points>
<connection>
<GID>4318</GID>
<name>clock</name></connection>
<connection>
<GID>4314</GID>
<name>clock</name></connection>
<connection>
<GID>4310</GID>
<name>clock</name></connection>
<connection>
<GID>4306</GID>
<name>clock</name></connection>
<connection>
<GID>4302</GID>
<name>clock</name></connection>
<connection>
<GID>4661</GID>
<name>clock</name></connection>
<connection>
<GID>4657</GID>
<name>clock</name></connection>
<connection>
<GID>4653</GID>
<name>clock</name></connection>
<connection>
<GID>4649</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-4024,178,-3859.5</points>
<connection>
<GID>253</GID>
<name>N_in1</name></connection>
<connection>
<GID>215</GID>
<name>N_in0</name></connection>
<intersection>-4008 6</intersection>
<intersection>-3989.5 7</intersection>
<intersection>-3970.5 8</intersection>
<intersection>-3952 9</intersection>
<intersection>-3930 10</intersection>
<intersection>-3911.5 11</intersection>
<intersection>-3892.5 12</intersection>
<intersection>-3874 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>175,-4008,178,-4008</points>
<intersection>175 15</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>175,-3989.5,178,-3989.5</points>
<intersection>175 16</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>175,-3970.5,178,-3970.5</points>
<intersection>175 17</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>175,-3952,178,-3952</points>
<intersection>175 18</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>175,-3930,178,-3930</points>
<intersection>175 21</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>175,-3911.5,178,-3911.5</points>
<intersection>175 22</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>175,-3892.5,178,-3892.5</points>
<intersection>175 23</intersection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>175,-3874,178,-3874</points>
<intersection>175 14</intersection>
<intersection>178 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>175,-3875.5,175,-3874</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-3874 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>175,-4009.5,175,-4008</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>-4008 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>175,-3991,175,-3989.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>175,-3972,175,-3970.5</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>175,-3953.5,175,-3952</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>-3952 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>175,-3931.5,175,-3930</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>-3930 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>175,-3913,175,-3911.5</points>
<connection>
<GID>329</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>175,-3894,175,-3892.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 12</intersection></vsegment></shape></wire>
<wire>
<ID>3275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-441.5,231.5,-441.5</points>
<connection>
<GID>4320</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4316</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4312</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4308</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4304</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4663</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4659</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4655</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4651</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-4024,183,-3859.5</points>
<connection>
<GID>255</GID>
<name>N_in1</name></connection>
<connection>
<GID>217</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 13</intersection>
<intersection>-3981 12</intersection>
<intersection>-3962 11</intersection>
<intersection>-3943.5 10</intersection>
<intersection>-3921.5 9</intersection>
<intersection>-3903 8</intersection>
<intersection>-3884 7</intersection>
<intersection>-3865.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>183,-3865.5,185,-3865.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>183,-3884,185,-3884</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>183,-3903,185,-3903</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>183,-3921.5,185,-3921.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183,-3943.5,185,-3943.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183,-3962,185,-3962</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183,-3981,185,-3981</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183,-3999.5,185,-3999.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>3276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-425.5,68.5,-425.5</points>
<connection>
<GID>4330</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-425.5,62.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-410,62.5,-410</points>
<connection>
<GID>4328</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-4023.5,201,-3859.5</points>
<connection>
<GID>257</GID>
<name>N_in1</name></connection>
<connection>
<GID>221</GID>
<name>N_in0</name></connection>
<intersection>-4008 16</intersection>
<intersection>-3989.5 15</intersection>
<intersection>-3970.5 14</intersection>
<intersection>-3952 13</intersection>
<intersection>-3930 12</intersection>
<intersection>-3911.5 11</intersection>
<intersection>-3892.5 10</intersection>
<intersection>-3874 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>198,-3874,201,-3874</points>
<intersection>198 17</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>198,-3892.5,201,-3892.5</points>
<intersection>198 26</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>198,-3911.5,201,-3911.5</points>
<intersection>198 25</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>198,-3930,201,-3930</points>
<intersection>198 24</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>198,-3952,201,-3952</points>
<intersection>198 21</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>198,-3970.5,201,-3970.5</points>
<intersection>198 20</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>198,-3989.5,201,-3989.5</points>
<intersection>198 19</intersection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>198,-4008,201,-4008</points>
<intersection>198 18</intersection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>198,-3875.5,198,-3874</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-3874 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>198,-4009.5,198,-4008</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-4008 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>198,-3991,198,-3989.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>198,-3972,198,-3970.5</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>198,-3953.5,198,-3952</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>-3952 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>198,-3931.5,198,-3930</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>-3930 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>198,-3913,198,-3911.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>198,-3894,198,-3892.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>3277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-425.5,91.5,-425.5</points>
<connection>
<GID>4335</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-425.5,85.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-410,85.5,-410</points>
<connection>
<GID>4333</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-4023.5,205.5,-3859.5</points>
<connection>
<GID>259</GID>
<name>N_in1</name></connection>
<connection>
<GID>219</GID>
<name>N_in0</name></connection>
<intersection>-3999.5 13</intersection>
<intersection>-3981 12</intersection>
<intersection>-3962 11</intersection>
<intersection>-3943.5 10</intersection>
<intersection>-3921.5 9</intersection>
<intersection>-3903 8</intersection>
<intersection>-3884 7</intersection>
<intersection>-3865.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>205.5,-3865.5,210,-3865.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205.5,-3884,210,-3884</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>205.5,-3903,210,-3903</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>205.5,-3921.5,210,-3921.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>205.5,-3943.5,210,-3943.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205.5,-3962,210,-3962</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>205.5,-3981,210,-3981</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>205.5,-3999.5,210,-3999.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-425.5,116.5,-425.5</points>
<connection>
<GID>4340</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-425.5,110.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-410,110.5,-410</points>
<connection>
<GID>4338</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-4023,226.5,-3860</points>
<connection>
<GID>261</GID>
<name>N_in1</name></connection>
<connection>
<GID>223</GID>
<name>N_in0</name></connection>
<intersection>-4008 6</intersection>
<intersection>-3989.5 7</intersection>
<intersection>-3970.5 8</intersection>
<intersection>-3952 9</intersection>
<intersection>-3930 10</intersection>
<intersection>-3911.5 11</intersection>
<intersection>-3892.5 12</intersection>
<intersection>-3874 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>223,-4008,226.5,-4008</points>
<intersection>223 15</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>223,-3989.5,226.5,-3989.5</points>
<intersection>223 16</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>223,-3970.5,226.5,-3970.5</points>
<intersection>223 17</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>223,-3952,226.5,-3952</points>
<intersection>223 18</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>223,-3930,226.5,-3930</points>
<intersection>223 21</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>223,-3911.5,226.5,-3911.5</points>
<intersection>223 22</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>223,-3892.5,226.5,-3892.5</points>
<intersection>223 23</intersection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>223,-3874,226.5,-3874</points>
<intersection>223 14</intersection>
<intersection>226.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>223,-3875.5,223,-3874</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-3874 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>223,-4009.5,223,-4008</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>-4008 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>223,-3991,223,-3989.5</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>223,-3972,223,-3970.5</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>223,-3953.5,223,-3952</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>-3952 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>223,-3931.5,223,-3930</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>-3930 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>223,-3913,223,-3911.5</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>223,-3894,223,-3892.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 12</intersection></vsegment></shape></wire>
<wire>
<ID>3279</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-425.5,139.5,-425.5</points>
<connection>
<GID>4345</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-425.5,133.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-410,133.5,-410</points>
<connection>
<GID>4343</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-4023,230,-3860</points>
<connection>
<GID>265</GID>
<name>N_in0</name></connection>
<connection>
<GID>263</GID>
<name>N_in1</name></connection>
<intersection>-3999.5 11</intersection>
<intersection>-3981 10</intersection>
<intersection>-3962 9</intersection>
<intersection>-3943.5 7</intersection>
<intersection>-3921.5 6</intersection>
<intersection>-3903 5</intersection>
<intersection>-3884 4</intersection>
<intersection>-3865.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>230,-3865.5,233,-3865.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>230,-3884,233,-3884</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>230,-3903,233,-3903</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>230,-3921.5,233,-3921.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>230,-3943.5,233,-3943.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>230,-3962,233,-3962</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>230,-3981,233,-3981</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>230,-3999.5,233,-3999.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>3280</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-425.5,162.5,-425.5</points>
<connection>
<GID>4350</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-425.5,156.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-410,156.5,-410</points>
<connection>
<GID>4348</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-4023,251,-3861</points>
<connection>
<GID>267</GID>
<name>N_in1</name></connection>
<connection>
<GID>225</GID>
<name>N_in0</name></connection>
<intersection>-4008 11</intersection>
<intersection>-3989.5 10</intersection>
<intersection>-3970.5 9</intersection>
<intersection>-3952 8</intersection>
<intersection>-3930 7</intersection>
<intersection>-3911.5 6</intersection>
<intersection>-3892.5 5</intersection>
<intersection>-3874 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>246,-3874,251,-3874</points>
<intersection>246 12</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>246,-3892.5,251,-3892.5</points>
<intersection>246 21</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>246,-3911.5,251,-3911.5</points>
<intersection>246 20</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>246,-3930,251,-3930</points>
<intersection>246 19</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>246,-3952,251,-3952</points>
<intersection>246 16</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>246,-3970.5,251,-3970.5</points>
<intersection>246 15</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>246,-3989.5,251,-3989.5</points>
<intersection>246 14</intersection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>246,-4008,251,-4008</points>
<intersection>246 13</intersection>
<intersection>251 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>246,-3875.5,246,-3874</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-3874 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>246,-4009.5,246,-4008</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-4008 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>246,-3991,246,-3989.5</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>-3989.5 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>246,-3972,246,-3970.5</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>-3970.5 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>246,-3953.5,246,-3952</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-3952 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>246,-3931.5,246,-3930</points>
<connection>
<GID>305</GID>
<name>OUT_0</name></connection>
<intersection>-3930 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>246,-3913,246,-3911.5</points>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection>
<intersection>-3911.5 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>246,-3894,246,-3892.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-3892.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>3281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-425.5,185.5,-425.5</points>
<connection>
<GID>4353</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-425.5,179.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-410,179.5,-410</points>
<connection>
<GID>4352</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-99,-3867.5,40.5,-3867.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-99 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-99,-3877,-99,-3851.5</points>
<intersection>-3877 4</intersection>
<intersection>-3867.5 2</intersection>
<intersection>-3851.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-99,-3877,52,-3877</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-99 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-106,-3851.5,-99,-3851.5</points>
<connection>
<GID>149</GID>
<name>OUT_7</name></connection>
<intersection>-99 3</intersection></hsegment></shape></wire>
<wire>
<ID>3282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-425.5,210.5,-425.5</points>
<connection>
<GID>4356</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-425.5,204.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-410,204.5,-410</points>
<connection>
<GID>4355</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-100,-3886,40.5,-3886</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-100 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-100,-3895.5,-100,-3852.5</points>
<intersection>-3895.5 5</intersection>
<intersection>-3886 2</intersection>
<intersection>-3852.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-100,-3895.5,52,-3895.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>-100 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-106,-3852.5,-100,-3852.5</points>
<connection>
<GID>149</GID>
<name>OUT_6</name></connection>
<intersection>-100 4</intersection></hsegment></shape></wire>
<wire>
<ID>3283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-425.5,233.5,-425.5</points>
<connection>
<GID>4358</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-425.5,227.5,-410</points>
<intersection>-425.5 1</intersection>
<intersection>-410 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-410,227.5,-410</points>
<connection>
<GID>4357</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-101,-3905,40.5,-3905</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>-101 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-101,-3914.5,-101,-3853.5</points>
<intersection>-3914.5 4</intersection>
<intersection>-3905 2</intersection>
<intersection>-3853.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-101,-3914.5,52,-3914.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-101 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-106,-3853.5,-101,-3853.5</points>
<connection>
<GID>149</GID>
<name>OUT_5</name></connection>
<intersection>-101 3</intersection></hsegment></shape></wire>
<wire>
<ID>3284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-413,220.5,-413</points>
<connection>
<GID>4357</GID>
<name>clock</name></connection>
<connection>
<GID>4355</GID>
<name>clock</name></connection>
<connection>
<GID>4352</GID>
<name>clock</name></connection>
<connection>
<GID>4348</GID>
<name>clock</name></connection>
<connection>
<GID>4343</GID>
<name>clock</name></connection>
<connection>
<GID>4338</GID>
<name>clock</name></connection>
<connection>
<GID>4333</GID>
<name>clock</name></connection>
<connection>
<GID>4328</GID>
<name>clock</name></connection>
<connection>
<GID>4323</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-102,-3923.5,40.5,-3923.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-102 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-102,-3933,-102,-3854.5</points>
<intersection>-3933 4</intersection>
<intersection>-3923.5 2</intersection>
<intersection>-3854.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-102,-3933,52,-3933</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>-102 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3854.5,-102,-3854.5</points>
<connection>
<GID>149</GID>
<name>OUT_4</name></connection>
<intersection>-102 3</intersection></hsegment></shape></wire>
<wire>
<ID>3285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-422.5,231.5,-422.5</points>
<connection>
<GID>4358</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4356</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4353</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4350</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4345</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4340</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4335</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4330</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4325</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-103,-3945.5,40.5,-3945.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-103 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-103,-3955,-103,-3855.5</points>
<intersection>-3955 4</intersection>
<intersection>-3945.5 1</intersection>
<intersection>-3855.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-103,-3955,51.5,-3955</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-103 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3855.5,-103,-3855.5</points>
<connection>
<GID>149</GID>
<name>OUT_3</name></connection>
<intersection>-103 3</intersection></hsegment></shape></wire>
<wire>
<ID>3286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-407,68.5,-407</points>
<connection>
<GID>4362</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-407,62.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-391.5,62.5,-391.5</points>
<connection>
<GID>4361</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104,-3964,40.5,-3964</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-104 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-104,-3973.5,-104,-3856.5</points>
<intersection>-3973.5 4</intersection>
<intersection>-3964 1</intersection>
<intersection>-3856.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-104,-3973.5,51.5,-3973.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-104 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3856.5,-104,-3856.5</points>
<connection>
<GID>149</GID>
<name>OUT_2</name></connection>
<intersection>-104 3</intersection></hsegment></shape></wire>
<wire>
<ID>3287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-407,91.5,-407</points>
<connection>
<GID>4364</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-407,85.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-391.5,85.5,-391.5</points>
<connection>
<GID>4363</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105,-3983,40.5,-3983</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-105 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-105,-3992.5,-105,-3857.5</points>
<intersection>-3992.5 4</intersection>
<intersection>-3983 1</intersection>
<intersection>-3857.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-105,-3992.5,51.5,-3992.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-105 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-106,-3857.5,-105,-3857.5</points>
<connection>
<GID>149</GID>
<name>OUT_1</name></connection>
<intersection>-105 3</intersection></hsegment></shape></wire>
<wire>
<ID>3288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-407,116.5,-407</points>
<connection>
<GID>4366</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-407,110.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-391.5,110.5,-391.5</points>
<connection>
<GID>4365</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-4001.5,40.5,-4001.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-106 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-106,-4011,-106,-3858.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>-4011 4</intersection>
<intersection>-4001.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-106,-4011,51.5,-4011</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-106 3</intersection></hsegment></shape></wire>
<wire>
<ID>3289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-407,139.5,-407</points>
<connection>
<GID>4368</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-407,133.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-391.5,133.5,-391.5</points>
<connection>
<GID>4367</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-4025,39.5,-3860</points>
<connection>
<GID>285</GID>
<name>N_in1</name></connection>
<connection>
<GID>277</GID>
<name>N_in0</name></connection>
<intersection>-4003.5 10</intersection>
<intersection>-3985 9</intersection>
<intersection>-3966 8</intersection>
<intersection>-3947.5 7</intersection>
<intersection>-3925.5 6</intersection>
<intersection>-3907 5</intersection>
<intersection>-3888 4</intersection>
<intersection>-3869.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>39.5,-3869.5,40.5,-3869.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39.5,-3888,40.5,-3888</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>39.5,-3907,40.5,-3907</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>39.5,-3925.5,40.5,-3925.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>39.5,-3947.5,40.5,-3947.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>39.5,-3966,40.5,-3966</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>39.5,-3985,40.5,-3985</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>39.5,-4003.5,40.5,-4003.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-407,162.5,-407</points>
<connection>
<GID>4370</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-407,156.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-391.5,156.5,-391.5</points>
<connection>
<GID>4369</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-4025,49.5,-3860</points>
<connection>
<GID>281</GID>
<name>N_in1</name></connection>
<connection>
<GID>273</GID>
<name>N_in0</name></connection>
<intersection>-4013 3</intersection>
<intersection>-3994.5 5</intersection>
<intersection>-3975.5 7</intersection>
<intersection>-3957 9</intersection>
<intersection>-3935 11</intersection>
<intersection>-3916.5 13</intersection>
<intersection>-3897.5 15</intersection>
<intersection>-3879 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49.5,-4013,51.5,-4013</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>49.5,-3994.5,51.5,-3994.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>49.5,-3975.5,51.5,-3975.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>49.5,-3957,51.5,-3957</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>49.5,-3935,52,-3935</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>49.5,-3916.5,52,-3916.5</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>49.5,-3897.5,52,-3897.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>49.5,-3879,52,-3879</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-407,185.5,-407</points>
<connection>
<GID>4372</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-407,179.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-391.5,179.5,-391.5</points>
<connection>
<GID>4371</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-3858,39.5,-3851.5</points>
<connection>
<GID>277</GID>
<name>N_in1</name></connection>
<connection>
<GID>147</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-407,210.5,-407</points>
<connection>
<GID>4374</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-407,204.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-391.5,204.5,-391.5</points>
<connection>
<GID>4373</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-3858,49.5,-3851.5</points>
<connection>
<GID>273</GID>
<name>N_in1</name></connection>
<connection>
<GID>146</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-407,233.5,-407</points>
<connection>
<GID>4376</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-407,227.5,-391.5</points>
<intersection>-407 1</intersection>
<intersection>-391.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-391.5,227.5,-391.5</points>
<connection>
<GID>4375</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-3858,62.5,-3851.5</points>
<connection>
<GID>204</GID>
<name>N_in1</name></connection>
<connection>
<GID>127</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-394.5,220.5,-394.5</points>
<connection>
<GID>4375</GID>
<name>clock</name></connection>
<connection>
<GID>4373</GID>
<name>clock</name></connection>
<connection>
<GID>4371</GID>
<name>clock</name></connection>
<connection>
<GID>4369</GID>
<name>clock</name></connection>
<connection>
<GID>4367</GID>
<name>clock</name></connection>
<connection>
<GID>4365</GID>
<name>clock</name></connection>
<connection>
<GID>4363</GID>
<name>clock</name></connection>
<connection>
<GID>4361</GID>
<name>clock</name></connection>
<connection>
<GID>4359</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-3857.5,85.5,-3851</points>
<connection>
<GID>205</GID>
<name>N_in1</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-404,231.5,-404</points>
<connection>
<GID>4376</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4374</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4372</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4370</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4368</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4366</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4364</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4362</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4360</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-3858,88.5,-3851</points>
<connection>
<GID>206</GID>
<name>N_in1</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-473,50,-308</points>
<connection>
<GID>4392</GID>
<name>N_in1</name></connection>
<connection>
<GID>4377</GID>
<name>N_in0</name></connection>
<intersection>-447.5 12</intersection>
<intersection>-429 11</intersection>
<intersection>-410 10</intersection>
<intersection>-391.5 9</intersection>
<intersection>-369.5 8</intersection>
<intersection>-351 7</intersection>
<intersection>-332 6</intersection>
<intersection>-313.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-313.5,55.5,-313.5</points>
<connection>
<GID>4581</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>50,-332,55.5,-332</points>
<connection>
<GID>4545</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>50,-351,55.5,-351</points>
<connection>
<GID>4509</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>50,-369.5,55.5,-369.5</points>
<connection>
<GID>4455</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>50,-391.5,55.5,-391.5</points>
<connection>
<GID>4361</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>50,-410,55.5,-410</points>
<connection>
<GID>4328</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>50,-429,55.5,-429</points>
<connection>
<GID>4653</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>50,-447.5,55.5,-447.5</points>
<connection>
<GID>4617</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-3857.5,108,-3851</points>
<connection>
<GID>207</GID>
<name>N_in1</name></connection>
<connection>
<GID>130</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-472.5,73,-307.5</points>
<connection>
<GID>4393</GID>
<name>N_in1</name></connection>
<connection>
<GID>4378</GID>
<name>N_in0</name></connection>
<intersection>-456.5 4</intersection>
<intersection>-438 5</intersection>
<intersection>-419 6</intersection>
<intersection>-400.5 7</intersection>
<intersection>-378.5 8</intersection>
<intersection>-360 9</intersection>
<intersection>-341 10</intersection>
<intersection>-322.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-456.5,73,-456.5</points>
<intersection>68.5 12</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68.5,-438,73,-438</points>
<intersection>68.5 13</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68.5,-419,73,-419</points>
<intersection>68.5 14</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68.5,-400.5,73,-400.5</points>
<intersection>68.5 15</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-378.5,73,-378.5</points>
<intersection>68.5 18</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68.5,-360,73,-360</points>
<intersection>68.5 19</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68.5,-341,73,-341</points>
<intersection>68.5 20</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>68.5,-322.5,73,-322.5</points>
<intersection>68.5 21</intersection>
<intersection>73 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>68.5,-457.5,68.5,-456.5</points>
<connection>
<GID>4619</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>68.5,-439,68.5,-438</points>
<connection>
<GID>4655</GID>
<name>OUT_0</name></connection>
<intersection>-438 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>68.5,-420,68.5,-419</points>
<connection>
<GID>4330</GID>
<name>OUT_0</name></connection>
<intersection>-419 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>68.5,-401.5,68.5,-400.5</points>
<connection>
<GID>4362</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>68.5,-379.5,68.5,-378.5</points>
<connection>
<GID>4461</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>68.5,-361,68.5,-360</points>
<connection>
<GID>4511</GID>
<name>OUT_0</name></connection>
<intersection>-360 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>68.5,-342,68.5,-341</points>
<connection>
<GID>4547</GID>
<name>OUT_0</name></connection>
<intersection>-341 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>68.5,-323.5,68.5,-322.5</points>
<connection>
<GID>4583</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-3857.5,111.5,-3851</points>
<connection>
<GID>208</GID>
<name>N_in1</name></connection>
<connection>
<GID>131</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-472.5,76,-308</points>
<connection>
<GID>4394</GID>
<name>N_in1</name></connection>
<connection>
<GID>4379</GID>
<name>N_in0</name></connection>
<intersection>-447.5 10</intersection>
<intersection>-429 9</intersection>
<intersection>-410 8</intersection>
<intersection>-391.5 7</intersection>
<intersection>-369.5 6</intersection>
<intersection>-351 5</intersection>
<intersection>-332 4</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>76,-313.5,78.5,-313.5</points>
<connection>
<GID>4585</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>76,-332,78.5,-332</points>
<connection>
<GID>4549</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>76,-351,78.5,-351</points>
<connection>
<GID>4513</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>76,-369.5,78.5,-369.5</points>
<connection>
<GID>4477</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>76,-391.5,78.5,-391.5</points>
<connection>
<GID>4363</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>76,-410,78.5,-410</points>
<connection>
<GID>4333</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>76,-429,78.5,-429</points>
<connection>
<GID>4657</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>76,-447.5,78.5,-447.5</points>
<connection>
<GID>4621</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-3858,132.5,-3851</points>
<connection>
<GID>209</GID>
<name>N_in1</name></connection>
<connection>
<GID>132</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-472.5,95.5,-307.5</points>
<connection>
<GID>4395</GID>
<name>N_in1</name></connection>
<connection>
<GID>4380</GID>
<name>N_in0</name></connection>
<intersection>-456.5 6</intersection>
<intersection>-438 7</intersection>
<intersection>-419 8</intersection>
<intersection>-400.5 9</intersection>
<intersection>-378.5 10</intersection>
<intersection>-360 11</intersection>
<intersection>-341 12</intersection>
<intersection>-322.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91.5,-456.5,95.5,-456.5</points>
<intersection>91.5 14</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>91.5,-438,95.5,-438</points>
<intersection>91.5 15</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>91.5,-419,95.5,-419</points>
<intersection>91.5 16</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>91.5,-400.5,95.5,-400.5</points>
<intersection>91.5 17</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>91.5,-378.5,95.5,-378.5</points>
<intersection>91.5 20</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>91.5,-360,95.5,-360</points>
<intersection>91.5 21</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>91.5,-341,95.5,-341</points>
<intersection>91.5 22</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>91.5,-322.5,95.5,-322.5</points>
<intersection>91.5 23</intersection>
<intersection>95.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>91.5,-457.5,91.5,-456.5</points>
<connection>
<GID>4623</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>91.5,-439,91.5,-438</points>
<connection>
<GID>4659</GID>
<name>OUT_0</name></connection>
<intersection>-438 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>91.5,-420,91.5,-419</points>
<connection>
<GID>4335</GID>
<name>OUT_0</name></connection>
<intersection>-419 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>91.5,-401.5,91.5,-400.5</points>
<connection>
<GID>4364</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>91.5,-379.5,91.5,-378.5</points>
<connection>
<GID>4479</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>91.5,-361,91.5,-360</points>
<connection>
<GID>4515</GID>
<name>OUT_0</name></connection>
<intersection>-360 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>91.5,-342,91.5,-341</points>
<connection>
<GID>4551</GID>
<name>OUT_0</name></connection>
<intersection>-341 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>91.5,-323.5,91.5,-322.5</points>
<connection>
<GID>4587</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-3857.5,136.5,-3851</points>
<connection>
<GID>210</GID>
<name>N_in1</name></connection>
<connection>
<GID>133</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-472.5,99,-307.5</points>
<connection>
<GID>4396</GID>
<name>N_in1</name></connection>
<connection>
<GID>4381</GID>
<name>N_in0</name></connection>
<intersection>-447.5 13</intersection>
<intersection>-429 12</intersection>
<intersection>-410 11</intersection>
<intersection>-391.5 10</intersection>
<intersection>-369.5 9</intersection>
<intersection>-351 8</intersection>
<intersection>-332 7</intersection>
<intersection>-313.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>99,-313.5,103.5,-313.5</points>
<connection>
<GID>4589</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>99,-332,103.5,-332</points>
<connection>
<GID>4553</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>99,-351,103.5,-351</points>
<connection>
<GID>4517</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>99,-369.5,103.5,-369.5</points>
<connection>
<GID>4481</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>99,-391.5,103.5,-391.5</points>
<connection>
<GID>4365</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>99,-410,103.5,-410</points>
<connection>
<GID>4338</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>99,-429,103.5,-429</points>
<connection>
<GID>4661</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>99,-447.5,103.5,-447.5</points>
<connection>
<GID>4625</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-3857.5,155,-3851</points>
<connection>
<GID>211</GID>
<name>N_in1</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-472.5,120,-308</points>
<connection>
<GID>4397</GID>
<name>N_in1</name></connection>
<connection>
<GID>4382</GID>
<name>N_in0</name></connection>
<intersection>-456.5 6</intersection>
<intersection>-438 7</intersection>
<intersection>-419 8</intersection>
<intersection>-400.5 9</intersection>
<intersection>-378.5 10</intersection>
<intersection>-360 11</intersection>
<intersection>-341 12</intersection>
<intersection>-322.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116.5,-456.5,120,-456.5</points>
<intersection>116.5 14</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116.5,-438,120,-438</points>
<intersection>116.5 15</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>116.5,-419,120,-419</points>
<intersection>116.5 16</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116.5,-400.5,120,-400.5</points>
<intersection>116.5 17</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116.5,-378.5,120,-378.5</points>
<intersection>116.5 20</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>116.5,-360,120,-360</points>
<intersection>116.5 21</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>116.5,-341,120,-341</points>
<intersection>116.5 22</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>116.5,-322.5,120,-322.5</points>
<intersection>116.5 23</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>116.5,-457.5,116.5,-456.5</points>
<connection>
<GID>4627</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>116.5,-439,116.5,-438</points>
<connection>
<GID>4663</GID>
<name>OUT_0</name></connection>
<intersection>-438 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>116.5,-420,116.5,-419</points>
<connection>
<GID>4340</GID>
<name>OUT_0</name></connection>
<intersection>-419 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>116.5,-401.5,116.5,-400.5</points>
<connection>
<GID>4366</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>116.5,-379.5,116.5,-378.5</points>
<connection>
<GID>4483</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>116.5,-361,116.5,-360</points>
<connection>
<GID>4519</GID>
<name>OUT_0</name></connection>
<intersection>-360 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>116.5,-342,116.5,-341</points>
<connection>
<GID>4555</GID>
<name>OUT_0</name></connection>
<intersection>-341 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>116.5,-323.5,116.5,-322.5</points>
<connection>
<GID>4591</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-3857.5,159,-3851</points>
<connection>
<GID>213</GID>
<name>N_in1</name></connection>
<connection>
<GID>135</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-472.5,124,-307.5</points>
<connection>
<GID>4398</GID>
<name>N_in1</name></connection>
<connection>
<GID>4383</GID>
<name>N_in0</name></connection>
<intersection>-447.5 13</intersection>
<intersection>-429 12</intersection>
<intersection>-410 11</intersection>
<intersection>-391.5 10</intersection>
<intersection>-369.5 9</intersection>
<intersection>-351 8</intersection>
<intersection>-332 7</intersection>
<intersection>-313.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>124,-313.5,126.5,-313.5</points>
<connection>
<GID>4593</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>124,-332,126.5,-332</points>
<connection>
<GID>4557</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>124,-351,126.5,-351</points>
<connection>
<GID>4521</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>124,-369.5,126.5,-369.5</points>
<connection>
<GID>4485</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>124,-391.5,126.5,-391.5</points>
<connection>
<GID>4367</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>124,-410,126.5,-410</points>
<connection>
<GID>4343</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>124,-429,126.5,-429</points>
<connection>
<GID>4302</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>124,-447.5,126.5,-447.5</points>
<connection>
<GID>4629</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-3857.5,178,-3850.5</points>
<connection>
<GID>215</GID>
<name>N_in1</name></connection>
<connection>
<GID>136</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-472.5,142.5,-307.5</points>
<connection>
<GID>4399</GID>
<name>N_in1</name></connection>
<connection>
<GID>4384</GID>
<name>N_in0</name></connection>
<intersection>-456.5 6</intersection>
<intersection>-438 7</intersection>
<intersection>-419 8</intersection>
<intersection>-400.5 9</intersection>
<intersection>-378.5 10</intersection>
<intersection>-360 11</intersection>
<intersection>-341 12</intersection>
<intersection>-322.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139.5,-456.5,142.5,-456.5</points>
<intersection>139.5 14</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139.5,-438,142.5,-438</points>
<intersection>139.5 15</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>139.5,-419,142.5,-419</points>
<intersection>139.5 16</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>139.5,-400.5,142.5,-400.5</points>
<intersection>139.5 17</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>139.5,-378.5,142.5,-378.5</points>
<intersection>139.5 20</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139.5,-360,142.5,-360</points>
<intersection>139.5 21</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>139.5,-341,142.5,-341</points>
<intersection>139.5 22</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>139.5,-322.5,142.5,-322.5</points>
<intersection>139.5 23</intersection>
<intersection>142.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>139.5,-457.5,139.5,-456.5</points>
<connection>
<GID>4631</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>139.5,-439,139.5,-438</points>
<connection>
<GID>4304</GID>
<name>OUT_0</name></connection>
<intersection>-438 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>139.5,-420,139.5,-419</points>
<connection>
<GID>4345</GID>
<name>OUT_0</name></connection>
<intersection>-419 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>139.5,-401.5,139.5,-400.5</points>
<connection>
<GID>4368</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>139.5,-379.5,139.5,-378.5</points>
<connection>
<GID>4487</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>139.5,-361,139.5,-360</points>
<connection>
<GID>4523</GID>
<name>OUT_0</name></connection>
<intersection>-360 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>139.5,-342,139.5,-341</points>
<connection>
<GID>4559</GID>
<name>OUT_0</name></connection>
<intersection>-341 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>139.5,-323.5,139.5,-322.5</points>
<connection>
<GID>4595</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-3857.5,183,-3850.5</points>
<connection>
<GID>217</GID>
<name>N_in1</name></connection>
<connection>
<GID>137</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-472.5,146.5,-307.5</points>
<connection>
<GID>4400</GID>
<name>N_in1</name></connection>
<connection>
<GID>4385</GID>
<name>N_in0</name></connection>
<intersection>-447.5 13</intersection>
<intersection>-429 12</intersection>
<intersection>-410 11</intersection>
<intersection>-391.5 10</intersection>
<intersection>-369.5 9</intersection>
<intersection>-351 8</intersection>
<intersection>-332 7</intersection>
<intersection>-313.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>146.5,-313.5,149.5,-313.5</points>
<connection>
<GID>4597</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>146.5,-332,149.5,-332</points>
<connection>
<GID>4561</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>146.5,-351,149.5,-351</points>
<connection>
<GID>4525</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>146.5,-369.5,149.5,-369.5</points>
<connection>
<GID>4489</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>146.5,-391.5,149.5,-391.5</points>
<connection>
<GID>4369</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>146.5,-410,149.5,-410</points>
<connection>
<GID>4348</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>146.5,-429,149.5,-429</points>
<connection>
<GID>4306</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>146.5,-447.5,149.5,-447.5</points>
<connection>
<GID>4633</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-3857.5,201,-3850</points>
<connection>
<GID>221</GID>
<name>N_in1</name></connection>
<connection>
<GID>138</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-472,165.5,-307.5</points>
<connection>
<GID>4401</GID>
<name>N_in1</name></connection>
<connection>
<GID>4386</GID>
<name>N_in0</name></connection>
<intersection>-456.5 6</intersection>
<intersection>-438 7</intersection>
<intersection>-419 8</intersection>
<intersection>-400.5 9</intersection>
<intersection>-378.5 10</intersection>
<intersection>-360 11</intersection>
<intersection>-341 12</intersection>
<intersection>-322.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>162.5,-456.5,165.5,-456.5</points>
<intersection>162.5 14</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162.5,-438,165.5,-438</points>
<intersection>162.5 15</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>162.5,-419,165.5,-419</points>
<intersection>162.5 16</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-400.5,165.5,-400.5</points>
<intersection>162.5 17</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>162.5,-378.5,165.5,-378.5</points>
<intersection>162.5 20</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>162.5,-360,165.5,-360</points>
<intersection>162.5 21</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>162.5,-341,165.5,-341</points>
<intersection>162.5 22</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>162.5,-322.5,165.5,-322.5</points>
<intersection>162.5 23</intersection>
<intersection>165.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>162.5,-457.5,162.5,-456.5</points>
<connection>
<GID>4635</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>162.5,-439,162.5,-438</points>
<connection>
<GID>4308</GID>
<name>OUT_0</name></connection>
<intersection>-438 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>162.5,-420,162.5,-419</points>
<connection>
<GID>4350</GID>
<name>OUT_0</name></connection>
<intersection>-419 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>162.5,-401.5,162.5,-400.5</points>
<connection>
<GID>4370</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>162.5,-379.5,162.5,-378.5</points>
<connection>
<GID>4491</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>162.5,-361,162.5,-360</points>
<connection>
<GID>4527</GID>
<name>OUT_0</name></connection>
<intersection>-360 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>162.5,-342,162.5,-341</points>
<connection>
<GID>4563</GID>
<name>OUT_0</name></connection>
<intersection>-341 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>162.5,-323.5,162.5,-322.5</points>
<connection>
<GID>4599</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-3857.5,205.5,-3850</points>
<connection>
<GID>219</GID>
<name>N_in1</name></connection>
<connection>
<GID>139</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-472,170.5,-307.5</points>
<connection>
<GID>4402</GID>
<name>N_in1</name></connection>
<connection>
<GID>4387</GID>
<name>N_in0</name></connection>
<intersection>-447.5 13</intersection>
<intersection>-429 12</intersection>
<intersection>-410 11</intersection>
<intersection>-391.5 10</intersection>
<intersection>-369.5 9</intersection>
<intersection>-351 8</intersection>
<intersection>-332 7</intersection>
<intersection>-313.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>170.5,-313.5,172.5,-313.5</points>
<connection>
<GID>4601</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>170.5,-332,172.5,-332</points>
<connection>
<GID>4565</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>170.5,-351,172.5,-351</points>
<connection>
<GID>4529</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>170.5,-369.5,172.5,-369.5</points>
<connection>
<GID>4493</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>170.5,-391.5,172.5,-391.5</points>
<connection>
<GID>4371</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>170.5,-410,172.5,-410</points>
<connection>
<GID>4352</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>170.5,-429,172.5,-429</points>
<connection>
<GID>4310</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>170.5,-447.5,172.5,-447.5</points>
<connection>
<GID>4637</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-3858,226.5,-3849.5</points>
<connection>
<GID>223</GID>
<name>N_in1</name></connection>
<connection>
<GID>140</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-471.5,188.5,-307.5</points>
<connection>
<GID>4403</GID>
<name>N_in1</name></connection>
<connection>
<GID>4389</GID>
<name>N_in0</name></connection>
<intersection>-456.5 16</intersection>
<intersection>-438 15</intersection>
<intersection>-419 14</intersection>
<intersection>-400.5 13</intersection>
<intersection>-378.5 12</intersection>
<intersection>-360 11</intersection>
<intersection>-341 10</intersection>
<intersection>-322.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>185.5,-322.5,188.5,-322.5</points>
<intersection>185.5 26</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>185.5,-341,188.5,-341</points>
<intersection>185.5 25</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>185.5,-360,188.5,-360</points>
<intersection>185.5 24</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185.5,-378.5,188.5,-378.5</points>
<intersection>185.5 23</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>185.5,-400.5,188.5,-400.5</points>
<intersection>185.5 20</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>185.5,-419,188.5,-419</points>
<intersection>185.5 19</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>185.5,-438,188.5,-438</points>
<intersection>185.5 18</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>185.5,-456.5,188.5,-456.5</points>
<intersection>185.5 17</intersection>
<intersection>188.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>185.5,-457.5,185.5,-456.5</points>
<connection>
<GID>4639</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>185.5,-439,185.5,-438</points>
<connection>
<GID>4312</GID>
<name>OUT_0</name></connection>
<intersection>-438 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>185.5,-420,185.5,-419</points>
<connection>
<GID>4353</GID>
<name>OUT_0</name></connection>
<intersection>-419 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>185.5,-401.5,185.5,-400.5</points>
<connection>
<GID>4372</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>185.5,-379.5,185.5,-378.5</points>
<connection>
<GID>4495</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>185.5,-361,185.5,-360</points>
<connection>
<GID>4531</GID>
<name>OUT_0</name></connection>
<intersection>-360 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>185.5,-342,185.5,-341</points>
<connection>
<GID>4567</GID>
<name>OUT_0</name></connection>
<intersection>-341 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>185.5,-323.5,185.5,-322.5</points>
<connection>
<GID>4603</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-3858,230,-3849.5</points>
<connection>
<GID>265</GID>
<name>N_in1</name></connection>
<connection>
<GID>141</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-471.5,193,-307.5</points>
<connection>
<GID>4404</GID>
<name>N_in1</name></connection>
<connection>
<GID>4388</GID>
<name>N_in0</name></connection>
<intersection>-447.5 13</intersection>
<intersection>-429 12</intersection>
<intersection>-410 11</intersection>
<intersection>-391.5 10</intersection>
<intersection>-369.5 9</intersection>
<intersection>-351 8</intersection>
<intersection>-332 7</intersection>
<intersection>-313.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>193,-313.5,197.5,-313.5</points>
<connection>
<GID>4605</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>193,-332,197.5,-332</points>
<connection>
<GID>4569</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>193,-351,197.5,-351</points>
<connection>
<GID>4533</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>193,-369.5,197.5,-369.5</points>
<connection>
<GID>4497</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>193,-391.5,197.5,-391.5</points>
<connection>
<GID>4373</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>193,-410,197.5,-410</points>
<connection>
<GID>4355</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>193,-429,197.5,-429</points>
<connection>
<GID>4314</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>193,-447.5,197.5,-447.5</points>
<connection>
<GID>4641</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-3859,251,-3849.5</points>
<connection>
<GID>225</GID>
<name>N_in1</name></connection>
<connection>
<GID>143</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-471,214,-308</points>
<connection>
<GID>4405</GID>
<name>N_in1</name></connection>
<connection>
<GID>4390</GID>
<name>N_in0</name></connection>
<intersection>-456.5 6</intersection>
<intersection>-438 7</intersection>
<intersection>-419 8</intersection>
<intersection>-400.5 9</intersection>
<intersection>-378.5 10</intersection>
<intersection>-360 11</intersection>
<intersection>-341 12</intersection>
<intersection>-322.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>210.5,-456.5,214,-456.5</points>
<intersection>210.5 14</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>210.5,-438,214,-438</points>
<intersection>210.5 15</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>210.5,-419,214,-419</points>
<intersection>210.5 16</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>210.5,-400.5,214,-400.5</points>
<intersection>210.5 17</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210.5,-378.5,214,-378.5</points>
<intersection>210.5 20</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>210.5,-360,214,-360</points>
<intersection>210.5 21</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>210.5,-341,214,-341</points>
<intersection>210.5 22</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>210.5,-322.5,214,-322.5</points>
<intersection>210.5 23</intersection>
<intersection>214 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>210.5,-457.5,210.5,-456.5</points>
<connection>
<GID>4643</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>210.5,-439,210.5,-438</points>
<connection>
<GID>4316</GID>
<name>OUT_0</name></connection>
<intersection>-438 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>210.5,-420,210.5,-419</points>
<connection>
<GID>4356</GID>
<name>OUT_0</name></connection>
<intersection>-419 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>210.5,-401.5,210.5,-400.5</points>
<connection>
<GID>4374</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>210.5,-379.5,210.5,-378.5</points>
<connection>
<GID>4499</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>210.5,-361,210.5,-360</points>
<connection>
<GID>4535</GID>
<name>OUT_0</name></connection>
<intersection>-360 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>210.5,-342,210.5,-341</points>
<connection>
<GID>4571</GID>
<name>OUT_0</name></connection>
<intersection>-341 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>210.5,-323.5,210.5,-322.5</points>
<connection>
<GID>4607</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-471,217.5,-308</points>
<connection>
<GID>4406</GID>
<name>N_in1</name></connection>
<connection>
<GID>4407</GID>
<name>N_in0</name></connection>
<intersection>-447.5 11</intersection>
<intersection>-429 10</intersection>
<intersection>-410 9</intersection>
<intersection>-391.5 7</intersection>
<intersection>-369.5 6</intersection>
<intersection>-351 5</intersection>
<intersection>-332 4</intersection>
<intersection>-313.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-313.5,220.5,-313.5</points>
<connection>
<GID>4609</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>217.5,-332,220.5,-332</points>
<connection>
<GID>4573</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-351,220.5,-351</points>
<connection>
<GID>4537</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>217.5,-369.5,220.5,-369.5</points>
<connection>
<GID>4501</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>217.5,-391.5,220.5,-391.5</points>
<connection>
<GID>4375</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>217.5,-410,220.5,-410</points>
<connection>
<GID>4357</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>217.5,-429,220.5,-429</points>
<connection>
<GID>4318</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>217.5,-447.5,220.5,-447.5</points>
<connection>
<GID>4645</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-471,238.5,-309</points>
<connection>
<GID>4408</GID>
<name>N_in1</name></connection>
<connection>
<GID>4391</GID>
<name>N_in0</name></connection>
<intersection>-456.5 11</intersection>
<intersection>-438 10</intersection>
<intersection>-419 9</intersection>
<intersection>-400.5 8</intersection>
<intersection>-378.5 7</intersection>
<intersection>-360 6</intersection>
<intersection>-341 5</intersection>
<intersection>-322.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>233.5,-322.5,238.5,-322.5</points>
<intersection>233.5 21</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>233.5,-341,238.5,-341</points>
<intersection>233.5 20</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>233.5,-360,238.5,-360</points>
<intersection>233.5 19</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>233.5,-378.5,238.5,-378.5</points>
<intersection>233.5 18</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>233.5,-400.5,238.5,-400.5</points>
<intersection>233.5 15</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>233.5,-419,238.5,-419</points>
<intersection>233.5 14</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>233.5,-438,238.5,-438</points>
<intersection>233.5 13</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>233.5,-456.5,238.5,-456.5</points>
<intersection>233.5 12</intersection>
<intersection>238.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>233.5,-457.5,233.5,-456.5</points>
<connection>
<GID>4647</GID>
<name>OUT_0</name></connection>
<intersection>-456.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>233.5,-439,233.5,-438</points>
<connection>
<GID>4320</GID>
<name>OUT_0</name></connection>
<intersection>-438 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>233.5,-420,233.5,-419</points>
<connection>
<GID>4358</GID>
<name>OUT_0</name></connection>
<intersection>-419 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>233.5,-401.5,233.5,-400.5</points>
<connection>
<GID>4376</GID>
<name>OUT_0</name></connection>
<intersection>-400.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>233.5,-379.5,233.5,-378.5</points>
<connection>
<GID>4503</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>233.5,-361,233.5,-360</points>
<connection>
<GID>4539</GID>
<name>OUT_0</name></connection>
<intersection>-360 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>233.5,-342,233.5,-341</points>
<connection>
<GID>4575</GID>
<name>OUT_0</name></connection>
<intersection>-341 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>233.5,-323.5,233.5,-322.5</points>
<connection>
<GID>4611</GID>
<name>OUT_0</name></connection>
<intersection>-322.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>3312</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-118.5,-315.5,28,-315.5</points>
<connection>
<GID>4577</GID>
<name>IN_0</name></connection>
<intersection>-118.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118.5,-467,-118.5,-315.5</points>
<connection>
<GID>4414</GID>
<name>OUT_15</name></connection>
<intersection>-325 4</intersection>
<intersection>-315.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118.5,-325,39.5,-325</points>
<connection>
<GID>4579</GID>
<name>IN_0</name></connection>
<intersection>-118.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3313</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-117.5,-334,28,-334</points>
<connection>
<GID>4541</GID>
<name>IN_0</name></connection>
<intersection>-117.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-117.5,-468,-117.5,-334</points>
<intersection>-468 6</intersection>
<intersection>-343.5 5</intersection>
<intersection>-334 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-117.5,-343.5,39.5,-343.5</points>
<connection>
<GID>4543</GID>
<name>IN_0</name></connection>
<intersection>-117.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118.5,-468,-117.5,-468</points>
<connection>
<GID>4414</GID>
<name>OUT_14</name></connection>
<intersection>-117.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3314</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-116.5,-353,28,-353</points>
<connection>
<GID>4505</GID>
<name>IN_0</name></connection>
<intersection>-116.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-116.5,-469,-116.5,-353</points>
<intersection>-469 6</intersection>
<intersection>-362.5 4</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-116.5,-362.5,39.5,-362.5</points>
<connection>
<GID>4507</GID>
<name>IN_0</name></connection>
<intersection>-116.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118.5,-469,-116.5,-469</points>
<connection>
<GID>4414</GID>
<name>OUT_13</name></connection>
<intersection>-116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3315</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-115.5,-371.5,28,-371.5</points>
<connection>
<GID>4445</GID>
<name>IN_0</name></connection>
<intersection>-115.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-115.5,-470,-115.5,-371.5</points>
<intersection>-470 5</intersection>
<intersection>-381 4</intersection>
<intersection>-371.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-115.5,-381,39.5,-381</points>
<connection>
<GID>4450</GID>
<name>IN_0</name></connection>
<intersection>-115.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-470,-115.5,-470</points>
<connection>
<GID>4414</GID>
<name>OUT_12</name></connection>
<intersection>-115.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114.5,-393.5,28,-393.5</points>
<connection>
<GID>4359</GID>
<name>IN_0</name></connection>
<intersection>-114.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114.5,-471,-114.5,-393.5</points>
<intersection>-471 6</intersection>
<intersection>-403 4</intersection>
<intersection>-393.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-114.5,-403,39,-403</points>
<connection>
<GID>4360</GID>
<name>IN_0</name></connection>
<intersection>-114.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118.5,-471,-114.5,-471</points>
<connection>
<GID>4414</GID>
<name>OUT_11</name></connection>
<intersection>-114.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,-412,28,-412</points>
<connection>
<GID>4323</GID>
<name>IN_0</name></connection>
<intersection>-113.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-113.5,-472,-113.5,-412</points>
<intersection>-472 5</intersection>
<intersection>-421.5 4</intersection>
<intersection>-412 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-113.5,-421.5,39,-421.5</points>
<connection>
<GID>4325</GID>
<name>IN_0</name></connection>
<intersection>-113.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-472,-113.5,-472</points>
<connection>
<GID>4414</GID>
<name>OUT_10</name></connection>
<intersection>-113.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-112.5,-431,28,-431</points>
<connection>
<GID>4649</GID>
<name>IN_0</name></connection>
<intersection>-112.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-112.5,-473,-112.5,-431</points>
<intersection>-473 5</intersection>
<intersection>-440.5 4</intersection>
<intersection>-431 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-112.5,-440.5,39,-440.5</points>
<connection>
<GID>4651</GID>
<name>IN_0</name></connection>
<intersection>-112.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-473,-112.5,-473</points>
<connection>
<GID>4414</GID>
<name>OUT_9</name></connection>
<intersection>-112.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-111.5,-449.5,28,-449.5</points>
<connection>
<GID>4613</GID>
<name>IN_0</name></connection>
<intersection>-111.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-111.5,-474,-111.5,-449.5</points>
<intersection>-474 5</intersection>
<intersection>-459 4</intersection>
<intersection>-449.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-111.5,-459,39,-459</points>
<connection>
<GID>4615</GID>
<name>IN_0</name></connection>
<intersection>-111.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-474,-111.5,-474</points>
<connection>
<GID>4414</GID>
<name>OUT_8</name></connection>
<intersection>-111.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-473,27,-308</points>
<connection>
<GID>4412</GID>
<name>N_in1</name></connection>
<connection>
<GID>4410</GID>
<name>N_in0</name></connection>
<intersection>-451.5 10</intersection>
<intersection>-433 9</intersection>
<intersection>-414 8</intersection>
<intersection>-395.5 7</intersection>
<intersection>-373.5 6</intersection>
<intersection>-355 5</intersection>
<intersection>-336 4</intersection>
<intersection>-317.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27,-317.5,28,-317.5</points>
<connection>
<GID>4577</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-336,28,-336</points>
<connection>
<GID>4541</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>27,-355,28,-355</points>
<connection>
<GID>4505</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-373.5,28,-373.5</points>
<connection>
<GID>4445</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27,-395.5,28,-395.5</points>
<connection>
<GID>4359</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>27,-414,28,-414</points>
<connection>
<GID>4323</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>27,-433,28,-433</points>
<connection>
<GID>4649</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>27,-451.5,28,-451.5</points>
<connection>
<GID>4613</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>3321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-473,37,-308</points>
<connection>
<GID>4411</GID>
<name>N_in1</name></connection>
<connection>
<GID>4409</GID>
<name>N_in0</name></connection>
<intersection>-461 3</intersection>
<intersection>-442.5 5</intersection>
<intersection>-423.5 7</intersection>
<intersection>-405 9</intersection>
<intersection>-383 11</intersection>
<intersection>-364.5 13</intersection>
<intersection>-345.5 15</intersection>
<intersection>-327 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>37,-461,39,-461</points>
<connection>
<GID>4615</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>37,-442.5,39,-442.5</points>
<connection>
<GID>4651</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>37,-423.5,39,-423.5</points>
<connection>
<GID>4325</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>37,-405,39,-405</points>
<connection>
<GID>4360</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>37,-383,39.5,-383</points>
<connection>
<GID>4450</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>37,-364.5,39.5,-364.5</points>
<connection>
<GID>4507</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>37,-345.5,39.5,-345.5</points>
<connection>
<GID>4543</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>37,-327,39.5,-327</points>
<connection>
<GID>4579</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>3322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-560.5,68.5,-560.5</points>
<connection>
<GID>4510</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-560.5,62.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-545,62.5,-545</points>
<connection>
<GID>4498</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-560.5,91.5,-560.5</points>
<connection>
<GID>4536</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-560.5,85.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-545,85.5,-545</points>
<connection>
<GID>4534</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-560.5,116.5,-560.5</points>
<connection>
<GID>4544</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-560.5,110.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-545,110.5,-545</points>
<connection>
<GID>4540</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-560.5,139.5,-560.5</points>
<connection>
<GID>4552</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-560.5,133.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-545,133.5,-545</points>
<connection>
<GID>4548</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3326</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-560.5,162.5,-560.5</points>
<connection>
<GID>4558</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-560.5,156.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-545,156.5,-545</points>
<connection>
<GID>4554</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-560.5,185.5,-560.5</points>
<connection>
<GID>4562</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-560.5,179.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-545,179.5,-545</points>
<connection>
<GID>4560</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-560.5,210.5,-560.5</points>
<connection>
<GID>4566</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-560.5,204.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-545,204.5,-545</points>
<connection>
<GID>4564</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-560.5,233.5,-560.5</points>
<connection>
<GID>4570</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-560.5,227.5,-545</points>
<intersection>-560.5 1</intersection>
<intersection>-545 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-545,227.5,-545</points>
<connection>
<GID>4568</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-548,220.5,-548</points>
<connection>
<GID>4568</GID>
<name>clock</name></connection>
<connection>
<GID>4564</GID>
<name>clock</name></connection>
<connection>
<GID>4560</GID>
<name>clock</name></connection>
<connection>
<GID>4554</GID>
<name>clock</name></connection>
<connection>
<GID>4548</GID>
<name>clock</name></connection>
<connection>
<GID>4540</GID>
<name>clock</name></connection>
<connection>
<GID>4534</GID>
<name>clock</name></connection>
<connection>
<GID>4498</GID>
<name>clock</name></connection>
<connection>
<GID>4492</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-557.5,231.5,-557.5</points>
<connection>
<GID>4570</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4566</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4562</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4558</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4552</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4544</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4536</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4510</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4494</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-542,68.5,-542</points>
<connection>
<GID>4578</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-542,62.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-526.5,62.5,-526.5</points>
<connection>
<GID>4576</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-542,91.5,-542</points>
<connection>
<GID>4582</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-542,85.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-526.5,85.5,-526.5</points>
<connection>
<GID>4580</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-542,116.5,-542</points>
<connection>
<GID>4586</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-542,110.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-526.5,110.5,-526.5</points>
<connection>
<GID>4584</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-542,139.5,-542</points>
<connection>
<GID>4590</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-542,133.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-526.5,133.5,-526.5</points>
<connection>
<GID>4588</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-542,162.5,-542</points>
<connection>
<GID>4594</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-542,156.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-526.5,156.5,-526.5</points>
<connection>
<GID>4592</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3337</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-542,185.5,-542</points>
<connection>
<GID>4598</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-542,179.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-526.5,179.5,-526.5</points>
<connection>
<GID>4596</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-542,210.5,-542</points>
<connection>
<GID>4602</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-542,204.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-526.5,204.5,-526.5</points>
<connection>
<GID>4600</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-542,233.5,-542</points>
<connection>
<GID>4606</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-542,227.5,-526.5</points>
<intersection>-542 1</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-526.5,227.5,-526.5</points>
<connection>
<GID>4604</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3340</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-529.5,220.5,-529.5</points>
<connection>
<GID>4604</GID>
<name>clock</name></connection>
<connection>
<GID>4600</GID>
<name>clock</name></connection>
<connection>
<GID>4596</GID>
<name>clock</name></connection>
<connection>
<GID>4592</GID>
<name>clock</name></connection>
<connection>
<GID>4588</GID>
<name>clock</name></connection>
<connection>
<GID>4584</GID>
<name>clock</name></connection>
<connection>
<GID>4580</GID>
<name>clock</name></connection>
<connection>
<GID>4576</GID>
<name>clock</name></connection>
<connection>
<GID>4572</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-539,231.5,-539</points>
<connection>
<GID>4606</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4602</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4598</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4594</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4590</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4586</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4582</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4578</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4574</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-523,68.5,-523</points>
<connection>
<GID>4614</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-523,62.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-507.5,62.5,-507.5</points>
<connection>
<GID>4612</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-523,91.5,-523</points>
<connection>
<GID>4618</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-523,85.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-507.5,85.5,-507.5</points>
<connection>
<GID>4616</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-523,116.5,-523</points>
<connection>
<GID>4622</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-523,110.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-507.5,110.5,-507.5</points>
<connection>
<GID>4620</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-523,139.5,-523</points>
<connection>
<GID>4626</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-523,133.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-507.5,133.5,-507.5</points>
<connection>
<GID>4624</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-523,162.5,-523</points>
<connection>
<GID>4630</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-523,156.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-507.5,156.5,-507.5</points>
<connection>
<GID>4628</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-523,185.5,-523</points>
<connection>
<GID>4634</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-523,179.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-507.5,179.5,-507.5</points>
<connection>
<GID>4632</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-523,210.5,-523</points>
<connection>
<GID>4638</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-523,204.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-507.5,204.5,-507.5</points>
<connection>
<GID>4636</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-523,233.5,-523</points>
<connection>
<GID>4642</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-523,227.5,-507.5</points>
<intersection>-523 1</intersection>
<intersection>-507.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-507.5,227.5,-507.5</points>
<connection>
<GID>4640</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-510.5,220.5,-510.5</points>
<connection>
<GID>4612</GID>
<name>clock</name></connection>
<connection>
<GID>4608</GID>
<name>OUT</name></connection>
<connection>
<GID>4640</GID>
<name>clock</name></connection>
<connection>
<GID>4636</GID>
<name>clock</name></connection>
<connection>
<GID>4632</GID>
<name>clock</name></connection>
<connection>
<GID>4628</GID>
<name>clock</name></connection>
<connection>
<GID>4624</GID>
<name>clock</name></connection>
<connection>
<GID>4620</GID>
<name>clock</name></connection>
<connection>
<GID>4616</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-520,231.5,-520</points>
<connection>
<GID>4610</GID>
<name>OUT</name></connection>
<connection>
<GID>4642</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4638</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4634</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4630</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4626</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4622</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4618</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4614</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-504.5,68.5,-504.5</points>
<connection>
<GID>4650</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-504.5,62.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-489,62.5,-489</points>
<connection>
<GID>4648</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-504.5,91.5,-504.5</points>
<connection>
<GID>4654</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-504.5,85.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-489,85.5,-489</points>
<connection>
<GID>4652</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-504.5,116.5,-504.5</points>
<connection>
<GID>4658</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-504.5,110.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-489,110.5,-489</points>
<connection>
<GID>4656</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3355</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-504.5,139.5,-504.5</points>
<connection>
<GID>4662</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-504.5,133.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-489,133.5,-489</points>
<connection>
<GID>4660</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3356</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-504.5,162.5,-504.5</points>
<connection>
<GID>4303</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-504.5,156.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-489,156.5,-489</points>
<connection>
<GID>4301</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-504.5,185.5,-504.5</points>
<connection>
<GID>4307</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-504.5,179.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-489,179.5,-489</points>
<connection>
<GID>4305</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3358</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-504.5,210.5,-504.5</points>
<connection>
<GID>4311</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-504.5,204.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-489,204.5,-489</points>
<connection>
<GID>4309</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3359</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-504.5,233.5,-504.5</points>
<connection>
<GID>4315</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-504.5,227.5,-489</points>
<intersection>-504.5 1</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-489,227.5,-489</points>
<connection>
<GID>4313</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-492,220.5,-492</points>
<connection>
<GID>4313</GID>
<name>clock</name></connection>
<connection>
<GID>4309</GID>
<name>clock</name></connection>
<connection>
<GID>4305</GID>
<name>clock</name></connection>
<connection>
<GID>4301</GID>
<name>clock</name></connection>
<connection>
<GID>4660</GID>
<name>clock</name></connection>
<connection>
<GID>4656</GID>
<name>clock</name></connection>
<connection>
<GID>4652</GID>
<name>clock</name></connection>
<connection>
<GID>4648</GID>
<name>clock</name></connection>
<connection>
<GID>4644</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3361</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-501.5,231.5,-501.5</points>
<connection>
<GID>4315</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4311</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4307</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4303</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4662</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4658</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4654</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4650</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4646</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3362</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-638.5,68.5,-638.5</points>
<connection>
<GID>4324</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-638.5,62.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-623,62.5,-623</points>
<connection>
<GID>4321</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-638.5,91.5,-638.5</points>
<connection>
<GID>4329</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-638.5,85.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-623,85.5,-623</points>
<connection>
<GID>4326</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-638.5,116.5,-638.5</points>
<connection>
<GID>4334</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-638.5,110.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-623,110.5,-623</points>
<connection>
<GID>4331</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-638.5,139.5,-638.5</points>
<connection>
<GID>4339</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-638.5,133.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-623,133.5,-623</points>
<connection>
<GID>4336</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3366</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-638.5,162.5,-638.5</points>
<connection>
<GID>4344</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-638.5,156.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-623,156.5,-623</points>
<connection>
<GID>4341</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3367</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-638.5,185.5,-638.5</points>
<connection>
<GID>4349</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-638.5,179.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-623,179.5,-623</points>
<connection>
<GID>4346</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-638.5,210.5,-638.5</points>
<connection>
<GID>4416</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-638.5,204.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-623,204.5,-623</points>
<connection>
<GID>4415</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-638.5,233.5,-638.5</points>
<connection>
<GID>4418</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-638.5,227.5,-623</points>
<intersection>-638.5 1</intersection>
<intersection>-623 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-623,227.5,-623</points>
<connection>
<GID>4417</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3370</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-626,220.5,-626</points>
<connection>
<GID>4417</GID>
<name>clock</name></connection>
<connection>
<GID>4415</GID>
<name>clock</name></connection>
<connection>
<GID>4346</GID>
<name>clock</name></connection>
<connection>
<GID>4341</GID>
<name>clock</name></connection>
<connection>
<GID>4336</GID>
<name>clock</name></connection>
<connection>
<GID>4331</GID>
<name>clock</name></connection>
<connection>
<GID>4326</GID>
<name>clock</name></connection>
<connection>
<GID>4321</GID>
<name>clock</name></connection>
<connection>
<GID>4317</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-635.5,231.5,-635.5</points>
<connection>
<GID>4418</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4416</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4349</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4344</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4339</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4334</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4329</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4324</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4319</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-620,68.5,-620</points>
<connection>
<GID>4422</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-620,62.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-604.5,62.5,-604.5</points>
<connection>
<GID>4421</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-620,91.5,-620</points>
<connection>
<GID>4424</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-620,85.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-604.5,85.5,-604.5</points>
<connection>
<GID>4423</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-620,116.5,-620</points>
<connection>
<GID>4426</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-620,110.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-604.5,110.5,-604.5</points>
<connection>
<GID>4425</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3375</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-620,139.5,-620</points>
<connection>
<GID>4428</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-620,133.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-604.5,133.5,-604.5</points>
<connection>
<GID>4427</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-620,162.5,-620</points>
<connection>
<GID>4430</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-620,156.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-604.5,156.5,-604.5</points>
<connection>
<GID>4429</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-620,185.5,-620</points>
<connection>
<GID>4432</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-620,179.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-604.5,179.5,-604.5</points>
<connection>
<GID>4431</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3378</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-620,210.5,-620</points>
<connection>
<GID>4434</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-620,204.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-604.5,204.5,-604.5</points>
<connection>
<GID>4433</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3379</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-620,233.5,-620</points>
<connection>
<GID>4436</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-620,227.5,-604.5</points>
<intersection>-620 1</intersection>
<intersection>-604.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-604.5,227.5,-604.5</points>
<connection>
<GID>4435</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-607.5,220.5,-607.5</points>
<connection>
<GID>4435</GID>
<name>clock</name></connection>
<connection>
<GID>4433</GID>
<name>clock</name></connection>
<connection>
<GID>4431</GID>
<name>clock</name></connection>
<connection>
<GID>4429</GID>
<name>clock</name></connection>
<connection>
<GID>4427</GID>
<name>clock</name></connection>
<connection>
<GID>4425</GID>
<name>clock</name></connection>
<connection>
<GID>4423</GID>
<name>clock</name></connection>
<connection>
<GID>4421</GID>
<name>clock</name></connection>
<connection>
<GID>4419</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3381</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-617,231.5,-617</points>
<connection>
<GID>4436</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4434</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4432</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4430</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4428</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4426</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4424</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4422</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4420</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3382</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-601,68.5,-601</points>
<connection>
<GID>4332</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-601,62.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-585.5,62.5,-585.5</points>
<connection>
<GID>4327</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3383</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-601,91.5,-601</points>
<connection>
<GID>4342</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-601,85.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-585.5,85.5,-585.5</points>
<connection>
<GID>4337</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3384</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-601,116.5,-601</points>
<connection>
<GID>4351</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-601,110.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-585.5,110.5,-585.5</points>
<connection>
<GID>4347</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-601,139.5,-601</points>
<connection>
<GID>4438</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-601,133.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-585.5,133.5,-585.5</points>
<connection>
<GID>4354</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-601,162.5,-601</points>
<connection>
<GID>4440</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-601,156.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-585.5,156.5,-585.5</points>
<connection>
<GID>4439</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3387</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-601,185.5,-601</points>
<connection>
<GID>4442</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-601,179.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-585.5,179.5,-585.5</points>
<connection>
<GID>4441</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-601,210.5,-601</points>
<connection>
<GID>4444</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-601,204.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-585.5,204.5,-585.5</points>
<connection>
<GID>4443</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-601,233.5,-601</points>
<connection>
<GID>4447</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-601,227.5,-585.5</points>
<intersection>-601 1</intersection>
<intersection>-585.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-585.5,227.5,-585.5</points>
<connection>
<GID>4446</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3390</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-588.5,220.5,-588.5</points>
<connection>
<GID>4446</GID>
<name>clock</name></connection>
<connection>
<GID>4443</GID>
<name>clock</name></connection>
<connection>
<GID>4441</GID>
<name>clock</name></connection>
<connection>
<GID>4439</GID>
<name>clock</name></connection>
<connection>
<GID>4437</GID>
<name>OUT</name></connection>
<connection>
<GID>4354</GID>
<name>clock</name></connection>
<connection>
<GID>4347</GID>
<name>clock</name></connection>
<connection>
<GID>4337</GID>
<name>clock</name></connection>
<connection>
<GID>4327</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3391</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-598,231.5,-598</points>
<connection>
<GID>4447</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4444</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4442</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4440</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4438</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4351</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4342</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4332</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4322</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-582.5,68.5,-582.5</points>
<connection>
<GID>4452</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,-582.5,62.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-567,62.5,-567</points>
<connection>
<GID>4451</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3393</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-582.5,91.5,-582.5</points>
<connection>
<GID>4454</GID>
<name>IN_0</name></connection>
<intersection>85.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-582.5,85.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-567,85.5,-567</points>
<connection>
<GID>4453</GID>
<name>OUT_0</name></connection>
<intersection>85.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-582.5,116.5,-582.5</points>
<connection>
<GID>4457</GID>
<name>IN_0</name></connection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-582.5,110.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-567,110.5,-567</points>
<connection>
<GID>4456</GID>
<name>OUT_0</name></connection>
<intersection>110.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3395</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-582.5,139.5,-582.5</points>
<connection>
<GID>4459</GID>
<name>IN_0</name></connection>
<intersection>133.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-582.5,133.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-567,133.5,-567</points>
<connection>
<GID>4458</GID>
<name>OUT_0</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-582.5,162.5,-582.5</points>
<connection>
<GID>4462</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-582.5,156.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-567,156.5,-567</points>
<connection>
<GID>4460</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-582.5,185.5,-582.5</points>
<connection>
<GID>4464</GID>
<name>IN_0</name></connection>
<intersection>179.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179.5,-582.5,179.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178.5,-567,179.5,-567</points>
<connection>
<GID>4463</GID>
<name>OUT_0</name></connection>
<intersection>179.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3398</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-582.5,210.5,-582.5</points>
<connection>
<GID>4466</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-582.5,204.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-567,204.5,-567</points>
<connection>
<GID>4465</GID>
<name>OUT_0</name></connection>
<intersection>204.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-582.5,233.5,-582.5</points>
<connection>
<GID>4468</GID>
<name>IN_0</name></connection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-582.5,227.5,-567</points>
<intersection>-582.5 1</intersection>
<intersection>-567 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-567,227.5,-567</points>
<connection>
<GID>4467</GID>
<name>OUT_0</name></connection>
<intersection>227.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3400</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-570,220.5,-570</points>
<connection>
<GID>4467</GID>
<name>clock</name></connection>
<connection>
<GID>4465</GID>
<name>clock</name></connection>
<connection>
<GID>4463</GID>
<name>clock</name></connection>
<connection>
<GID>4460</GID>
<name>clock</name></connection>
<connection>
<GID>4458</GID>
<name>clock</name></connection>
<connection>
<GID>4456</GID>
<name>clock</name></connection>
<connection>
<GID>4453</GID>
<name>clock</name></connection>
<connection>
<GID>4451</GID>
<name>clock</name></connection>
<connection>
<GID>4448</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-579.5,231.5,-579.5</points>
<connection>
<GID>4468</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4466</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4464</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4462</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4459</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4457</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4454</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4452</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4449</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-648.5,50,-483.5</points>
<connection>
<GID>4496</GID>
<name>N_in1</name></connection>
<connection>
<GID>4469</GID>
<name>N_in0</name></connection>
<intersection>-623 12</intersection>
<intersection>-604.5 11</intersection>
<intersection>-585.5 10</intersection>
<intersection>-567 9</intersection>
<intersection>-545 8</intersection>
<intersection>-526.5 7</intersection>
<intersection>-507.5 6</intersection>
<intersection>-489 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-489,55.5,-489</points>
<connection>
<GID>4648</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>50,-507.5,55.5,-507.5</points>
<connection>
<GID>4612</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>50,-526.5,55.5,-526.5</points>
<connection>
<GID>4576</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>50,-545,55.5,-545</points>
<connection>
<GID>4498</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>50,-567,55.5,-567</points>
<connection>
<GID>4451</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>50,-585.5,55.5,-585.5</points>
<connection>
<GID>4327</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>50,-604.5,55.5,-604.5</points>
<connection>
<GID>4421</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>50,-623,55.5,-623</points>
<connection>
<GID>4321</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>3403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-648,73,-483</points>
<connection>
<GID>4500</GID>
<name>N_in1</name></connection>
<connection>
<GID>4470</GID>
<name>N_in0</name></connection>
<intersection>-631.5 4</intersection>
<intersection>-613 5</intersection>
<intersection>-594 6</intersection>
<intersection>-575.5 7</intersection>
<intersection>-553.5 8</intersection>
<intersection>-535 9</intersection>
<intersection>-516 10</intersection>
<intersection>-497.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-631.5,73,-631.5</points>
<intersection>68.5 12</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68.5,-613,73,-613</points>
<intersection>68.5 14</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68.5,-594,73,-594</points>
<intersection>68.5 13</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68.5,-575.5,73,-575.5</points>
<intersection>68.5 15</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-553.5,73,-553.5</points>
<intersection>68.5 18</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68.5,-535,73,-535</points>
<intersection>68.5 19</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68.5,-516,73,-516</points>
<intersection>68.5 20</intersection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>68.5,-497.5,73,-497.5</points>
<intersection>68.5 21</intersection>
<intersection>73 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>68.5,-633,68.5,-631.5</points>
<connection>
<GID>4324</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>68.5,-595.5,68.5,-594</points>
<connection>
<GID>4332</GID>
<name>OUT_0</name></connection>
<intersection>-594 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>68.5,-614.5,68.5,-613</points>
<connection>
<GID>4422</GID>
<name>OUT_0</name></connection>
<intersection>-613 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>68.5,-577,68.5,-575.5</points>
<connection>
<GID>4452</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>68.5,-555,68.5,-553.5</points>
<connection>
<GID>4510</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>68.5,-536.5,68.5,-535</points>
<connection>
<GID>4578</GID>
<name>OUT_0</name></connection>
<intersection>-535 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>68.5,-517.5,68.5,-516</points>
<connection>
<GID>4614</GID>
<name>OUT_0</name></connection>
<intersection>-516 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>68.5,-499,68.5,-497.5</points>
<connection>
<GID>4650</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>3404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-648,76,-483.5</points>
<connection>
<GID>4502</GID>
<name>N_in1</name></connection>
<connection>
<GID>4471</GID>
<name>N_in0</name></connection>
<intersection>-623 10</intersection>
<intersection>-604.5 9</intersection>
<intersection>-585.5 8</intersection>
<intersection>-567 7</intersection>
<intersection>-545 6</intersection>
<intersection>-526.5 5</intersection>
<intersection>-507.5 4</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>76,-489,78.5,-489</points>
<connection>
<GID>4652</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>76,-507.5,78.5,-507.5</points>
<connection>
<GID>4616</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>76,-526.5,78.5,-526.5</points>
<connection>
<GID>4580</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>76,-545,78.5,-545</points>
<connection>
<GID>4534</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>76,-567,78.5,-567</points>
<connection>
<GID>4453</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>76,-585.5,78.5,-585.5</points>
<connection>
<GID>4337</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>76,-604.5,78.5,-604.5</points>
<connection>
<GID>4423</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>76,-623,78.5,-623</points>
<connection>
<GID>4326</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>3405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-648,95.5,-483</points>
<connection>
<GID>4504</GID>
<name>N_in1</name></connection>
<connection>
<GID>4472</GID>
<name>N_in0</name></connection>
<intersection>-631.5 6</intersection>
<intersection>-613 7</intersection>
<intersection>-594 8</intersection>
<intersection>-575.5 9</intersection>
<intersection>-553.5 10</intersection>
<intersection>-535 11</intersection>
<intersection>-516 12</intersection>
<intersection>-497.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91.5,-631.5,95.5,-631.5</points>
<intersection>91.5 14</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>91.5,-613,95.5,-613</points>
<intersection>91.5 16</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>91.5,-594,95.5,-594</points>
<intersection>91.5 15</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>91.5,-575.5,95.5,-575.5</points>
<intersection>91.5 17</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>91.5,-553.5,95.5,-553.5</points>
<intersection>91.5 20</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>91.5,-535,95.5,-535</points>
<intersection>91.5 21</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>91.5,-516,95.5,-516</points>
<intersection>91.5 22</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>91.5,-497.5,95.5,-497.5</points>
<intersection>91.5 23</intersection>
<intersection>95.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>91.5,-633,91.5,-631.5</points>
<connection>
<GID>4329</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>91.5,-595.5,91.5,-594</points>
<connection>
<GID>4342</GID>
<name>OUT_0</name></connection>
<intersection>-594 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>91.5,-614.5,91.5,-613</points>
<connection>
<GID>4424</GID>
<name>OUT_0</name></connection>
<intersection>-613 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>91.5,-577,91.5,-575.5</points>
<connection>
<GID>4454</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>91.5,-555,91.5,-553.5</points>
<connection>
<GID>4536</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>91.5,-536.5,91.5,-535</points>
<connection>
<GID>4582</GID>
<name>OUT_0</name></connection>
<intersection>-535 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>91.5,-517.5,91.5,-516</points>
<connection>
<GID>4618</GID>
<name>OUT_0</name></connection>
<intersection>-516 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>91.5,-499,91.5,-497.5</points>
<connection>
<GID>4654</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-648,99,-483</points>
<connection>
<GID>4506</GID>
<name>N_in1</name></connection>
<connection>
<GID>4473</GID>
<name>N_in0</name></connection>
<intersection>-623 13</intersection>
<intersection>-604.5 12</intersection>
<intersection>-585.5 11</intersection>
<intersection>-567 10</intersection>
<intersection>-545 9</intersection>
<intersection>-526.5 8</intersection>
<intersection>-507.5 7</intersection>
<intersection>-489 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>99,-489,103.5,-489</points>
<connection>
<GID>4656</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>99,-507.5,103.5,-507.5</points>
<connection>
<GID>4620</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>99,-526.5,103.5,-526.5</points>
<connection>
<GID>4584</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>99,-545,103.5,-545</points>
<connection>
<GID>4540</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>99,-567,103.5,-567</points>
<connection>
<GID>4456</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>99,-585.5,103.5,-585.5</points>
<connection>
<GID>4347</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>99,-604.5,103.5,-604.5</points>
<connection>
<GID>4425</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>99,-623,103.5,-623</points>
<connection>
<GID>4331</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>3407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-648,120,-483.5</points>
<connection>
<GID>4508</GID>
<name>N_in1</name></connection>
<connection>
<GID>4474</GID>
<name>N_in0</name></connection>
<intersection>-631.5 6</intersection>
<intersection>-613 7</intersection>
<intersection>-594 8</intersection>
<intersection>-575.5 9</intersection>
<intersection>-553.5 10</intersection>
<intersection>-535 11</intersection>
<intersection>-516 12</intersection>
<intersection>-497.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116.5,-631.5,120,-631.5</points>
<intersection>116.5 14</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116.5,-613,120,-613</points>
<intersection>116.5 16</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>116.5,-594,120,-594</points>
<intersection>116.5 15</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116.5,-575.5,120,-575.5</points>
<intersection>116.5 17</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116.5,-553.5,120,-553.5</points>
<intersection>116.5 20</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>116.5,-535,120,-535</points>
<intersection>116.5 21</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>116.5,-516,120,-516</points>
<intersection>116.5 22</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>116.5,-497.5,120,-497.5</points>
<intersection>116.5 23</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>116.5,-633,116.5,-631.5</points>
<connection>
<GID>4334</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>116.5,-595.5,116.5,-594</points>
<connection>
<GID>4351</GID>
<name>OUT_0</name></connection>
<intersection>-594 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>116.5,-614.5,116.5,-613</points>
<connection>
<GID>4426</GID>
<name>OUT_0</name></connection>
<intersection>-613 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>116.5,-577,116.5,-575.5</points>
<connection>
<GID>4457</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>116.5,-555,116.5,-553.5</points>
<connection>
<GID>4544</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>116.5,-536.5,116.5,-535</points>
<connection>
<GID>4586</GID>
<name>OUT_0</name></connection>
<intersection>-535 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>116.5,-517.5,116.5,-516</points>
<connection>
<GID>4622</GID>
<name>OUT_0</name></connection>
<intersection>-516 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>116.5,-499,116.5,-497.5</points>
<connection>
<GID>4658</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-648,124,-483</points>
<connection>
<GID>4512</GID>
<name>N_in1</name></connection>
<connection>
<GID>4475</GID>
<name>N_in0</name></connection>
<intersection>-623 13</intersection>
<intersection>-604.5 12</intersection>
<intersection>-585.5 11</intersection>
<intersection>-567 10</intersection>
<intersection>-545 9</intersection>
<intersection>-526.5 8</intersection>
<intersection>-507.5 7</intersection>
<intersection>-489 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>124,-489,126.5,-489</points>
<connection>
<GID>4660</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>124,-507.5,126.5,-507.5</points>
<connection>
<GID>4624</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>124,-526.5,126.5,-526.5</points>
<connection>
<GID>4588</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>124,-545,126.5,-545</points>
<connection>
<GID>4548</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>124,-567,126.5,-567</points>
<connection>
<GID>4458</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>124,-585.5,126.5,-585.5</points>
<connection>
<GID>4354</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>124,-604.5,126.5,-604.5</points>
<connection>
<GID>4427</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>124,-623,126.5,-623</points>
<connection>
<GID>4336</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>3409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-648,142.5,-483</points>
<connection>
<GID>4514</GID>
<name>N_in1</name></connection>
<connection>
<GID>4476</GID>
<name>N_in0</name></connection>
<intersection>-631.5 6</intersection>
<intersection>-613 7</intersection>
<intersection>-594 8</intersection>
<intersection>-575.5 9</intersection>
<intersection>-553.5 10</intersection>
<intersection>-535 11</intersection>
<intersection>-516 12</intersection>
<intersection>-497.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139.5,-631.5,142.5,-631.5</points>
<intersection>139.5 14</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139.5,-613,142.5,-613</points>
<intersection>139.5 15</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>139.5,-594,142.5,-594</points>
<intersection>139.5 16</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>139.5,-575.5,142.5,-575.5</points>
<intersection>139.5 17</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>139.5,-553.5,142.5,-553.5</points>
<intersection>139.5 20</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139.5,-535,142.5,-535</points>
<intersection>139.5 21</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>139.5,-516,142.5,-516</points>
<intersection>139.5 22</intersection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>139.5,-497.5,142.5,-497.5</points>
<intersection>139.5 23</intersection>
<intersection>142.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>139.5,-633,139.5,-631.5</points>
<connection>
<GID>4339</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>139.5,-614.5,139.5,-613</points>
<connection>
<GID>4428</GID>
<name>OUT_0</name></connection>
<intersection>-613 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>139.5,-595.5,139.5,-594</points>
<connection>
<GID>4438</GID>
<name>OUT_0</name></connection>
<intersection>-594 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>139.5,-577,139.5,-575.5</points>
<connection>
<GID>4459</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>139.5,-555,139.5,-553.5</points>
<connection>
<GID>4552</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>139.5,-536.5,139.5,-535</points>
<connection>
<GID>4590</GID>
<name>OUT_0</name></connection>
<intersection>-535 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>139.5,-517.5,139.5,-516</points>
<connection>
<GID>4626</GID>
<name>OUT_0</name></connection>
<intersection>-516 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>139.5,-499,139.5,-497.5</points>
<connection>
<GID>4662</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-648,146.5,-483</points>
<connection>
<GID>4516</GID>
<name>N_in1</name></connection>
<connection>
<GID>4478</GID>
<name>N_in0</name></connection>
<intersection>-623 13</intersection>
<intersection>-604.5 12</intersection>
<intersection>-585.5 11</intersection>
<intersection>-567 10</intersection>
<intersection>-545 9</intersection>
<intersection>-526.5 8</intersection>
<intersection>-507.5 7</intersection>
<intersection>-489 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>146.5,-489,149.5,-489</points>
<connection>
<GID>4301</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>146.5,-507.5,149.5,-507.5</points>
<connection>
<GID>4628</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>146.5,-526.5,149.5,-526.5</points>
<connection>
<GID>4592</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>146.5,-545,149.5,-545</points>
<connection>
<GID>4554</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>146.5,-567,149.5,-567</points>
<connection>
<GID>4460</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>146.5,-585.5,149.5,-585.5</points>
<connection>
<GID>4439</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>146.5,-604.5,149.5,-604.5</points>
<connection>
<GID>4429</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>146.5,-623,149.5,-623</points>
<connection>
<GID>4341</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-647.5,165.5,-483</points>
<connection>
<GID>4518</GID>
<name>N_in1</name></connection>
<connection>
<GID>4480</GID>
<name>N_in0</name></connection>
<intersection>-631.5 6</intersection>
<intersection>-613 7</intersection>
<intersection>-594 8</intersection>
<intersection>-575.5 9</intersection>
<intersection>-553.5 10</intersection>
<intersection>-535 11</intersection>
<intersection>-516 12</intersection>
<intersection>-497.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>162.5,-631.5,165.5,-631.5</points>
<intersection>162.5 15</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162.5,-613,165.5,-613</points>
<intersection>162.5 16</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>162.5,-594,165.5,-594</points>
<intersection>162.5 17</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-575.5,165.5,-575.5</points>
<intersection>162.5 18</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>162.5,-553.5,165.5,-553.5</points>
<intersection>162.5 21</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>162.5,-535,165.5,-535</points>
<intersection>162.5 22</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>162.5,-516,165.5,-516</points>
<intersection>162.5 23</intersection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>162.5,-497.5,165.5,-497.5</points>
<intersection>162.5 14</intersection>
<intersection>165.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>162.5,-499,162.5,-497.5</points>
<connection>
<GID>4303</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>162.5,-633,162.5,-631.5</points>
<connection>
<GID>4344</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>162.5,-614.5,162.5,-613</points>
<connection>
<GID>4430</GID>
<name>OUT_0</name></connection>
<intersection>-613 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>162.5,-595.5,162.5,-594</points>
<connection>
<GID>4440</GID>
<name>OUT_0</name></connection>
<intersection>-594 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>162.5,-577,162.5,-575.5</points>
<connection>
<GID>4462</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>162.5,-555,162.5,-553.5</points>
<connection>
<GID>4558</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>162.5,-536.5,162.5,-535</points>
<connection>
<GID>4594</GID>
<name>OUT_0</name></connection>
<intersection>-535 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>162.5,-517.5,162.5,-516</points>
<connection>
<GID>4630</GID>
<name>OUT_0</name></connection>
<intersection>-516 12</intersection></vsegment></shape></wire>
<wire>
<ID>3412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-647.5,170.5,-483</points>
<connection>
<GID>4520</GID>
<name>N_in1</name></connection>
<connection>
<GID>4482</GID>
<name>N_in0</name></connection>
<intersection>-623 13</intersection>
<intersection>-604.5 12</intersection>
<intersection>-585.5 11</intersection>
<intersection>-567 10</intersection>
<intersection>-545 9</intersection>
<intersection>-526.5 8</intersection>
<intersection>-507.5 7</intersection>
<intersection>-489 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>170.5,-489,172.5,-489</points>
<connection>
<GID>4305</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>170.5,-507.5,172.5,-507.5</points>
<connection>
<GID>4632</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>170.5,-526.5,172.5,-526.5</points>
<connection>
<GID>4596</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>170.5,-545,172.5,-545</points>
<connection>
<GID>4560</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>170.5,-567,172.5,-567</points>
<connection>
<GID>4463</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>170.5,-585.5,172.5,-585.5</points>
<connection>
<GID>4441</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>170.5,-604.5,172.5,-604.5</points>
<connection>
<GID>4431</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>170.5,-623,172.5,-623</points>
<connection>
<GID>4346</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-647,188.5,-483</points>
<connection>
<GID>4522</GID>
<name>N_in1</name></connection>
<connection>
<GID>4486</GID>
<name>N_in0</name></connection>
<intersection>-631.5 16</intersection>
<intersection>-613 15</intersection>
<intersection>-594 14</intersection>
<intersection>-575.5 13</intersection>
<intersection>-553.5 12</intersection>
<intersection>-535 11</intersection>
<intersection>-516 10</intersection>
<intersection>-497.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>185.5,-497.5,188.5,-497.5</points>
<intersection>185.5 17</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>185.5,-516,188.5,-516</points>
<intersection>185.5 26</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>185.5,-535,188.5,-535</points>
<intersection>185.5 25</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185.5,-553.5,188.5,-553.5</points>
<intersection>185.5 24</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>185.5,-575.5,188.5,-575.5</points>
<intersection>185.5 21</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>185.5,-594,188.5,-594</points>
<intersection>185.5 20</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>185.5,-613,188.5,-613</points>
<intersection>185.5 19</intersection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>185.5,-631.5,188.5,-631.5</points>
<intersection>185.5 18</intersection>
<intersection>188.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>185.5,-499,185.5,-497.5</points>
<connection>
<GID>4307</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>185.5,-633,185.5,-631.5</points>
<connection>
<GID>4349</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>185.5,-614.5,185.5,-613</points>
<connection>
<GID>4432</GID>
<name>OUT_0</name></connection>
<intersection>-613 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>185.5,-595.5,185.5,-594</points>
<connection>
<GID>4442</GID>
<name>OUT_0</name></connection>
<intersection>-594 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>185.5,-577,185.5,-575.5</points>
<connection>
<GID>4464</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>185.5,-555,185.5,-553.5</points>
<connection>
<GID>4562</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>185.5,-536.5,185.5,-535</points>
<connection>
<GID>4598</GID>
<name>OUT_0</name></connection>
<intersection>-535 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>185.5,-517.5,185.5,-516</points>
<connection>
<GID>4634</GID>
<name>OUT_0</name></connection>
<intersection>-516 10</intersection></vsegment></shape></wire>
<wire>
<ID>3414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-647,193,-483</points>
<connection>
<GID>4524</GID>
<name>N_in1</name></connection>
<connection>
<GID>4484</GID>
<name>N_in0</name></connection>
<intersection>-623 13</intersection>
<intersection>-604.5 12</intersection>
<intersection>-585.5 11</intersection>
<intersection>-567 10</intersection>
<intersection>-545 9</intersection>
<intersection>-526.5 8</intersection>
<intersection>-507.5 7</intersection>
<intersection>-489 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>193,-489,197.5,-489</points>
<connection>
<GID>4309</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>193,-507.5,197.5,-507.5</points>
<connection>
<GID>4636</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>193,-526.5,197.5,-526.5</points>
<connection>
<GID>4600</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>193,-545,197.5,-545</points>
<connection>
<GID>4564</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>193,-567,197.5,-567</points>
<connection>
<GID>4465</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>193,-585.5,197.5,-585.5</points>
<connection>
<GID>4443</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>193,-604.5,197.5,-604.5</points>
<connection>
<GID>4433</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>193,-623,197.5,-623</points>
<connection>
<GID>4415</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>3415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-646.5,214,-483.5</points>
<connection>
<GID>4526</GID>
<name>N_in1</name></connection>
<connection>
<GID>4488</GID>
<name>N_in0</name></connection>
<intersection>-631.5 6</intersection>
<intersection>-613 7</intersection>
<intersection>-594 8</intersection>
<intersection>-575.5 9</intersection>
<intersection>-553.5 10</intersection>
<intersection>-535 11</intersection>
<intersection>-516 12</intersection>
<intersection>-497.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>210.5,-631.5,214,-631.5</points>
<intersection>210.5 15</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>210.5,-613,214,-613</points>
<intersection>210.5 16</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>210.5,-594,214,-594</points>
<intersection>210.5 17</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>210.5,-575.5,214,-575.5</points>
<intersection>210.5 18</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210.5,-553.5,214,-553.5</points>
<intersection>210.5 21</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>210.5,-535,214,-535</points>
<intersection>210.5 22</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>210.5,-516,214,-516</points>
<intersection>210.5 23</intersection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>210.5,-497.5,214,-497.5</points>
<intersection>210.5 14</intersection>
<intersection>214 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>210.5,-499,210.5,-497.5</points>
<connection>
<GID>4311</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>210.5,-633,210.5,-631.5</points>
<connection>
<GID>4416</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>210.5,-614.5,210.5,-613</points>
<connection>
<GID>4434</GID>
<name>OUT_0</name></connection>
<intersection>-613 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>210.5,-595.5,210.5,-594</points>
<connection>
<GID>4444</GID>
<name>OUT_0</name></connection>
<intersection>-594 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>210.5,-577,210.5,-575.5</points>
<connection>
<GID>4466</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>210.5,-555,210.5,-553.5</points>
<connection>
<GID>4566</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>210.5,-536.5,210.5,-535</points>
<connection>
<GID>4602</GID>
<name>OUT_0</name></connection>
<intersection>-535 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>210.5,-517.5,210.5,-516</points>
<connection>
<GID>4638</GID>
<name>OUT_0</name></connection>
<intersection>-516 12</intersection></vsegment></shape></wire>
<wire>
<ID>3416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-646.5,217.5,-483.5</points>
<connection>
<GID>4528</GID>
<name>N_in1</name></connection>
<connection>
<GID>4530</GID>
<name>N_in0</name></connection>
<intersection>-623 11</intersection>
<intersection>-604.5 10</intersection>
<intersection>-585.5 9</intersection>
<intersection>-567 7</intersection>
<intersection>-545 6</intersection>
<intersection>-526.5 5</intersection>
<intersection>-507.5 4</intersection>
<intersection>-489 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217.5,-489,220.5,-489</points>
<connection>
<GID>4313</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>217.5,-507.5,220.5,-507.5</points>
<connection>
<GID>4640</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217.5,-526.5,220.5,-526.5</points>
<connection>
<GID>4604</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>217.5,-545,220.5,-545</points>
<connection>
<GID>4568</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>217.5,-567,220.5,-567</points>
<connection>
<GID>4467</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>217.5,-585.5,220.5,-585.5</points>
<connection>
<GID>4446</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>217.5,-604.5,220.5,-604.5</points>
<connection>
<GID>4435</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>217.5,-623,220.5,-623</points>
<connection>
<GID>4417</GID>
<name>IN_0</name></connection>
<intersection>217.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-646.5,238.5,-484.5</points>
<connection>
<GID>4532</GID>
<name>N_in1</name></connection>
<connection>
<GID>4490</GID>
<name>N_in0</name></connection>
<intersection>-631.5 11</intersection>
<intersection>-613 10</intersection>
<intersection>-594 9</intersection>
<intersection>-575.5 8</intersection>
<intersection>-553.5 7</intersection>
<intersection>-535 6</intersection>
<intersection>-516 5</intersection>
<intersection>-497.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>233.5,-497.5,238.5,-497.5</points>
<intersection>233.5 12</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>233.5,-516,238.5,-516</points>
<intersection>233.5 21</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>233.5,-535,238.5,-535</points>
<intersection>233.5 20</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>233.5,-553.5,238.5,-553.5</points>
<intersection>233.5 19</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>233.5,-575.5,238.5,-575.5</points>
<intersection>233.5 16</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>233.5,-594,238.5,-594</points>
<intersection>233.5 15</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>233.5,-613,238.5,-613</points>
<intersection>233.5 14</intersection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>233.5,-631.5,238.5,-631.5</points>
<intersection>233.5 13</intersection>
<intersection>238.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>233.5,-499,233.5,-497.5</points>
<connection>
<GID>4315</GID>
<name>OUT_0</name></connection>
<intersection>-497.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>233.5,-633,233.5,-631.5</points>
<connection>
<GID>4418</GID>
<name>OUT_0</name></connection>
<intersection>-631.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>233.5,-614.5,233.5,-613</points>
<connection>
<GID>4436</GID>
<name>OUT_0</name></connection>
<intersection>-613 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>233.5,-595.5,233.5,-594</points>
<connection>
<GID>4447</GID>
<name>OUT_0</name></connection>
<intersection>-594 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>233.5,-577,233.5,-575.5</points>
<connection>
<GID>4468</GID>
<name>OUT_0</name></connection>
<intersection>-575.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>233.5,-555,233.5,-553.5</points>
<connection>
<GID>4570</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>233.5,-536.5,233.5,-535</points>
<connection>
<GID>4606</GID>
<name>OUT_0</name></connection>
<intersection>-535 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>233.5,-517.5,233.5,-516</points>
<connection>
<GID>4642</GID>
<name>OUT_0</name></connection>
<intersection>-516 5</intersection></vsegment></shape></wire>
<wire>
<ID>3418</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-111.5,-491,28,-491</points>
<connection>
<GID>4644</GID>
<name>IN_0</name></connection>
<intersection>-111.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-111.5,-500.5,-111.5,-475</points>
<intersection>-500.5 4</intersection>
<intersection>-491 2</intersection>
<intersection>-475 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-111.5,-500.5,39.5,-500.5</points>
<connection>
<GID>4646</GID>
<name>IN_0</name></connection>
<intersection>-111.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118.5,-475,-111.5,-475</points>
<connection>
<GID>4414</GID>
<name>OUT_7</name></connection>
<intersection>-111.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3419</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-112.5,-509.5,28,-509.5</points>
<connection>
<GID>4608</GID>
<name>IN_0</name></connection>
<intersection>-112.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-112.5,-519,-112.5,-476</points>
<intersection>-519 5</intersection>
<intersection>-509.5 2</intersection>
<intersection>-476 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-112.5,-519,39.5,-519</points>
<connection>
<GID>4610</GID>
<name>IN_0</name></connection>
<intersection>-112.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118.5,-476,-112.5,-476</points>
<connection>
<GID>4414</GID>
<name>OUT_6</name></connection>
<intersection>-112.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3420</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-113.5,-528.5,28,-528.5</points>
<connection>
<GID>4572</GID>
<name>IN_0</name></connection>
<intersection>-113.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-113.5,-538,-113.5,-477</points>
<intersection>-538 4</intersection>
<intersection>-528.5 2</intersection>
<intersection>-477 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-113.5,-538,39.5,-538</points>
<connection>
<GID>4574</GID>
<name>IN_0</name></connection>
<intersection>-113.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118.5,-477,-113.5,-477</points>
<connection>
<GID>4414</GID>
<name>OUT_5</name></connection>
<intersection>-113.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3421</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-114.5,-547,28,-547</points>
<connection>
<GID>4492</GID>
<name>IN_0</name></connection>
<intersection>-114.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114.5,-556.5,-114.5,-478</points>
<intersection>-556.5 4</intersection>
<intersection>-547 2</intersection>
<intersection>-478 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-114.5,-556.5,39.5,-556.5</points>
<connection>
<GID>4494</GID>
<name>IN_0</name></connection>
<intersection>-114.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-478,-114.5,-478</points>
<connection>
<GID>4414</GID>
<name>OUT_4</name></connection>
<intersection>-114.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-569,28,-569</points>
<connection>
<GID>4448</GID>
<name>IN_0</name></connection>
<intersection>-115.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-115.5,-578.5,-115.5,-479</points>
<intersection>-578.5 4</intersection>
<intersection>-569 1</intersection>
<intersection>-479 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-115.5,-578.5,39,-578.5</points>
<connection>
<GID>4449</GID>
<name>IN_0</name></connection>
<intersection>-115.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-479,-115.5,-479</points>
<connection>
<GID>4414</GID>
<name>OUT_3</name></connection>
<intersection>-115.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116.5,-587.5,28,-587.5</points>
<connection>
<GID>4437</GID>
<name>IN_0</name></connection>
<intersection>-116.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-116.5,-597,-116.5,-480</points>
<intersection>-597 4</intersection>
<intersection>-587.5 1</intersection>
<intersection>-480 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-116.5,-597,39,-597</points>
<connection>
<GID>4322</GID>
<name>IN_0</name></connection>
<intersection>-116.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-480,-116.5,-480</points>
<connection>
<GID>4414</GID>
<name>OUT_2</name></connection>
<intersection>-116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-117.5,-606.5,28,-606.5</points>
<connection>
<GID>4419</GID>
<name>IN_0</name></connection>
<intersection>-117.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117.5,-616,-117.5,-481</points>
<intersection>-616 4</intersection>
<intersection>-606.5 1</intersection>
<intersection>-481 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117.5,-616,39,-616</points>
<connection>
<GID>4420</GID>
<name>IN_0</name></connection>
<intersection>-117.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-481,-117.5,-481</points>
<connection>
<GID>4414</GID>
<name>OUT_1</name></connection>
<intersection>-117.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-625,28,-625</points>
<connection>
<GID>4317</GID>
<name>IN_0</name></connection>
<intersection>-118.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118.5,-634.5,-118.5,-482</points>
<connection>
<GID>4414</GID>
<name>OUT_0</name></connection>
<intersection>-634.5 4</intersection>
<intersection>-625 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118.5,-634.5,39,-634.5</points>
<connection>
<GID>4319</GID>
<name>IN_0</name></connection>
<intersection>-118.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-648.5,27,-483.5</points>
<connection>
<GID>4550</GID>
<name>N_in1</name></connection>
<connection>
<GID>4542</GID>
<name>N_in0</name></connection>
<intersection>-627 10</intersection>
<intersection>-608.5 9</intersection>
<intersection>-589.5 8</intersection>
<intersection>-571 7</intersection>
<intersection>-549 6</intersection>
<intersection>-530.5 5</intersection>
<intersection>-511.5 4</intersection>
<intersection>-493 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27,-493,28,-493</points>
<connection>
<GID>4644</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-511.5,28,-511.5</points>
<connection>
<GID>4608</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>27,-530.5,28,-530.5</points>
<connection>
<GID>4572</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-549,28,-549</points>
<connection>
<GID>4492</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27,-571,28,-571</points>
<connection>
<GID>4448</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>27,-589.5,28,-589.5</points>
<connection>
<GID>4437</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>27,-608.5,28,-608.5</points>
<connection>
<GID>4419</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>27,-627,28,-627</points>
<connection>
<GID>4317</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>3427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-648.5,37,-483.5</points>
<connection>
<GID>4546</GID>
<name>N_in1</name></connection>
<connection>
<GID>4538</GID>
<name>N_in0</name></connection>
<intersection>-636.5 3</intersection>
<intersection>-618 5</intersection>
<intersection>-599 7</intersection>
<intersection>-580.5 9</intersection>
<intersection>-558.5 11</intersection>
<intersection>-540 13</intersection>
<intersection>-521 15</intersection>
<intersection>-502.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>37,-636.5,39,-636.5</points>
<connection>
<GID>4319</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>37,-618,39,-618</points>
<connection>
<GID>4420</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>37,-599,39,-599</points>
<connection>
<GID>4322</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>37,-580.5,39,-580.5</points>
<connection>
<GID>4449</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>37,-558.5,39.5,-558.5</points>
<connection>
<GID>4494</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>37,-540,39.5,-540</points>
<connection>
<GID>4574</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>37,-521,39.5,-521</points>
<connection>
<GID>4610</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>37,-502.5,39.5,-502.5</points>
<connection>
<GID>4646</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>3428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-481.5,27,-475</points>
<connection>
<GID>4542</GID>
<name>N_in1</name></connection>
<connection>
<GID>4412</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-481.5,37,-475</points>
<connection>
<GID>4538</GID>
<name>N_in1</name></connection>
<connection>
<GID>4411</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-481.5,50,-475</points>
<connection>
<GID>4469</GID>
<name>N_in1</name></connection>
<connection>
<GID>4392</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-481,73,-474.5</points>
<connection>
<GID>4470</GID>
<name>N_in1</name></connection>
<connection>
<GID>4393</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-481.5,76,-474.5</points>
<connection>
<GID>4471</GID>
<name>N_in1</name></connection>
<connection>
<GID>4394</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-481,95.5,-474.5</points>
<connection>
<GID>4472</GID>
<name>N_in1</name></connection>
<connection>
<GID>4395</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-481,99,-474.5</points>
<connection>
<GID>4473</GID>
<name>N_in1</name></connection>
<connection>
<GID>4396</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-481.5,120,-474.5</points>
<connection>
<GID>4474</GID>
<name>N_in1</name></connection>
<connection>
<GID>4397</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-481,124,-474.5</points>
<connection>
<GID>4475</GID>
<name>N_in1</name></connection>
<connection>
<GID>4398</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-481,142.5,-474.5</points>
<connection>
<GID>4476</GID>
<name>N_in1</name></connection>
<connection>
<GID>4399</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-481,146.5,-474.5</points>
<connection>
<GID>4478</GID>
<name>N_in1</name></connection>
<connection>
<GID>4400</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-481,165.5,-474</points>
<connection>
<GID>4480</GID>
<name>N_in1</name></connection>
<connection>
<GID>4401</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-481,170.5,-474</points>
<connection>
<GID>4482</GID>
<name>N_in1</name></connection>
<connection>
<GID>4402</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-481,188.5,-473.5</points>
<connection>
<GID>4486</GID>
<name>N_in1</name></connection>
<connection>
<GID>4403</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-481,193,-473.5</points>
<connection>
<GID>4484</GID>
<name>N_in1</name></connection>
<connection>
<GID>4404</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-481.5,214,-473</points>
<connection>
<GID>4488</GID>
<name>N_in1</name></connection>
<connection>
<GID>4405</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-481.5,217.5,-473</points>
<connection>
<GID>4530</GID>
<name>N_in1</name></connection>
<connection>
<GID>4406</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-482.5,238.5,-473</points>
<connection>
<GID>4490</GID>
<name>N_in1</name></connection>
<connection>
<GID>4408</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>3906</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-755.5,66,-755.5</points>
<connection>
<GID>5589</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-755.5,60,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-740,60,-740</points>
<connection>
<GID>5583</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3907</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-755.5,89,-755.5</points>
<connection>
<GID>5607</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-755.5,83,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-740,83,-740</points>
<connection>
<GID>5605</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3908</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-755.5,114,-755.5</points>
<connection>
<GID>5611</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-755.5,108,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-740,108,-740</points>
<connection>
<GID>5609</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3909</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-755.5,137,-755.5</points>
<connection>
<GID>5615</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-755.5,131,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-740,131,-740</points>
<connection>
<GID>5613</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3910</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-755.5,160,-755.5</points>
<connection>
<GID>5619</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-755.5,154,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-740,154,-740</points>
<connection>
<GID>5617</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3911</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-755.5,183,-755.5</points>
<connection>
<GID>5623</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-755.5,177,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-740,177,-740</points>
<connection>
<GID>5621</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3912</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-755.5,208,-755.5</points>
<connection>
<GID>5627</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-755.5,202,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-740,202,-740</points>
<connection>
<GID>5625</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3913</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-755.5,231,-755.5</points>
<connection>
<GID>5631</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-755.5,225,-740</points>
<intersection>-755.5 1</intersection>
<intersection>-740 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-740,225,-740</points>
<connection>
<GID>5629</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3914</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-743,218,-743</points>
<connection>
<GID>5629</GID>
<name>clock</name></connection>
<connection>
<GID>5625</GID>
<name>clock</name></connection>
<connection>
<GID>5621</GID>
<name>clock</name></connection>
<connection>
<GID>5617</GID>
<name>clock</name></connection>
<connection>
<GID>5613</GID>
<name>clock</name></connection>
<connection>
<GID>5609</GID>
<name>clock</name></connection>
<connection>
<GID>5605</GID>
<name>clock</name></connection>
<connection>
<GID>5583</GID>
<name>clock</name></connection>
<connection>
<GID>5573</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3915</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-752.5,229,-752.5</points>
<connection>
<GID>5631</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5627</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5623</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5619</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5615</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5611</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5607</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5589</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5578</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3916</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-737,66,-737</points>
<connection>
<GID>5639</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-737,60,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-721.5,60,-721.5</points>
<connection>
<GID>5637</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3917</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-737,89,-737</points>
<connection>
<GID>5643</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-737,83,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-721.5,83,-721.5</points>
<connection>
<GID>5641</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3918</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-737,114,-737</points>
<connection>
<GID>5647</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-737,108,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-721.5,108,-721.5</points>
<connection>
<GID>5645</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3919</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-737,137,-737</points>
<connection>
<GID>5651</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-737,131,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-721.5,131,-721.5</points>
<connection>
<GID>5649</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3920</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-737,160,-737</points>
<connection>
<GID>5655</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-737,154,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-721.5,154,-721.5</points>
<connection>
<GID>5653</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3921</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-737,183,-737</points>
<connection>
<GID>5659</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-737,177,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-721.5,177,-721.5</points>
<connection>
<GID>5657</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3922</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-737,208,-737</points>
<connection>
<GID>5663</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-737,202,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-721.5,202,-721.5</points>
<connection>
<GID>5661</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3923</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-737,231,-737</points>
<connection>
<GID>5667</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-737,225,-721.5</points>
<intersection>-737 1</intersection>
<intersection>-721.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-721.5,225,-721.5</points>
<connection>
<GID>5665</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3924</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-724.5,218,-724.5</points>
<connection>
<GID>5665</GID>
<name>clock</name></connection>
<connection>
<GID>5661</GID>
<name>clock</name></connection>
<connection>
<GID>5657</GID>
<name>clock</name></connection>
<connection>
<GID>5653</GID>
<name>clock</name></connection>
<connection>
<GID>5649</GID>
<name>clock</name></connection>
<connection>
<GID>5645</GID>
<name>clock</name></connection>
<connection>
<GID>5641</GID>
<name>clock</name></connection>
<connection>
<GID>5637</GID>
<name>clock</name></connection>
<connection>
<GID>5633</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3925</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-734,229,-734</points>
<connection>
<GID>5667</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5663</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5659</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5655</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5651</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5647</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5643</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5639</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5635</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3926</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-718,66,-718</points>
<connection>
<GID>5675</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-718,60,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-702.5,60,-702.5</points>
<connection>
<GID>5673</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3927</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-718,89,-718</points>
<connection>
<GID>5679</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-718,83,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-702.5,83,-702.5</points>
<connection>
<GID>5677</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-718,114,-718</points>
<connection>
<GID>5683</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-718,108,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-702.5,108,-702.5</points>
<connection>
<GID>5681</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3929</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-718,137,-718</points>
<connection>
<GID>5687</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-718,131,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-702.5,131,-702.5</points>
<connection>
<GID>5685</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3930</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-718,160,-718</points>
<connection>
<GID>5691</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-718,154,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-702.5,154,-702.5</points>
<connection>
<GID>5689</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3931</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-718,183,-718</points>
<connection>
<GID>5695</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-718,177,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-702.5,177,-702.5</points>
<connection>
<GID>5693</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3932</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-718,208,-718</points>
<connection>
<GID>5699</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-718,202,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-702.5,202,-702.5</points>
<connection>
<GID>5697</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3933</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-718,231,-718</points>
<connection>
<GID>5703</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-718,225,-702.5</points>
<intersection>-718 1</intersection>
<intersection>-702.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-702.5,225,-702.5</points>
<connection>
<GID>5701</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3934</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-705.5,218,-705.5</points>
<connection>
<GID>5701</GID>
<name>clock</name></connection>
<connection>
<GID>5697</GID>
<name>clock</name></connection>
<connection>
<GID>5693</GID>
<name>clock</name></connection>
<connection>
<GID>5689</GID>
<name>clock</name></connection>
<connection>
<GID>5685</GID>
<name>clock</name></connection>
<connection>
<GID>5681</GID>
<name>clock</name></connection>
<connection>
<GID>5677</GID>
<name>clock</name></connection>
<connection>
<GID>5673</GID>
<name>clock</name></connection>
<connection>
<GID>5669</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3935</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-715,229,-715</points>
<connection>
<GID>5703</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5699</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5695</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5691</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5687</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5683</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5679</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5675</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5671</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3936</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-699.5,66,-699.5</points>
<connection>
<GID>5711</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-699.5,60,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-684,60,-684</points>
<connection>
<GID>5709</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3937</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-699.5,89,-699.5</points>
<connection>
<GID>5715</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-699.5,83,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-684,83,-684</points>
<connection>
<GID>5713</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3938</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-699.5,114,-699.5</points>
<connection>
<GID>5719</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-699.5,108,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-684,108,-684</points>
<connection>
<GID>5717</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3939</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-699.5,137,-699.5</points>
<connection>
<GID>5723</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-699.5,131,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-684,131,-684</points>
<connection>
<GID>5721</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3940</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-699.5,160,-699.5</points>
<connection>
<GID>5727</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-699.5,154,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-684,154,-684</points>
<connection>
<GID>5725</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3941</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-699.5,183,-699.5</points>
<connection>
<GID>5731</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-699.5,177,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-684,177,-684</points>
<connection>
<GID>5729</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-699.5,208,-699.5</points>
<connection>
<GID>5735</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-699.5,202,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-684,202,-684</points>
<connection>
<GID>5733</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3943</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-699.5,231,-699.5</points>
<connection>
<GID>5739</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-699.5,225,-684</points>
<intersection>-699.5 1</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-684,225,-684</points>
<connection>
<GID>5737</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3944</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-687,218,-687</points>
<connection>
<GID>5737</GID>
<name>clock</name></connection>
<connection>
<GID>5733</GID>
<name>clock</name></connection>
<connection>
<GID>5729</GID>
<name>clock</name></connection>
<connection>
<GID>5725</GID>
<name>clock</name></connection>
<connection>
<GID>5721</GID>
<name>clock</name></connection>
<connection>
<GID>5717</GID>
<name>clock</name></connection>
<connection>
<GID>5713</GID>
<name>clock</name></connection>
<connection>
<GID>5709</GID>
<name>clock</name></connection>
<connection>
<GID>5705</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3945</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-696.5,229,-696.5</points>
<connection>
<GID>5739</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5735</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5731</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5727</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5723</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5719</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5715</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5711</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5707</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3946</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-833.5,66,-833.5</points>
<connection>
<GID>5747</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-833.5,60,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-818,60,-818</points>
<connection>
<GID>5745</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3947</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-833.5,89,-833.5</points>
<connection>
<GID>5751</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-833.5,83,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-818,83,-818</points>
<connection>
<GID>5749</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3948</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-833.5,114,-833.5</points>
<connection>
<GID>5755</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-833.5,108,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-818,108,-818</points>
<connection>
<GID>5753</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3949</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-833.5,137,-833.5</points>
<connection>
<GID>5396</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-833.5,131,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-818,131,-818</points>
<connection>
<GID>5394</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3950</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-833.5,160,-833.5</points>
<connection>
<GID>5400</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-833.5,154,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-818,154,-818</points>
<connection>
<GID>5398</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3951</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-833.5,183,-833.5</points>
<connection>
<GID>5404</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-833.5,177,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-818,177,-818</points>
<connection>
<GID>5402</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3952</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-833.5,208,-833.5</points>
<connection>
<GID>5408</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-833.5,202,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-818,202,-818</points>
<connection>
<GID>5406</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3953</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-833.5,231,-833.5</points>
<connection>
<GID>5412</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-833.5,225,-818</points>
<intersection>-833.5 1</intersection>
<intersection>-818 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-818,225,-818</points>
<connection>
<GID>5410</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-821,218,-821</points>
<connection>
<GID>5753</GID>
<name>clock</name></connection>
<connection>
<GID>5749</GID>
<name>clock</name></connection>
<connection>
<GID>5745</GID>
<name>clock</name></connection>
<connection>
<GID>5741</GID>
<name>OUT</name></connection>
<connection>
<GID>5410</GID>
<name>clock</name></connection>
<connection>
<GID>5406</GID>
<name>clock</name></connection>
<connection>
<GID>5402</GID>
<name>clock</name></connection>
<connection>
<GID>5398</GID>
<name>clock</name></connection>
<connection>
<GID>5394</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3955</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-830.5,229,-830.5</points>
<connection>
<GID>5755</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5751</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5747</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5743</GID>
<name>OUT</name></connection>
<connection>
<GID>5412</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5408</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5404</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5400</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5396</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3956</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-815,66,-815</points>
<connection>
<GID>5420</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-815,60,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-799.5,60,-799.5</points>
<connection>
<GID>5418</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3957</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-815,89,-815</points>
<connection>
<GID>5424</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-815,83,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-799.5,83,-799.5</points>
<connection>
<GID>5422</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3958</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-815,114,-815</points>
<connection>
<GID>5428</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-815,108,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-799.5,108,-799.5</points>
<connection>
<GID>5426</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-815,137,-815</points>
<connection>
<GID>5432</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-815,131,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-799.5,131,-799.5</points>
<connection>
<GID>5430</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3960</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-815,160,-815</points>
<connection>
<GID>5436</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-815,154,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-799.5,154,-799.5</points>
<connection>
<GID>5434</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3961</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-815,183,-815</points>
<connection>
<GID>5440</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-815,177,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-799.5,177,-799.5</points>
<connection>
<GID>5438</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3962</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-815,208,-815</points>
<connection>
<GID>5444</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-815,202,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-799.5,202,-799.5</points>
<connection>
<GID>5442</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3963</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-815,231,-815</points>
<connection>
<GID>5448</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-815,225,-799.5</points>
<intersection>-815 1</intersection>
<intersection>-799.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-799.5,225,-799.5</points>
<connection>
<GID>5446</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3964</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-802.5,218,-802.5</points>
<connection>
<GID>5446</GID>
<name>clock</name></connection>
<connection>
<GID>5442</GID>
<name>clock</name></connection>
<connection>
<GID>5438</GID>
<name>clock</name></connection>
<connection>
<GID>5434</GID>
<name>clock</name></connection>
<connection>
<GID>5430</GID>
<name>clock</name></connection>
<connection>
<GID>5426</GID>
<name>clock</name></connection>
<connection>
<GID>5422</GID>
<name>clock</name></connection>
<connection>
<GID>5418</GID>
<name>clock</name></connection>
<connection>
<GID>5414</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3965</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-812,229,-812</points>
<connection>
<GID>5448</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5444</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5440</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5436</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5432</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5428</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5424</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5420</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5416</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-796,66,-796</points>
<connection>
<GID>5458</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-796,60,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-780.5,60,-780.5</points>
<connection>
<GID>5456</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3967</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-796,89,-796</points>
<connection>
<GID>5463</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-796,83,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-780.5,83,-780.5</points>
<connection>
<GID>5461</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3968</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-796,114,-796</points>
<connection>
<GID>5468</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-796,108,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-780.5,108,-780.5</points>
<connection>
<GID>5466</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-796,137,-796</points>
<connection>
<GID>5473</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-796,131,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-780.5,131,-780.5</points>
<connection>
<GID>5471</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3970</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-796,160,-796</points>
<connection>
<GID>5478</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-796,154,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-780.5,154,-780.5</points>
<connection>
<GID>5476</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3971</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-796,183,-796</points>
<connection>
<GID>5481</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-796,177,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-780.5,177,-780.5</points>
<connection>
<GID>5480</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3972</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-796,208,-796</points>
<connection>
<GID>5484</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-796,202,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-780.5,202,-780.5</points>
<connection>
<GID>5483</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-796,231,-796</points>
<connection>
<GID>5486</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-796,225,-780.5</points>
<intersection>-796 1</intersection>
<intersection>-780.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-780.5,225,-780.5</points>
<connection>
<GID>5485</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-783.5,218,-783.5</points>
<connection>
<GID>5485</GID>
<name>clock</name></connection>
<connection>
<GID>5483</GID>
<name>clock</name></connection>
<connection>
<GID>5480</GID>
<name>clock</name></connection>
<connection>
<GID>5476</GID>
<name>clock</name></connection>
<connection>
<GID>5471</GID>
<name>clock</name></connection>
<connection>
<GID>5466</GID>
<name>clock</name></connection>
<connection>
<GID>5461</GID>
<name>clock</name></connection>
<connection>
<GID>5456</GID>
<name>clock</name></connection>
<connection>
<GID>5451</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3975</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-793,229,-793</points>
<connection>
<GID>5486</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5484</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5481</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5478</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5473</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5468</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5463</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5458</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5453</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3976</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-777.5,66,-777.5</points>
<connection>
<GID>5490</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-777.5,60,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-762,60,-762</points>
<connection>
<GID>5489</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>3977</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-777.5,89,-777.5</points>
<connection>
<GID>5492</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-777.5,83,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-762,83,-762</points>
<connection>
<GID>5491</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>3978</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-777.5,114,-777.5</points>
<connection>
<GID>5494</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-777.5,108,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-762,108,-762</points>
<connection>
<GID>5493</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>3979</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-777.5,137,-777.5</points>
<connection>
<GID>5496</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-777.5,131,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-762,131,-762</points>
<connection>
<GID>5495</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>3980</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-777.5,160,-777.5</points>
<connection>
<GID>5498</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-777.5,154,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-762,154,-762</points>
<connection>
<GID>5497</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>3981</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-777.5,183,-777.5</points>
<connection>
<GID>5500</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-777.5,177,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-762,177,-762</points>
<connection>
<GID>5499</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>3982</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-777.5,208,-777.5</points>
<connection>
<GID>5502</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-777.5,202,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-762,202,-762</points>
<connection>
<GID>5501</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>3983</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-777.5,231,-777.5</points>
<connection>
<GID>5504</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-777.5,225,-762</points>
<intersection>-777.5 1</intersection>
<intersection>-762 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-762,225,-762</points>
<connection>
<GID>5503</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>3984</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-765,218,-765</points>
<connection>
<GID>5503</GID>
<name>clock</name></connection>
<connection>
<GID>5501</GID>
<name>clock</name></connection>
<connection>
<GID>5499</GID>
<name>clock</name></connection>
<connection>
<GID>5497</GID>
<name>clock</name></connection>
<connection>
<GID>5495</GID>
<name>clock</name></connection>
<connection>
<GID>5493</GID>
<name>clock</name></connection>
<connection>
<GID>5491</GID>
<name>clock</name></connection>
<connection>
<GID>5489</GID>
<name>clock</name></connection>
<connection>
<GID>5487</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3985</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-774.5,229,-774.5</points>
<connection>
<GID>5504</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5502</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5500</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5498</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5496</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5494</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5492</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5490</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5488</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-843.5,47.5,-678.5</points>
<connection>
<GID>5520</GID>
<name>N_in1</name></connection>
<connection>
<GID>5505</GID>
<name>N_in0</name></connection>
<intersection>-818 12</intersection>
<intersection>-799.5 11</intersection>
<intersection>-780.5 10</intersection>
<intersection>-762 9</intersection>
<intersection>-740 8</intersection>
<intersection>-721.5 7</intersection>
<intersection>-702.5 6</intersection>
<intersection>-684 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-684,53,-684</points>
<connection>
<GID>5709</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>47.5,-702.5,53,-702.5</points>
<connection>
<GID>5673</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>47.5,-721.5,53,-721.5</points>
<connection>
<GID>5637</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>47.5,-740,53,-740</points>
<connection>
<GID>5583</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>47.5,-762,53,-762</points>
<connection>
<GID>5489</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>47.5,-780.5,53,-780.5</points>
<connection>
<GID>5456</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>47.5,-799.5,53,-799.5</points>
<connection>
<GID>5418</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>47.5,-818,53,-818</points>
<connection>
<GID>5745</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-843,70.5,-678</points>
<connection>
<GID>5521</GID>
<name>N_in1</name></connection>
<connection>
<GID>5506</GID>
<name>N_in0</name></connection>
<intersection>-826 4</intersection>
<intersection>-807.5 5</intersection>
<intersection>-788.5 6</intersection>
<intersection>-770 7</intersection>
<intersection>-748 8</intersection>
<intersection>-729.5 9</intersection>
<intersection>-710.5 10</intersection>
<intersection>-692 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>66,-826,70.5,-826</points>
<intersection>66 12</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66,-807.5,70.5,-807.5</points>
<intersection>66 13</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66,-788.5,70.5,-788.5</points>
<intersection>66 14</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66,-770,70.5,-770</points>
<intersection>66 15</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66,-748,70.5,-748</points>
<intersection>66 18</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66,-729.5,70.5,-729.5</points>
<intersection>66 19</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>66,-710.5,70.5,-710.5</points>
<intersection>66 20</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>66,-692,70.5,-692</points>
<intersection>66 21</intersection>
<intersection>70.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>66,-828,66,-826</points>
<connection>
<GID>5747</GID>
<name>OUT_0</name></connection>
<intersection>-826 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>66,-809.5,66,-807.5</points>
<connection>
<GID>5420</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>66,-790.5,66,-788.5</points>
<connection>
<GID>5458</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>66,-772,66,-770</points>
<connection>
<GID>5490</GID>
<name>OUT_0</name></connection>
<intersection>-770 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>66,-750,66,-748</points>
<connection>
<GID>5589</GID>
<name>OUT_0</name></connection>
<intersection>-748 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>66,-731.5,66,-729.5</points>
<connection>
<GID>5639</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>66,-712.5,66,-710.5</points>
<connection>
<GID>5675</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>66,-694,66,-692</points>
<connection>
<GID>5711</GID>
<name>OUT_0</name></connection>
<intersection>-692 11</intersection></vsegment></shape></wire>
<wire>
<ID>3988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-843,73.5,-678.5</points>
<connection>
<GID>5522</GID>
<name>N_in1</name></connection>
<connection>
<GID>5507</GID>
<name>N_in0</name></connection>
<intersection>-818 10</intersection>
<intersection>-799.5 9</intersection>
<intersection>-780.5 8</intersection>
<intersection>-762 7</intersection>
<intersection>-740 6</intersection>
<intersection>-721.5 5</intersection>
<intersection>-702.5 4</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73.5,-684,76,-684</points>
<connection>
<GID>5713</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-702.5,76,-702.5</points>
<connection>
<GID>5677</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>73.5,-721.5,76,-721.5</points>
<connection>
<GID>5641</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>73.5,-740,76,-740</points>
<connection>
<GID>5605</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>73.5,-762,76,-762</points>
<connection>
<GID>5491</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>73.5,-780.5,76,-780.5</points>
<connection>
<GID>5461</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>73.5,-799.5,76,-799.5</points>
<connection>
<GID>5422</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>73.5,-818,76,-818</points>
<connection>
<GID>5749</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-843,93,-678</points>
<connection>
<GID>5523</GID>
<name>N_in1</name></connection>
<connection>
<GID>5508</GID>
<name>N_in0</name></connection>
<intersection>-826 6</intersection>
<intersection>-807.5 7</intersection>
<intersection>-788.5 8</intersection>
<intersection>-770 9</intersection>
<intersection>-748 10</intersection>
<intersection>-729.5 11</intersection>
<intersection>-710.5 12</intersection>
<intersection>-692 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89,-826,93,-826</points>
<intersection>89 14</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89,-807.5,93,-807.5</points>
<intersection>89 15</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89,-788.5,93,-788.5</points>
<intersection>89 16</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89,-770,93,-770</points>
<intersection>89 17</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>89,-748,93,-748</points>
<intersection>89 20</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89,-729.5,93,-729.5</points>
<intersection>89 21</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>89,-710.5,93,-710.5</points>
<intersection>89 22</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>89,-692,93,-692</points>
<intersection>89 23</intersection>
<intersection>93 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>89,-828,89,-826</points>
<connection>
<GID>5751</GID>
<name>OUT_0</name></connection>
<intersection>-826 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>89,-809.5,89,-807.5</points>
<connection>
<GID>5424</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>89,-790.5,89,-788.5</points>
<connection>
<GID>5463</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>89,-772,89,-770</points>
<connection>
<GID>5492</GID>
<name>OUT_0</name></connection>
<intersection>-770 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>89,-750,89,-748</points>
<connection>
<GID>5607</GID>
<name>OUT_0</name></connection>
<intersection>-748 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>89,-731.5,89,-729.5</points>
<connection>
<GID>5643</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>89,-712.5,89,-710.5</points>
<connection>
<GID>5679</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>89,-694,89,-692</points>
<connection>
<GID>5715</GID>
<name>OUT_0</name></connection>
<intersection>-692 13</intersection></vsegment></shape></wire>
<wire>
<ID>3990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-843,96.5,-678</points>
<connection>
<GID>5524</GID>
<name>N_in1</name></connection>
<connection>
<GID>5509</GID>
<name>N_in0</name></connection>
<intersection>-818 13</intersection>
<intersection>-799.5 12</intersection>
<intersection>-780.5 11</intersection>
<intersection>-762 10</intersection>
<intersection>-740 9</intersection>
<intersection>-721.5 8</intersection>
<intersection>-702.5 7</intersection>
<intersection>-684 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>96.5,-684,101,-684</points>
<connection>
<GID>5717</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>96.5,-702.5,101,-702.5</points>
<connection>
<GID>5681</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>96.5,-721.5,101,-721.5</points>
<connection>
<GID>5645</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>96.5,-740,101,-740</points>
<connection>
<GID>5609</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>96.5,-762,101,-762</points>
<connection>
<GID>5493</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>96.5,-780.5,101,-780.5</points>
<connection>
<GID>5466</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>96.5,-799.5,101,-799.5</points>
<connection>
<GID>5426</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>96.5,-818,101,-818</points>
<connection>
<GID>5753</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-843,117.5,-678.5</points>
<connection>
<GID>5525</GID>
<name>N_in1</name></connection>
<connection>
<GID>5510</GID>
<name>N_in0</name></connection>
<intersection>-826 6</intersection>
<intersection>-807.5 7</intersection>
<intersection>-788.5 8</intersection>
<intersection>-770 9</intersection>
<intersection>-748 10</intersection>
<intersection>-729.5 11</intersection>
<intersection>-710.5 12</intersection>
<intersection>-692 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>114,-826,117.5,-826</points>
<intersection>114 14</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114,-807.5,117.5,-807.5</points>
<intersection>114 15</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114,-788.5,117.5,-788.5</points>
<intersection>114 16</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114,-770,117.5,-770</points>
<intersection>114 17</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114,-748,117.5,-748</points>
<intersection>114 20</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>114,-729.5,117.5,-729.5</points>
<intersection>114 21</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114,-710.5,117.5,-710.5</points>
<intersection>114 22</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>114,-692,117.5,-692</points>
<intersection>114 23</intersection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>114,-828,114,-826</points>
<connection>
<GID>5755</GID>
<name>OUT_0</name></connection>
<intersection>-826 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>114,-809.5,114,-807.5</points>
<connection>
<GID>5428</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>114,-790.5,114,-788.5</points>
<connection>
<GID>5468</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>114,-772,114,-770</points>
<connection>
<GID>5494</GID>
<name>OUT_0</name></connection>
<intersection>-770 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>114,-750,114,-748</points>
<connection>
<GID>5611</GID>
<name>OUT_0</name></connection>
<intersection>-748 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>114,-731.5,114,-729.5</points>
<connection>
<GID>5647</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>114,-712.5,114,-710.5</points>
<connection>
<GID>5683</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>114,-694,114,-692</points>
<connection>
<GID>5719</GID>
<name>OUT_0</name></connection>
<intersection>-692 13</intersection></vsegment></shape></wire>
<wire>
<ID>3992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-843,121.5,-678</points>
<connection>
<GID>5526</GID>
<name>N_in1</name></connection>
<connection>
<GID>5511</GID>
<name>N_in0</name></connection>
<intersection>-818 13</intersection>
<intersection>-799.5 12</intersection>
<intersection>-780.5 11</intersection>
<intersection>-762 10</intersection>
<intersection>-740 9</intersection>
<intersection>-721.5 8</intersection>
<intersection>-702.5 7</intersection>
<intersection>-684 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>121.5,-684,124,-684</points>
<connection>
<GID>5721</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>121.5,-702.5,124,-702.5</points>
<connection>
<GID>5685</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121.5,-721.5,124,-721.5</points>
<connection>
<GID>5649</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>121.5,-740,124,-740</points>
<connection>
<GID>5613</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>121.5,-762,124,-762</points>
<connection>
<GID>5495</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>121.5,-780.5,124,-780.5</points>
<connection>
<GID>5471</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>121.5,-799.5,124,-799.5</points>
<connection>
<GID>5430</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>121.5,-818,124,-818</points>
<connection>
<GID>5394</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3993</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-843,140,-678</points>
<connection>
<GID>5527</GID>
<name>N_in1</name></connection>
<connection>
<GID>5512</GID>
<name>N_in0</name></connection>
<intersection>-826 6</intersection>
<intersection>-807.5 7</intersection>
<intersection>-788.5 8</intersection>
<intersection>-770 9</intersection>
<intersection>-748 10</intersection>
<intersection>-729.5 11</intersection>
<intersection>-710.5 12</intersection>
<intersection>-692 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>137,-826,140,-826</points>
<intersection>137 14</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137,-807.5,140,-807.5</points>
<intersection>137 15</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-788.5,140,-788.5</points>
<intersection>137 16</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137,-770,140,-770</points>
<intersection>137 17</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-748,140,-748</points>
<intersection>137 20</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>137,-729.5,140,-729.5</points>
<intersection>137 21</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137,-710.5,140,-710.5</points>
<intersection>137 22</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-692,140,-692</points>
<intersection>137 23</intersection>
<intersection>140 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>137,-828,137,-826</points>
<connection>
<GID>5396</GID>
<name>OUT_0</name></connection>
<intersection>-826 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>137,-809.5,137,-807.5</points>
<connection>
<GID>5432</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>137,-790.5,137,-788.5</points>
<connection>
<GID>5473</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>137,-772,137,-770</points>
<connection>
<GID>5496</GID>
<name>OUT_0</name></connection>
<intersection>-770 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>137,-750,137,-748</points>
<connection>
<GID>5615</GID>
<name>OUT_0</name></connection>
<intersection>-748 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>137,-731.5,137,-729.5</points>
<connection>
<GID>5651</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>137,-712.5,137,-710.5</points>
<connection>
<GID>5687</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>137,-694,137,-692</points>
<connection>
<GID>5723</GID>
<name>OUT_0</name></connection>
<intersection>-692 13</intersection></vsegment></shape></wire>
<wire>
<ID>3994</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-843,144,-678</points>
<connection>
<GID>5528</GID>
<name>N_in1</name></connection>
<connection>
<GID>5513</GID>
<name>N_in0</name></connection>
<intersection>-818 13</intersection>
<intersection>-799.5 12</intersection>
<intersection>-780.5 11</intersection>
<intersection>-762 10</intersection>
<intersection>-740 9</intersection>
<intersection>-721.5 8</intersection>
<intersection>-702.5 7</intersection>
<intersection>-684 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>144,-684,147,-684</points>
<connection>
<GID>5725</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>144,-702.5,147,-702.5</points>
<connection>
<GID>5689</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>144,-721.5,147,-721.5</points>
<connection>
<GID>5653</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>144,-740,147,-740</points>
<connection>
<GID>5617</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>144,-762,147,-762</points>
<connection>
<GID>5497</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>144,-780.5,147,-780.5</points>
<connection>
<GID>5476</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>144,-799.5,147,-799.5</points>
<connection>
<GID>5434</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>144,-818,147,-818</points>
<connection>
<GID>5398</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>3995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-842.5,163,-678</points>
<connection>
<GID>5529</GID>
<name>N_in1</name></connection>
<connection>
<GID>5514</GID>
<name>N_in0</name></connection>
<intersection>-826 6</intersection>
<intersection>-807.5 7</intersection>
<intersection>-788.5 8</intersection>
<intersection>-770 9</intersection>
<intersection>-748 10</intersection>
<intersection>-729.5 11</intersection>
<intersection>-710.5 12</intersection>
<intersection>-692 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>160,-826,163,-826</points>
<intersection>160 14</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>160,-807.5,163,-807.5</points>
<intersection>160 15</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>160,-788.5,163,-788.5</points>
<intersection>160 16</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>160,-770,163,-770</points>
<intersection>160 17</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>160,-748,163,-748</points>
<intersection>160 20</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>160,-729.5,163,-729.5</points>
<intersection>160 21</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>160,-710.5,163,-710.5</points>
<intersection>160 22</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>160,-692,163,-692</points>
<intersection>160 23</intersection>
<intersection>163 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>160,-828,160,-826</points>
<connection>
<GID>5400</GID>
<name>OUT_0</name></connection>
<intersection>-826 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>160,-809.5,160,-807.5</points>
<connection>
<GID>5436</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>160,-790.5,160,-788.5</points>
<connection>
<GID>5478</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>160,-772,160,-770</points>
<connection>
<GID>5498</GID>
<name>OUT_0</name></connection>
<intersection>-770 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>160,-750,160,-748</points>
<connection>
<GID>5619</GID>
<name>OUT_0</name></connection>
<intersection>-748 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>160,-731.5,160,-729.5</points>
<connection>
<GID>5655</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>160,-712.5,160,-710.5</points>
<connection>
<GID>5691</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>160,-694,160,-692</points>
<connection>
<GID>5727</GID>
<name>OUT_0</name></connection>
<intersection>-692 13</intersection></vsegment></shape></wire>
<wire>
<ID>3996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-842.5,168,-678</points>
<connection>
<GID>5530</GID>
<name>N_in1</name></connection>
<connection>
<GID>5515</GID>
<name>N_in0</name></connection>
<intersection>-818 13</intersection>
<intersection>-799.5 12</intersection>
<intersection>-780.5 11</intersection>
<intersection>-762 10</intersection>
<intersection>-740 9</intersection>
<intersection>-721.5 8</intersection>
<intersection>-702.5 7</intersection>
<intersection>-684 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>168,-684,170,-684</points>
<connection>
<GID>5729</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>168,-702.5,170,-702.5</points>
<connection>
<GID>5693</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>168,-721.5,170,-721.5</points>
<connection>
<GID>5657</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>168,-740,170,-740</points>
<connection>
<GID>5621</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>168,-762,170,-762</points>
<connection>
<GID>5499</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>168,-780.5,170,-780.5</points>
<connection>
<GID>5480</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>168,-799.5,170,-799.5</points>
<connection>
<GID>5438</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>168,-818,170,-818</points>
<connection>
<GID>5402</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>3997</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-842,186,-678</points>
<connection>
<GID>5531</GID>
<name>N_in1</name></connection>
<connection>
<GID>5517</GID>
<name>N_in0</name></connection>
<intersection>-826 16</intersection>
<intersection>-807.5 15</intersection>
<intersection>-788.5 14</intersection>
<intersection>-770 13</intersection>
<intersection>-748 12</intersection>
<intersection>-729.5 11</intersection>
<intersection>-710.5 10</intersection>
<intersection>-692 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>183,-692,186,-692</points>
<intersection>183 26</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183,-710.5,186,-710.5</points>
<intersection>183 25</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183,-729.5,186,-729.5</points>
<intersection>183 24</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183,-748,186,-748</points>
<intersection>183 23</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183,-770,186,-770</points>
<intersection>183 20</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>183,-788.5,186,-788.5</points>
<intersection>183 19</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>183,-807.5,186,-807.5</points>
<intersection>183 18</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>183,-826,186,-826</points>
<intersection>183 17</intersection>
<intersection>186 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>183,-828,183,-826</points>
<connection>
<GID>5404</GID>
<name>OUT_0</name></connection>
<intersection>-826 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>183,-809.5,183,-807.5</points>
<connection>
<GID>5440</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>183,-790.5,183,-788.5</points>
<connection>
<GID>5481</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>183,-772,183,-770</points>
<connection>
<GID>5500</GID>
<name>OUT_0</name></connection>
<intersection>-770 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>183,-750,183,-748</points>
<connection>
<GID>5623</GID>
<name>OUT_0</name></connection>
<intersection>-748 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>183,-731.5,183,-729.5</points>
<connection>
<GID>5659</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>183,-712.5,183,-710.5</points>
<connection>
<GID>5695</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>183,-694,183,-692</points>
<connection>
<GID>5731</GID>
<name>OUT_0</name></connection>
<intersection>-692 9</intersection></vsegment></shape></wire>
<wire>
<ID>3998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-842,190.5,-678</points>
<connection>
<GID>5532</GID>
<name>N_in1</name></connection>
<connection>
<GID>5516</GID>
<name>N_in0</name></connection>
<intersection>-818 13</intersection>
<intersection>-799.5 12</intersection>
<intersection>-780.5 11</intersection>
<intersection>-762 10</intersection>
<intersection>-740 9</intersection>
<intersection>-721.5 8</intersection>
<intersection>-702.5 7</intersection>
<intersection>-684 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>190.5,-684,195,-684</points>
<connection>
<GID>5733</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>190.5,-702.5,195,-702.5</points>
<connection>
<GID>5697</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>190.5,-721.5,195,-721.5</points>
<connection>
<GID>5661</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>190.5,-740,195,-740</points>
<connection>
<GID>5625</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>190.5,-762,195,-762</points>
<connection>
<GID>5501</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>190.5,-780.5,195,-780.5</points>
<connection>
<GID>5483</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>190.5,-799.5,195,-799.5</points>
<connection>
<GID>5442</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>190.5,-818,195,-818</points>
<connection>
<GID>5406</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,-841.5,211.5,-678.5</points>
<connection>
<GID>5533</GID>
<name>N_in1</name></connection>
<connection>
<GID>5518</GID>
<name>N_in0</name></connection>
<intersection>-826 6</intersection>
<intersection>-807.5 7</intersection>
<intersection>-788.5 8</intersection>
<intersection>-770 9</intersection>
<intersection>-748 10</intersection>
<intersection>-729.5 11</intersection>
<intersection>-710.5 12</intersection>
<intersection>-692 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>208,-826,211.5,-826</points>
<intersection>208 14</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>208,-807.5,211.5,-807.5</points>
<intersection>208 15</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>208,-788.5,211.5,-788.5</points>
<intersection>208 16</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>208,-770,211.5,-770</points>
<intersection>208 17</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>208,-748,211.5,-748</points>
<intersection>208 20</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>208,-729.5,211.5,-729.5</points>
<intersection>208 21</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>208,-710.5,211.5,-710.5</points>
<intersection>208 22</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>208,-692,211.5,-692</points>
<intersection>208 23</intersection>
<intersection>211.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>208,-828,208,-826</points>
<connection>
<GID>5408</GID>
<name>OUT_0</name></connection>
<intersection>-826 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>208,-809.5,208,-807.5</points>
<connection>
<GID>5444</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>208,-790.5,208,-788.5</points>
<connection>
<GID>5484</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>208,-772,208,-770</points>
<connection>
<GID>5502</GID>
<name>OUT_0</name></connection>
<intersection>-770 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>208,-750,208,-748</points>
<connection>
<GID>5627</GID>
<name>OUT_0</name></connection>
<intersection>-748 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>208,-731.5,208,-729.5</points>
<connection>
<GID>5663</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>208,-712.5,208,-710.5</points>
<connection>
<GID>5699</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>208,-694,208,-692</points>
<connection>
<GID>5735</GID>
<name>OUT_0</name></connection>
<intersection>-692 13</intersection></vsegment></shape></wire>
<wire>
<ID>4000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215,-841.5,215,-678.5</points>
<connection>
<GID>5534</GID>
<name>N_in1</name></connection>
<connection>
<GID>5535</GID>
<name>N_in0</name></connection>
<intersection>-818 11</intersection>
<intersection>-799.5 10</intersection>
<intersection>-780.5 9</intersection>
<intersection>-762 7</intersection>
<intersection>-740 6</intersection>
<intersection>-721.5 5</intersection>
<intersection>-702.5 4</intersection>
<intersection>-684 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-684,218,-684</points>
<connection>
<GID>5737</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>215,-702.5,218,-702.5</points>
<connection>
<GID>5701</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>215,-721.5,218,-721.5</points>
<connection>
<GID>5665</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>215,-740,218,-740</points>
<connection>
<GID>5629</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>215,-762,218,-762</points>
<connection>
<GID>5503</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>215,-780.5,218,-780.5</points>
<connection>
<GID>5485</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>215,-799.5,218,-799.5</points>
<connection>
<GID>5446</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>215,-818,218,-818</points>
<connection>
<GID>5410</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment></shape></wire>
<wire>
<ID>4001</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-841.5,236,-679.5</points>
<connection>
<GID>5536</GID>
<name>N_in1</name></connection>
<connection>
<GID>5519</GID>
<name>N_in0</name></connection>
<intersection>-826 11</intersection>
<intersection>-807.5 10</intersection>
<intersection>-788.5 9</intersection>
<intersection>-770 8</intersection>
<intersection>-748 7</intersection>
<intersection>-729.5 6</intersection>
<intersection>-710.5 5</intersection>
<intersection>-692 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>231,-692,236,-692</points>
<intersection>231 21</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>231,-710.5,236,-710.5</points>
<intersection>231 20</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>231,-729.5,236,-729.5</points>
<intersection>231 19</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>231,-748,236,-748</points>
<intersection>231 18</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>231,-770,236,-770</points>
<intersection>231 15</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>231,-788.5,236,-788.5</points>
<intersection>231 14</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>231,-807.5,236,-807.5</points>
<intersection>231 13</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>231,-826,236,-826</points>
<intersection>231 12</intersection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>231,-828,231,-826</points>
<connection>
<GID>5412</GID>
<name>OUT_0</name></connection>
<intersection>-826 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>231,-809.5,231,-807.5</points>
<connection>
<GID>5448</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>231,-790.5,231,-788.5</points>
<connection>
<GID>5486</GID>
<name>OUT_0</name></connection>
<intersection>-788.5 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>231,-772,231,-770</points>
<connection>
<GID>5504</GID>
<name>OUT_0</name></connection>
<intersection>-770 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>231,-750,231,-748</points>
<connection>
<GID>5631</GID>
<name>OUT_0</name></connection>
<intersection>-748 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>231,-731.5,231,-729.5</points>
<connection>
<GID>5667</GID>
<name>OUT_0</name></connection>
<intersection>-729.5 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>231,-712.5,231,-710.5</points>
<connection>
<GID>5703</GID>
<name>OUT_0</name></connection>
<intersection>-710.5 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>231,-694,231,-692</points>
<connection>
<GID>5739</GID>
<name>OUT_0</name></connection>
<intersection>-692 4</intersection></vsegment></shape></wire>
<wire>
<ID>4002</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-121,-686,25.5,-686</points>
<connection>
<GID>5705</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-837.5,-121,-686</points>
<connection>
<GID>5542</GID>
<name>OUT_15</name></connection>
<intersection>-695.5 4</intersection>
<intersection>-686 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-695.5,37,-695.5</points>
<connection>
<GID>5707</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4003</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-120,-704.5,25.5,-704.5</points>
<connection>
<GID>5669</GID>
<name>IN_0</name></connection>
<intersection>-120 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-120,-838.5,-120,-704.5</points>
<intersection>-838.5 6</intersection>
<intersection>-714 5</intersection>
<intersection>-704.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-120,-714,37,-714</points>
<connection>
<GID>5671</GID>
<name>IN_0</name></connection>
<intersection>-120 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-121,-838.5,-120,-838.5</points>
<connection>
<GID>5542</GID>
<name>OUT_14</name></connection>
<intersection>-120 4</intersection></hsegment></shape></wire>
<wire>
<ID>4004</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-119,-723.5,25.5,-723.5</points>
<connection>
<GID>5633</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-839.5,-119,-723.5</points>
<intersection>-839.5 6</intersection>
<intersection>-733 4</intersection>
<intersection>-723.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-733,37,-733</points>
<connection>
<GID>5635</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-121,-839.5,-119,-839.5</points>
<connection>
<GID>5542</GID>
<name>OUT_13</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>4005</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-118,-742,25.5,-742</points>
<connection>
<GID>5573</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118,-840.5,-118,-742</points>
<intersection>-840.5 5</intersection>
<intersection>-751.5 4</intersection>
<intersection>-742 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118,-751.5,37,-751.5</points>
<connection>
<GID>5578</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-840.5,-118,-840.5</points>
<connection>
<GID>5542</GID>
<name>OUT_12</name></connection>
<intersection>-118 3</intersection></hsegment></shape></wire>
<wire>
<ID>4006</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-117,-764,25.5,-764</points>
<connection>
<GID>5487</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-841.5,-117,-764</points>
<intersection>-841.5 6</intersection>
<intersection>-773.5 4</intersection>
<intersection>-764 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-773.5,36.5,-773.5</points>
<connection>
<GID>5488</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-121,-841.5,-117,-841.5</points>
<connection>
<GID>5542</GID>
<name>OUT_11</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>4007</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,-782.5,25.5,-782.5</points>
<connection>
<GID>5451</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-116,-842.5,-116,-782.5</points>
<intersection>-842.5 5</intersection>
<intersection>-792 4</intersection>
<intersection>-782.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-116,-792,36.5,-792</points>
<connection>
<GID>5453</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-842.5,-116,-842.5</points>
<connection>
<GID>5542</GID>
<name>OUT_10</name></connection>
<intersection>-116 3</intersection></hsegment></shape></wire>
<wire>
<ID>4008</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115,-801.5,25.5,-801.5</points>
<connection>
<GID>5414</GID>
<name>IN_0</name></connection>
<intersection>-115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-115,-843.5,-115,-801.5</points>
<intersection>-843.5 5</intersection>
<intersection>-811 4</intersection>
<intersection>-801.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-115,-811,36.5,-811</points>
<connection>
<GID>5416</GID>
<name>IN_0</name></connection>
<intersection>-115 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-843.5,-115,-843.5</points>
<connection>
<GID>5542</GID>
<name>OUT_9</name></connection>
<intersection>-115 3</intersection></hsegment></shape></wire>
<wire>
<ID>4009</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-820,25.5,-820</points>
<connection>
<GID>5741</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114,-844.5,-114,-820</points>
<intersection>-844.5 5</intersection>
<intersection>-829.5 4</intersection>
<intersection>-820 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-114,-829.5,36.5,-829.5</points>
<connection>
<GID>5743</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-844.5,-114,-844.5</points>
<connection>
<GID>5542</GID>
<name>OUT_8</name></connection>
<intersection>-114 3</intersection></hsegment></shape></wire>
<wire>
<ID>4010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-843.5,24.5,-678.5</points>
<connection>
<GID>5540</GID>
<name>N_in1</name></connection>
<connection>
<GID>5538</GID>
<name>N_in0</name></connection>
<intersection>-822 10</intersection>
<intersection>-803.5 9</intersection>
<intersection>-784.5 8</intersection>
<intersection>-766 7</intersection>
<intersection>-744 6</intersection>
<intersection>-725.5 5</intersection>
<intersection>-706.5 4</intersection>
<intersection>-688 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-688,25.5,-688</points>
<connection>
<GID>5705</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-706.5,25.5,-706.5</points>
<connection>
<GID>5669</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>24.5,-725.5,25.5,-725.5</points>
<connection>
<GID>5633</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>24.5,-744,25.5,-744</points>
<connection>
<GID>5573</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>24.5,-766,25.5,-766</points>
<connection>
<GID>5487</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>24.5,-784.5,25.5,-784.5</points>
<connection>
<GID>5451</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>24.5,-803.5,25.5,-803.5</points>
<connection>
<GID>5414</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>24.5,-822,25.5,-822</points>
<connection>
<GID>5741</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-843.5,34.5,-678.5</points>
<connection>
<GID>5539</GID>
<name>N_in1</name></connection>
<connection>
<GID>5537</GID>
<name>N_in0</name></connection>
<intersection>-831.5 3</intersection>
<intersection>-813 5</intersection>
<intersection>-794 7</intersection>
<intersection>-775.5 9</intersection>
<intersection>-753.5 11</intersection>
<intersection>-735 13</intersection>
<intersection>-716 15</intersection>
<intersection>-697.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34.5,-831.5,36.5,-831.5</points>
<connection>
<GID>5743</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>34.5,-813,36.5,-813</points>
<connection>
<GID>5416</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>34.5,-794,36.5,-794</points>
<connection>
<GID>5453</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>34.5,-775.5,36.5,-775.5</points>
<connection>
<GID>5488</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>34.5,-753.5,37,-753.5</points>
<connection>
<GID>5578</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>34.5,-735,37,-735</points>
<connection>
<GID>5635</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>34.5,-716,37,-716</points>
<connection>
<GID>5671</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>34.5,-697.5,37,-697.5</points>
<connection>
<GID>5707</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4012</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-931,66,-931</points>
<connection>
<GID>5638</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-931,60,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-915.5,60,-915.5</points>
<connection>
<GID>5626</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4013</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-931,89,-931</points>
<connection>
<GID>5664</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-931,83,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-915.5,83,-915.5</points>
<connection>
<GID>5662</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4014</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-931,114,-931</points>
<connection>
<GID>5672</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-931,108,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-915.5,108,-915.5</points>
<connection>
<GID>5668</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4015</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-931,137,-931</points>
<connection>
<GID>5680</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-931,131,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-915.5,131,-915.5</points>
<connection>
<GID>5676</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4016</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-931,160,-931</points>
<connection>
<GID>5686</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-931,154,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-915.5,154,-915.5</points>
<connection>
<GID>5682</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4017</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-931,183,-931</points>
<connection>
<GID>5690</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-931,177,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-915.5,177,-915.5</points>
<connection>
<GID>5688</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4018</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-931,208,-931</points>
<connection>
<GID>5694</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-931,202,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-915.5,202,-915.5</points>
<connection>
<GID>5692</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4019</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-931,231,-931</points>
<connection>
<GID>5698</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-931,225,-915.5</points>
<intersection>-931 1</intersection>
<intersection>-915.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-915.5,225,-915.5</points>
<connection>
<GID>5696</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4020</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-918.5,218,-918.5</points>
<connection>
<GID>5696</GID>
<name>clock</name></connection>
<connection>
<GID>5692</GID>
<name>clock</name></connection>
<connection>
<GID>5688</GID>
<name>clock</name></connection>
<connection>
<GID>5682</GID>
<name>clock</name></connection>
<connection>
<GID>5676</GID>
<name>clock</name></connection>
<connection>
<GID>5668</GID>
<name>clock</name></connection>
<connection>
<GID>5662</GID>
<name>clock</name></connection>
<connection>
<GID>5626</GID>
<name>clock</name></connection>
<connection>
<GID>5620</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4021</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-928,229,-928</points>
<connection>
<GID>5698</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5694</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5690</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5686</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5672</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5664</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5638</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5622</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4022</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-912.5,66,-912.5</points>
<connection>
<GID>5706</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-912.5,60,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-897,60,-897</points>
<connection>
<GID>5704</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4023</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-912.5,89,-912.5</points>
<connection>
<GID>5710</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-912.5,83,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-897,83,-897</points>
<connection>
<GID>5708</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4024</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-912.5,114,-912.5</points>
<connection>
<GID>5714</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-912.5,108,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-897,108,-897</points>
<connection>
<GID>5712</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4025</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-912.5,137,-912.5</points>
<connection>
<GID>5718</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-912.5,131,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-897,131,-897</points>
<connection>
<GID>5716</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4026</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-912.5,160,-912.5</points>
<connection>
<GID>5722</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-912.5,154,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-897,154,-897</points>
<connection>
<GID>5720</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4027</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-912.5,183,-912.5</points>
<connection>
<GID>5726</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-912.5,177,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-897,177,-897</points>
<connection>
<GID>5724</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4028</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-912.5,208,-912.5</points>
<connection>
<GID>5730</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-912.5,202,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-897,202,-897</points>
<connection>
<GID>5728</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4029</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-912.5,231,-912.5</points>
<connection>
<GID>5734</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-912.5,225,-897</points>
<intersection>-912.5 1</intersection>
<intersection>-897 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-897,225,-897</points>
<connection>
<GID>5732</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4030</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-900,218,-900</points>
<connection>
<GID>5732</GID>
<name>clock</name></connection>
<connection>
<GID>5728</GID>
<name>clock</name></connection>
<connection>
<GID>5724</GID>
<name>clock</name></connection>
<connection>
<GID>5720</GID>
<name>clock</name></connection>
<connection>
<GID>5716</GID>
<name>clock</name></connection>
<connection>
<GID>5712</GID>
<name>clock</name></connection>
<connection>
<GID>5708</GID>
<name>clock</name></connection>
<connection>
<GID>5704</GID>
<name>clock</name></connection>
<connection>
<GID>5700</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4031</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-909.5,229,-909.5</points>
<connection>
<GID>5734</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5730</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5726</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5722</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5718</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5714</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5710</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5706</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5702</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4032</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-893.5,66,-893.5</points>
<connection>
<GID>5742</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-893.5,60,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-878,60,-878</points>
<connection>
<GID>5740</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-893.5,89,-893.5</points>
<connection>
<GID>5746</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-893.5,83,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-878,83,-878</points>
<connection>
<GID>5744</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4034</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-893.5,114,-893.5</points>
<connection>
<GID>5750</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-893.5,108,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-878,108,-878</points>
<connection>
<GID>5748</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4035</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-893.5,137,-893.5</points>
<connection>
<GID>5754</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-893.5,131,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-878,131,-878</points>
<connection>
<GID>5752</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-893.5,160,-893.5</points>
<connection>
<GID>5395</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-893.5,154,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-878,154,-878</points>
<connection>
<GID>5756</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-893.5,183,-893.5</points>
<connection>
<GID>5399</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-893.5,177,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-878,177,-878</points>
<connection>
<GID>5397</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4038</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-893.5,208,-893.5</points>
<connection>
<GID>5403</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-893.5,202,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-878,202,-878</points>
<connection>
<GID>5401</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4039</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-893.5,231,-893.5</points>
<connection>
<GID>5407</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-893.5,225,-878</points>
<intersection>-893.5 1</intersection>
<intersection>-878 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-878,225,-878</points>
<connection>
<GID>5405</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4040</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-881,218,-881</points>
<connection>
<GID>5756</GID>
<name>clock</name></connection>
<connection>
<GID>5752</GID>
<name>clock</name></connection>
<connection>
<GID>5748</GID>
<name>clock</name></connection>
<connection>
<GID>5744</GID>
<name>clock</name></connection>
<connection>
<GID>5740</GID>
<name>clock</name></connection>
<connection>
<GID>5736</GID>
<name>OUT</name></connection>
<connection>
<GID>5405</GID>
<name>clock</name></connection>
<connection>
<GID>5401</GID>
<name>clock</name></connection>
<connection>
<GID>5397</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-890.5,229,-890.5</points>
<connection>
<GID>5754</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5746</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5742</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5738</GID>
<name>OUT</name></connection>
<connection>
<GID>5407</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5403</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5399</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5395</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4042</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-875,66,-875</points>
<connection>
<GID>5415</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-875,60,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-859.5,60,-859.5</points>
<connection>
<GID>5413</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4043</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-875,89,-875</points>
<connection>
<GID>5419</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-875,83,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-859.5,83,-859.5</points>
<connection>
<GID>5417</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4044</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-875,114,-875</points>
<connection>
<GID>5423</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-875,108,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-859.5,108,-859.5</points>
<connection>
<GID>5421</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-875,137,-875</points>
<connection>
<GID>5427</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-875,131,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-859.5,131,-859.5</points>
<connection>
<GID>5425</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4046</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-875,160,-875</points>
<connection>
<GID>5431</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-875,154,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-859.5,154,-859.5</points>
<connection>
<GID>5429</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4047</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-875,183,-875</points>
<connection>
<GID>5435</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-875,177,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-859.5,177,-859.5</points>
<connection>
<GID>5433</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4048</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-875,208,-875</points>
<connection>
<GID>5439</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-875,202,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-859.5,202,-859.5</points>
<connection>
<GID>5437</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-875,231,-875</points>
<connection>
<GID>5443</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-875,225,-859.5</points>
<intersection>-875 1</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-859.5,225,-859.5</points>
<connection>
<GID>5441</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4050</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-862.5,218,-862.5</points>
<connection>
<GID>5441</GID>
<name>clock</name></connection>
<connection>
<GID>5437</GID>
<name>clock</name></connection>
<connection>
<GID>5433</GID>
<name>clock</name></connection>
<connection>
<GID>5429</GID>
<name>clock</name></connection>
<connection>
<GID>5425</GID>
<name>clock</name></connection>
<connection>
<GID>5421</GID>
<name>clock</name></connection>
<connection>
<GID>5417</GID>
<name>clock</name></connection>
<connection>
<GID>5413</GID>
<name>clock</name></connection>
<connection>
<GID>5409</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4051</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-872,229,-872</points>
<connection>
<GID>5443</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5439</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5435</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5431</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5427</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5423</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5419</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5415</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5411</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4052</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-1009,66,-1009</points>
<connection>
<GID>5452</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-1009,60,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-993.5,60,-993.5</points>
<connection>
<GID>5449</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-1009,89,-1009</points>
<connection>
<GID>5457</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-1009,83,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-993.5,83,-993.5</points>
<connection>
<GID>5454</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-1009,114,-1009</points>
<connection>
<GID>5462</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-1009,108,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-993.5,108,-993.5</points>
<connection>
<GID>5459</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4055</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-1009,137,-1009</points>
<connection>
<GID>5467</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-1009,131,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-993.5,131,-993.5</points>
<connection>
<GID>5464</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4056</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-1009,160,-1009</points>
<connection>
<GID>5472</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-1009,154,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-993.5,154,-993.5</points>
<connection>
<GID>5469</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-1009,183,-1009</points>
<connection>
<GID>5477</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-1009,177,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-993.5,177,-993.5</points>
<connection>
<GID>5474</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4058</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-1009,208,-1009</points>
<connection>
<GID>5544</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-1009,202,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-993.5,202,-993.5</points>
<connection>
<GID>5543</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4059</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-1009,231,-1009</points>
<connection>
<GID>5546</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-1009,225,-993.5</points>
<intersection>-1009 1</intersection>
<intersection>-993.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-993.5,225,-993.5</points>
<connection>
<GID>5545</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-996.5,218,-996.5</points>
<connection>
<GID>5545</GID>
<name>clock</name></connection>
<connection>
<GID>5543</GID>
<name>clock</name></connection>
<connection>
<GID>5474</GID>
<name>clock</name></connection>
<connection>
<GID>5469</GID>
<name>clock</name></connection>
<connection>
<GID>5464</GID>
<name>clock</name></connection>
<connection>
<GID>5459</GID>
<name>clock</name></connection>
<connection>
<GID>5454</GID>
<name>clock</name></connection>
<connection>
<GID>5449</GID>
<name>clock</name></connection>
<connection>
<GID>5445</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-1006,229,-1006</points>
<connection>
<GID>5546</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5544</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5477</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5472</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5467</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5462</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5457</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5452</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5447</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-990.5,66,-990.5</points>
<connection>
<GID>5550</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-990.5,60,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-975,60,-975</points>
<connection>
<GID>5549</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-990.5,89,-990.5</points>
<connection>
<GID>5552</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-990.5,83,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-975,83,-975</points>
<connection>
<GID>5551</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-990.5,114,-990.5</points>
<connection>
<GID>5554</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-990.5,108,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-975,108,-975</points>
<connection>
<GID>5553</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-990.5,137,-990.5</points>
<connection>
<GID>5556</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-990.5,131,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-975,131,-975</points>
<connection>
<GID>5555</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-990.5,160,-990.5</points>
<connection>
<GID>5558</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-990.5,154,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-975,154,-975</points>
<connection>
<GID>5557</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-990.5,183,-990.5</points>
<connection>
<GID>5560</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-990.5,177,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-975,177,-975</points>
<connection>
<GID>5559</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-990.5,208,-990.5</points>
<connection>
<GID>5562</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-990.5,202,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-975,202,-975</points>
<connection>
<GID>5561</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-990.5,231,-990.5</points>
<connection>
<GID>5564</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-990.5,225,-975</points>
<intersection>-990.5 1</intersection>
<intersection>-975 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-975,225,-975</points>
<connection>
<GID>5563</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4070</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-978,218,-978</points>
<connection>
<GID>5563</GID>
<name>clock</name></connection>
<connection>
<GID>5561</GID>
<name>clock</name></connection>
<connection>
<GID>5559</GID>
<name>clock</name></connection>
<connection>
<GID>5557</GID>
<name>clock</name></connection>
<connection>
<GID>5555</GID>
<name>clock</name></connection>
<connection>
<GID>5553</GID>
<name>clock</name></connection>
<connection>
<GID>5551</GID>
<name>clock</name></connection>
<connection>
<GID>5549</GID>
<name>clock</name></connection>
<connection>
<GID>5547</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4071</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-987.5,229,-987.5</points>
<connection>
<GID>5564</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5562</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5560</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5558</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5556</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5554</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5552</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5550</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5548</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-971.5,66,-971.5</points>
<connection>
<GID>5460</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-971.5,60,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-956,60,-956</points>
<connection>
<GID>5455</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-971.5,89,-971.5</points>
<connection>
<GID>5470</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-971.5,83,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-956,83,-956</points>
<connection>
<GID>5465</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4074</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-971.5,114,-971.5</points>
<connection>
<GID>5479</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-971.5,108,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-956,108,-956</points>
<connection>
<GID>5475</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4075</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-971.5,137,-971.5</points>
<connection>
<GID>5566</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-971.5,131,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-956,131,-956</points>
<connection>
<GID>5482</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-971.5,160,-971.5</points>
<connection>
<GID>5568</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-971.5,154,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-956,154,-956</points>
<connection>
<GID>5567</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-971.5,183,-971.5</points>
<connection>
<GID>5570</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-971.5,177,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-956,177,-956</points>
<connection>
<GID>5569</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4078</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-971.5,208,-971.5</points>
<connection>
<GID>5572</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-971.5,202,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-956,202,-956</points>
<connection>
<GID>5571</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4079</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-971.5,231,-971.5</points>
<connection>
<GID>5575</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-971.5,225,-956</points>
<intersection>-971.5 1</intersection>
<intersection>-956 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-956,225,-956</points>
<connection>
<GID>5574</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>4080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-959,218,-959</points>
<connection>
<GID>5574</GID>
<name>clock</name></connection>
<connection>
<GID>5571</GID>
<name>clock</name></connection>
<connection>
<GID>5569</GID>
<name>clock</name></connection>
<connection>
<GID>5567</GID>
<name>clock</name></connection>
<connection>
<GID>5565</GID>
<name>OUT</name></connection>
<connection>
<GID>5482</GID>
<name>clock</name></connection>
<connection>
<GID>5475</GID>
<name>clock</name></connection>
<connection>
<GID>5465</GID>
<name>clock</name></connection>
<connection>
<GID>5455</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4081</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-968.5,229,-968.5</points>
<connection>
<GID>5575</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5572</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5570</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5568</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5566</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5479</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5470</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5460</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5450</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-953,66,-953</points>
<connection>
<GID>5580</GID>
<name>IN_0</name></connection>
<intersection>60 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-953,60,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-937.5,60,-937.5</points>
<connection>
<GID>5579</GID>
<name>OUT_0</name></connection>
<intersection>60 2</intersection></hsegment></shape></wire>
<wire>
<ID>4083</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-953,89,-953</points>
<connection>
<GID>5582</GID>
<name>IN_0</name></connection>
<intersection>83 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,-953,83,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-937.5,83,-937.5</points>
<connection>
<GID>5581</GID>
<name>OUT_0</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>4084</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-953,114,-953</points>
<connection>
<GID>5585</GID>
<name>IN_0</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-953,108,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-937.5,108,-937.5</points>
<connection>
<GID>5584</GID>
<name>OUT_0</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>4085</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-953,137,-953</points>
<connection>
<GID>5587</GID>
<name>IN_0</name></connection>
<intersection>131 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131,-953,131,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-937.5,131,-937.5</points>
<connection>
<GID>5586</GID>
<name>OUT_0</name></connection>
<intersection>131 2</intersection></hsegment></shape></wire>
<wire>
<ID>4086</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-953,160,-953</points>
<connection>
<GID>5590</GID>
<name>IN_0</name></connection>
<intersection>154 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154,-953,154,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-937.5,154,-937.5</points>
<connection>
<GID>5588</GID>
<name>OUT_0</name></connection>
<intersection>154 2</intersection></hsegment></shape></wire>
<wire>
<ID>4087</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-953,183,-953</points>
<connection>
<GID>5592</GID>
<name>IN_0</name></connection>
<intersection>177 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>177,-953,177,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>176,-937.5,177,-937.5</points>
<connection>
<GID>5591</GID>
<name>OUT_0</name></connection>
<intersection>177 2</intersection></hsegment></shape></wire>
<wire>
<ID>4088</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-953,208,-953</points>
<connection>
<GID>5594</GID>
<name>IN_0</name></connection>
<intersection>202 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>202,-953,202,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>201,-937.5,202,-937.5</points>
<connection>
<GID>5593</GID>
<name>OUT_0</name></connection>
<intersection>202 2</intersection></hsegment></shape></wire>
<wire>
<ID>4089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-953,231,-953</points>
<connection>
<GID>5596</GID>
<name>IN_0</name></connection>
<intersection>225 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225,-953,225,-937.5</points>
<intersection>-953 1</intersection>
<intersection>-937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>224,-937.5,225,-937.5</points>
<connection>
<GID>5595</GID>
<name>OUT_0</name></connection>
<intersection>225 2</intersection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-25,68,-25</points>
<connection>
<GID>1447</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-25,62,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-9.5,62,-9.5</points>
<connection>
<GID>1442</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4090</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-940.5,218,-940.5</points>
<connection>
<GID>5595</GID>
<name>clock</name></connection>
<connection>
<GID>5593</GID>
<name>clock</name></connection>
<connection>
<GID>5591</GID>
<name>clock</name></connection>
<connection>
<GID>5588</GID>
<name>clock</name></connection>
<connection>
<GID>5586</GID>
<name>clock</name></connection>
<connection>
<GID>5584</GID>
<name>clock</name></connection>
<connection>
<GID>5581</GID>
<name>clock</name></connection>
<connection>
<GID>5579</GID>
<name>clock</name></connection>
<connection>
<GID>5576</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-25,91,-25</points>
<connection>
<GID>1463</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-25,85,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-9.5,85,-9.5</points>
<connection>
<GID>1462</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4091</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-950,229,-950</points>
<connection>
<GID>5596</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5594</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5592</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5590</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5587</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5585</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5582</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5580</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5577</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-25,116,-25</points>
<connection>
<GID>1465</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-25,110,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-9.5,110,-9.5</points>
<connection>
<GID>1464</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-1019,47.5,-854</points>
<connection>
<GID>5624</GID>
<name>N_in1</name></connection>
<connection>
<GID>5597</GID>
<name>N_in0</name></connection>
<intersection>-993.5 12</intersection>
<intersection>-975 11</intersection>
<intersection>-956 10</intersection>
<intersection>-937.5 9</intersection>
<intersection>-915.5 8</intersection>
<intersection>-897 7</intersection>
<intersection>-878 6</intersection>
<intersection>-859.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-859.5,53,-859.5</points>
<connection>
<GID>5413</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>47.5,-878,53,-878</points>
<connection>
<GID>5740</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>47.5,-897,53,-897</points>
<connection>
<GID>5704</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>47.5,-915.5,53,-915.5</points>
<connection>
<GID>5626</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>47.5,-937.5,53,-937.5</points>
<connection>
<GID>5579</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>47.5,-956,53,-956</points>
<connection>
<GID>5455</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>47.5,-975,53,-975</points>
<connection>
<GID>5549</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>47.5,-993.5,53,-993.5</points>
<connection>
<GID>5449</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-25,139,-25</points>
<connection>
<GID>1467</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-25,133,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-9.5,133,-9.5</points>
<connection>
<GID>1466</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-1018.5,70.5,-853.5</points>
<connection>
<GID>5628</GID>
<name>N_in1</name></connection>
<connection>
<GID>5598</GID>
<name>N_in0</name></connection>
<intersection>-1001 4</intersection>
<intersection>-982.5 5</intersection>
<intersection>-963.5 6</intersection>
<intersection>-945 7</intersection>
<intersection>-923 8</intersection>
<intersection>-904.5 9</intersection>
<intersection>-885.5 10</intersection>
<intersection>-867 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>66,-1001,70.5,-1001</points>
<intersection>66 12</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66,-982.5,70.5,-982.5</points>
<intersection>66 14</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66,-963.5,70.5,-963.5</points>
<intersection>66 13</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66,-945,70.5,-945</points>
<intersection>66 15</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66,-923,70.5,-923</points>
<intersection>66 18</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66,-904.5,70.5,-904.5</points>
<intersection>66 19</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>66,-885.5,70.5,-885.5</points>
<intersection>66 20</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>66,-867,70.5,-867</points>
<intersection>66 21</intersection>
<intersection>70.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>66,-1003.5,66,-1001</points>
<connection>
<GID>5452</GID>
<name>OUT_0</name></connection>
<intersection>-1001 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>66,-966,66,-963.5</points>
<connection>
<GID>5460</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>66,-985,66,-982.5</points>
<connection>
<GID>5550</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>66,-947.5,66,-945</points>
<connection>
<GID>5580</GID>
<name>OUT_0</name></connection>
<intersection>-945 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>66,-925.5,66,-923</points>
<connection>
<GID>5638</GID>
<name>OUT_0</name></connection>
<intersection>-923 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>66,-907,66,-904.5</points>
<connection>
<GID>5706</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>66,-888,66,-885.5</points>
<connection>
<GID>5742</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>66,-869.5,66,-867</points>
<connection>
<GID>5415</GID>
<name>OUT_0</name></connection>
<intersection>-867 11</intersection></vsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-25,162,-25</points>
<connection>
<GID>1469</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-25,156,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-9.5,156,-9.5</points>
<connection>
<GID>1468</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-1018.5,73.5,-854</points>
<connection>
<GID>5630</GID>
<name>N_in1</name></connection>
<connection>
<GID>5599</GID>
<name>N_in0</name></connection>
<intersection>-993.5 10</intersection>
<intersection>-975 9</intersection>
<intersection>-956 8</intersection>
<intersection>-937.5 7</intersection>
<intersection>-915.5 6</intersection>
<intersection>-897 5</intersection>
<intersection>-878 4</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73.5,-859.5,76,-859.5</points>
<connection>
<GID>5417</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-878,76,-878</points>
<connection>
<GID>5744</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>73.5,-897,76,-897</points>
<connection>
<GID>5708</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>73.5,-915.5,76,-915.5</points>
<connection>
<GID>5662</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>73.5,-937.5,76,-937.5</points>
<connection>
<GID>5581</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>73.5,-956,76,-956</points>
<connection>
<GID>5465</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>73.5,-975,76,-975</points>
<connection>
<GID>5551</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>73.5,-993.5,76,-993.5</points>
<connection>
<GID>5454</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-25,185,-25</points>
<connection>
<GID>1471</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-25,179,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-9.5,179,-9.5</points>
<connection>
<GID>1470</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-1018.5,93,-853.5</points>
<connection>
<GID>5632</GID>
<name>N_in1</name></connection>
<connection>
<GID>5600</GID>
<name>N_in0</name></connection>
<intersection>-1001 6</intersection>
<intersection>-982.5 7</intersection>
<intersection>-963.5 8</intersection>
<intersection>-945 9</intersection>
<intersection>-923 10</intersection>
<intersection>-904.5 11</intersection>
<intersection>-885.5 12</intersection>
<intersection>-867 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89,-1001,93,-1001</points>
<intersection>89 14</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89,-982.5,93,-982.5</points>
<intersection>89 16</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89,-963.5,93,-963.5</points>
<intersection>89 15</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89,-945,93,-945</points>
<intersection>89 17</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>89,-923,93,-923</points>
<intersection>89 20</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89,-904.5,93,-904.5</points>
<intersection>89 21</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>89,-885.5,93,-885.5</points>
<intersection>89 22</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>89,-867,93,-867</points>
<intersection>89 23</intersection>
<intersection>93 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>89,-1003.5,89,-1001</points>
<connection>
<GID>5457</GID>
<name>OUT_0</name></connection>
<intersection>-1001 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>89,-966,89,-963.5</points>
<connection>
<GID>5470</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>89,-985,89,-982.5</points>
<connection>
<GID>5552</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>89,-947.5,89,-945</points>
<connection>
<GID>5582</GID>
<name>OUT_0</name></connection>
<intersection>-945 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>89,-925.5,89,-923</points>
<connection>
<GID>5664</GID>
<name>OUT_0</name></connection>
<intersection>-923 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>89,-907,89,-904.5</points>
<connection>
<GID>5710</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>89,-888,89,-885.5</points>
<connection>
<GID>5746</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>89,-869.5,89,-867</points>
<connection>
<GID>5419</GID>
<name>OUT_0</name></connection>
<intersection>-867 13</intersection></vsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-25,210,-25</points>
<connection>
<GID>1473</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-25,204,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-9.5,204,-9.5</points>
<connection>
<GID>1472</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-1018.5,96.5,-853.5</points>
<connection>
<GID>5634</GID>
<name>N_in1</name></connection>
<connection>
<GID>5601</GID>
<name>N_in0</name></connection>
<intersection>-993.5 13</intersection>
<intersection>-975 12</intersection>
<intersection>-956 11</intersection>
<intersection>-937.5 10</intersection>
<intersection>-915.5 9</intersection>
<intersection>-897 8</intersection>
<intersection>-878 7</intersection>
<intersection>-859.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>96.5,-859.5,101,-859.5</points>
<connection>
<GID>5421</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>96.5,-878,101,-878</points>
<connection>
<GID>5748</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>96.5,-897,101,-897</points>
<connection>
<GID>5712</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>96.5,-915.5,101,-915.5</points>
<connection>
<GID>5668</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>96.5,-937.5,101,-937.5</points>
<connection>
<GID>5584</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>96.5,-956,101,-956</points>
<connection>
<GID>5475</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>96.5,-975,101,-975</points>
<connection>
<GID>5553</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>96.5,-993.5,101,-993.5</points>
<connection>
<GID>5459</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-25,233,-25</points>
<connection>
<GID>1475</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-25,227,-9.5</points>
<intersection>-25 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-9.5,227,-9.5</points>
<connection>
<GID>1474</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-1018.5,117.5,-854</points>
<connection>
<GID>5636</GID>
<name>N_in1</name></connection>
<connection>
<GID>5602</GID>
<name>N_in0</name></connection>
<intersection>-1001 6</intersection>
<intersection>-982.5 7</intersection>
<intersection>-963.5 8</intersection>
<intersection>-945 9</intersection>
<intersection>-923 10</intersection>
<intersection>-904.5 11</intersection>
<intersection>-885.5 12</intersection>
<intersection>-867 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>114,-1001,117.5,-1001</points>
<intersection>114 14</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114,-982.5,117.5,-982.5</points>
<intersection>114 16</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114,-963.5,117.5,-963.5</points>
<intersection>114 15</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114,-945,117.5,-945</points>
<intersection>114 17</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114,-923,117.5,-923</points>
<intersection>114 20</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>114,-904.5,117.5,-904.5</points>
<intersection>114 21</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114,-885.5,117.5,-885.5</points>
<intersection>114 22</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>114,-867,117.5,-867</points>
<intersection>114 23</intersection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>114,-1003.5,114,-1001</points>
<connection>
<GID>5462</GID>
<name>OUT_0</name></connection>
<intersection>-1001 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>114,-966,114,-963.5</points>
<connection>
<GID>5479</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>114,-985,114,-982.5</points>
<connection>
<GID>5554</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>114,-947.5,114,-945</points>
<connection>
<GID>5585</GID>
<name>OUT_0</name></connection>
<intersection>-945 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>114,-925.5,114,-923</points>
<connection>
<GID>5672</GID>
<name>OUT_0</name></connection>
<intersection>-923 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>114,-907,114,-904.5</points>
<connection>
<GID>5714</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>114,-888,114,-885.5</points>
<connection>
<GID>5750</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>114,-869.5,114,-867</points>
<connection>
<GID>5423</GID>
<name>OUT_0</name></connection>
<intersection>-867 13</intersection></vsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-12.5,220,-12.5</points>
<connection>
<GID>1474</GID>
<name>clock</name></connection>
<connection>
<GID>1472</GID>
<name>clock</name></connection>
<connection>
<GID>1470</GID>
<name>clock</name></connection>
<connection>
<GID>1468</GID>
<name>clock</name></connection>
<connection>
<GID>1466</GID>
<name>clock</name></connection>
<connection>
<GID>1464</GID>
<name>clock</name></connection>
<connection>
<GID>1462</GID>
<name>clock</name></connection>
<connection>
<GID>1442</GID>
<name>clock</name></connection>
<connection>
<GID>1434</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-1018.5,121.5,-853.5</points>
<connection>
<GID>5640</GID>
<name>N_in1</name></connection>
<connection>
<GID>5603</GID>
<name>N_in0</name></connection>
<intersection>-993.5 13</intersection>
<intersection>-975 12</intersection>
<intersection>-956 11</intersection>
<intersection>-937.5 10</intersection>
<intersection>-915.5 9</intersection>
<intersection>-897 8</intersection>
<intersection>-878 7</intersection>
<intersection>-859.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>121.5,-859.5,124,-859.5</points>
<connection>
<GID>5425</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>121.5,-878,124,-878</points>
<connection>
<GID>5752</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121.5,-897,124,-897</points>
<connection>
<GID>5716</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>121.5,-915.5,124,-915.5</points>
<connection>
<GID>5676</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>121.5,-937.5,124,-937.5</points>
<connection>
<GID>5586</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>121.5,-956,124,-956</points>
<connection>
<GID>5482</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>121.5,-975,124,-975</points>
<connection>
<GID>5555</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>121.5,-993.5,124,-993.5</points>
<connection>
<GID>5464</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-22,231,-22</points>
<connection>
<GID>1447</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1463</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1465</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1467</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1469</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1471</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1473</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1475</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1438</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-1018.5,140,-853.5</points>
<connection>
<GID>5642</GID>
<name>N_in1</name></connection>
<connection>
<GID>5604</GID>
<name>N_in0</name></connection>
<intersection>-1001 6</intersection>
<intersection>-982.5 7</intersection>
<intersection>-963.5 8</intersection>
<intersection>-945 9</intersection>
<intersection>-923 10</intersection>
<intersection>-904.5 11</intersection>
<intersection>-885.5 12</intersection>
<intersection>-867 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>137,-1001,140,-1001</points>
<intersection>137 14</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137,-982.5,140,-982.5</points>
<intersection>137 15</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-963.5,140,-963.5</points>
<intersection>137 16</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137,-945,140,-945</points>
<intersection>137 17</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-923,140,-923</points>
<intersection>137 20</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>137,-904.5,140,-904.5</points>
<intersection>137 21</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137,-885.5,140,-885.5</points>
<intersection>137 22</intersection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-867,140,-867</points>
<intersection>137 23</intersection>
<intersection>140 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>137,-1003.5,137,-1001</points>
<connection>
<GID>5467</GID>
<name>OUT_0</name></connection>
<intersection>-1001 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>137,-985,137,-982.5</points>
<connection>
<GID>5556</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>137,-966,137,-963.5</points>
<connection>
<GID>5566</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>137,-947.5,137,-945</points>
<connection>
<GID>5587</GID>
<name>OUT_0</name></connection>
<intersection>-945 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>137,-925.5,137,-923</points>
<connection>
<GID>5680</GID>
<name>OUT_0</name></connection>
<intersection>-923 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>137,-907,137,-904.5</points>
<connection>
<GID>5718</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>137,-888,137,-885.5</points>
<connection>
<GID>5754</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>137,-869.5,137,-867</points>
<connection>
<GID>5427</GID>
<name>OUT_0</name></connection>
<intersection>-867 13</intersection></vsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-6.5,68,-6.5</points>
<connection>
<GID>1479</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-6.5,62,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,9,62,9</points>
<connection>
<GID>1478</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-1018.5,144,-853.5</points>
<connection>
<GID>5644</GID>
<name>N_in1</name></connection>
<connection>
<GID>5606</GID>
<name>N_in0</name></connection>
<intersection>-993.5 13</intersection>
<intersection>-975 12</intersection>
<intersection>-956 11</intersection>
<intersection>-937.5 10</intersection>
<intersection>-915.5 9</intersection>
<intersection>-897 8</intersection>
<intersection>-878 7</intersection>
<intersection>-859.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>144,-859.5,147,-859.5</points>
<connection>
<GID>5429</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>144,-878,147,-878</points>
<connection>
<GID>5756</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>144,-897,147,-897</points>
<connection>
<GID>5720</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>144,-915.5,147,-915.5</points>
<connection>
<GID>5682</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>144,-937.5,147,-937.5</points>
<connection>
<GID>5588</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>144,-956,147,-956</points>
<connection>
<GID>5567</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>144,-975,147,-975</points>
<connection>
<GID>5557</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>144,-993.5,147,-993.5</points>
<connection>
<GID>5469</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-6.5,91,-6.5</points>
<connection>
<GID>1481</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-6.5,85,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,9,85,9</points>
<connection>
<GID>1480</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-1018,163,-853.5</points>
<connection>
<GID>5646</GID>
<name>N_in1</name></connection>
<connection>
<GID>5608</GID>
<name>N_in0</name></connection>
<intersection>-1001 6</intersection>
<intersection>-982.5 7</intersection>
<intersection>-963.5 8</intersection>
<intersection>-945 9</intersection>
<intersection>-923 10</intersection>
<intersection>-904.5 11</intersection>
<intersection>-885.5 12</intersection>
<intersection>-867 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>160,-1001,163,-1001</points>
<intersection>160 15</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>160,-982.5,163,-982.5</points>
<intersection>160 16</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>160,-963.5,163,-963.5</points>
<intersection>160 17</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>160,-945,163,-945</points>
<intersection>160 18</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>160,-923,163,-923</points>
<intersection>160 21</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>160,-904.5,163,-904.5</points>
<intersection>160 22</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>160,-885.5,163,-885.5</points>
<intersection>160 23</intersection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>160,-867,163,-867</points>
<intersection>160 14</intersection>
<intersection>163 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>160,-869.5,160,-867</points>
<connection>
<GID>5431</GID>
<name>OUT_0</name></connection>
<intersection>-867 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>160,-1003.5,160,-1001</points>
<connection>
<GID>5472</GID>
<name>OUT_0</name></connection>
<intersection>-1001 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>160,-985,160,-982.5</points>
<connection>
<GID>5558</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>160,-966,160,-963.5</points>
<connection>
<GID>5568</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>160,-947.5,160,-945</points>
<connection>
<GID>5590</GID>
<name>OUT_0</name></connection>
<intersection>-945 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>160,-925.5,160,-923</points>
<connection>
<GID>5686</GID>
<name>OUT_0</name></connection>
<intersection>-923 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>160,-907,160,-904.5</points>
<connection>
<GID>5722</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>160,-888,160,-885.5</points>
<connection>
<GID>5395</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 12</intersection></vsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-6.5,116,-6.5</points>
<connection>
<GID>1483</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-6.5,110,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,9,110,9</points>
<connection>
<GID>1482</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-1018,168,-853.5</points>
<connection>
<GID>5648</GID>
<name>N_in1</name></connection>
<connection>
<GID>5610</GID>
<name>N_in0</name></connection>
<intersection>-993.5 13</intersection>
<intersection>-975 12</intersection>
<intersection>-956 11</intersection>
<intersection>-937.5 10</intersection>
<intersection>-915.5 9</intersection>
<intersection>-897 8</intersection>
<intersection>-878 7</intersection>
<intersection>-859.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>168,-859.5,170,-859.5</points>
<connection>
<GID>5433</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>168,-878,170,-878</points>
<connection>
<GID>5397</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>168,-897,170,-897</points>
<connection>
<GID>5724</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>168,-915.5,170,-915.5</points>
<connection>
<GID>5688</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>168,-937.5,170,-937.5</points>
<connection>
<GID>5591</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>168,-956,170,-956</points>
<connection>
<GID>5569</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>168,-975,170,-975</points>
<connection>
<GID>5559</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>168,-993.5,170,-993.5</points>
<connection>
<GID>5474</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-6.5,139,-6.5</points>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-6.5,133,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,9,133,9</points>
<connection>
<GID>1484</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-1017.5,186,-853.5</points>
<connection>
<GID>5650</GID>
<name>N_in1</name></connection>
<connection>
<GID>5614</GID>
<name>N_in0</name></connection>
<intersection>-1001 16</intersection>
<intersection>-982.5 15</intersection>
<intersection>-963.5 14</intersection>
<intersection>-945 13</intersection>
<intersection>-923 12</intersection>
<intersection>-904.5 11</intersection>
<intersection>-885.5 10</intersection>
<intersection>-867 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>183,-867,186,-867</points>
<intersection>183 17</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183,-885.5,186,-885.5</points>
<intersection>183 26</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183,-904.5,186,-904.5</points>
<intersection>183 25</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183,-923,186,-923</points>
<intersection>183 24</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183,-945,186,-945</points>
<intersection>183 21</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>183,-963.5,186,-963.5</points>
<intersection>183 20</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>183,-982.5,186,-982.5</points>
<intersection>183 19</intersection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>183,-1001,186,-1001</points>
<intersection>183 18</intersection>
<intersection>186 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>183,-869.5,183,-867</points>
<connection>
<GID>5435</GID>
<name>OUT_0</name></connection>
<intersection>-867 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>183,-1003.5,183,-1001</points>
<connection>
<GID>5477</GID>
<name>OUT_0</name></connection>
<intersection>-1001 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>183,-985,183,-982.5</points>
<connection>
<GID>5560</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>183,-966,183,-963.5</points>
<connection>
<GID>5570</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>183,-947.5,183,-945</points>
<connection>
<GID>5592</GID>
<name>OUT_0</name></connection>
<intersection>-945 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>183,-925.5,183,-923</points>
<connection>
<GID>5690</GID>
<name>OUT_0</name></connection>
<intersection>-923 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>183,-907,183,-904.5</points>
<connection>
<GID>5726</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>183,-888,183,-885.5</points>
<connection>
<GID>5399</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-6.5,162,-6.5</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-6.5,156,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,9,156,9</points>
<connection>
<GID>1486</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-1017.5,190.5,-853.5</points>
<connection>
<GID>5652</GID>
<name>N_in1</name></connection>
<connection>
<GID>5612</GID>
<name>N_in0</name></connection>
<intersection>-993.5 13</intersection>
<intersection>-975 12</intersection>
<intersection>-956 11</intersection>
<intersection>-937.5 10</intersection>
<intersection>-915.5 9</intersection>
<intersection>-897 8</intersection>
<intersection>-878 7</intersection>
<intersection>-859.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>190.5,-859.5,195,-859.5</points>
<connection>
<GID>5437</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>190.5,-878,195,-878</points>
<connection>
<GID>5401</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>190.5,-897,195,-897</points>
<connection>
<GID>5728</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>190.5,-915.5,195,-915.5</points>
<connection>
<GID>5692</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>190.5,-937.5,195,-937.5</points>
<connection>
<GID>5593</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>190.5,-956,195,-956</points>
<connection>
<GID>5571</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>190.5,-975,195,-975</points>
<connection>
<GID>5561</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>190.5,-993.5,195,-993.5</points>
<connection>
<GID>5543</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-6.5,185,-6.5</points>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-6.5,179,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,9,179,9</points>
<connection>
<GID>1488</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,-1017,211.5,-854</points>
<connection>
<GID>5654</GID>
<name>N_in1</name></connection>
<connection>
<GID>5616</GID>
<name>N_in0</name></connection>
<intersection>-1001 6</intersection>
<intersection>-982.5 7</intersection>
<intersection>-963.5 8</intersection>
<intersection>-945 9</intersection>
<intersection>-923 10</intersection>
<intersection>-904.5 11</intersection>
<intersection>-885.5 12</intersection>
<intersection>-867 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>208,-1001,211.5,-1001</points>
<intersection>208 15</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>208,-982.5,211.5,-982.5</points>
<intersection>208 16</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>208,-963.5,211.5,-963.5</points>
<intersection>208 17</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>208,-945,211.5,-945</points>
<intersection>208 18</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>208,-923,211.5,-923</points>
<intersection>208 21</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>208,-904.5,211.5,-904.5</points>
<intersection>208 22</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>208,-885.5,211.5,-885.5</points>
<intersection>208 23</intersection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>208,-867,211.5,-867</points>
<intersection>208 14</intersection>
<intersection>211.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>208,-869.5,208,-867</points>
<connection>
<GID>5439</GID>
<name>OUT_0</name></connection>
<intersection>-867 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>208,-1003.5,208,-1001</points>
<connection>
<GID>5544</GID>
<name>OUT_0</name></connection>
<intersection>-1001 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>208,-985,208,-982.5</points>
<connection>
<GID>5562</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>208,-966,208,-963.5</points>
<connection>
<GID>5572</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>208,-947.5,208,-945</points>
<connection>
<GID>5594</GID>
<name>OUT_0</name></connection>
<intersection>-945 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>208,-925.5,208,-923</points>
<connection>
<GID>5694</GID>
<name>OUT_0</name></connection>
<intersection>-923 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>208,-907,208,-904.5</points>
<connection>
<GID>5730</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>208,-888,208,-885.5</points>
<connection>
<GID>5403</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 12</intersection></vsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-6.5,210,-6.5</points>
<connection>
<GID>1491</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-6.5,204,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,9,204,9</points>
<connection>
<GID>1490</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215,-1017,215,-854</points>
<connection>
<GID>5656</GID>
<name>N_in1</name></connection>
<connection>
<GID>5658</GID>
<name>N_in0</name></connection>
<intersection>-993.5 11</intersection>
<intersection>-975 10</intersection>
<intersection>-956 9</intersection>
<intersection>-937.5 7</intersection>
<intersection>-915.5 6</intersection>
<intersection>-897 5</intersection>
<intersection>-878 4</intersection>
<intersection>-859.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-859.5,218,-859.5</points>
<connection>
<GID>5441</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>215,-878,218,-878</points>
<connection>
<GID>5405</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>215,-897,218,-897</points>
<connection>
<GID>5732</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>215,-915.5,218,-915.5</points>
<connection>
<GID>5696</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>215,-937.5,218,-937.5</points>
<connection>
<GID>5595</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>215,-956,218,-956</points>
<connection>
<GID>5574</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>215,-975,218,-975</points>
<connection>
<GID>5563</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>215,-993.5,218,-993.5</points>
<connection>
<GID>5545</GID>
<name>IN_0</name></connection>
<intersection>215 0</intersection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-6.5,233,-6.5</points>
<connection>
<GID>1493</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-6.5,227,9</points>
<intersection>-6.5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,9,227,9</points>
<connection>
<GID>1492</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-1017,236,-855</points>
<connection>
<GID>5660</GID>
<name>N_in1</name></connection>
<connection>
<GID>5618</GID>
<name>N_in0</name></connection>
<intersection>-1001 11</intersection>
<intersection>-982.5 10</intersection>
<intersection>-963.5 9</intersection>
<intersection>-945 8</intersection>
<intersection>-923 7</intersection>
<intersection>-904.5 6</intersection>
<intersection>-885.5 5</intersection>
<intersection>-867 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>231,-867,236,-867</points>
<intersection>231 12</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>231,-885.5,236,-885.5</points>
<intersection>231 21</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>231,-904.5,236,-904.5</points>
<intersection>231 20</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>231,-923,236,-923</points>
<intersection>231 19</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>231,-945,236,-945</points>
<intersection>231 16</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>231,-963.5,236,-963.5</points>
<intersection>231 15</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>231,-982.5,236,-982.5</points>
<intersection>231 14</intersection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>231,-1001,236,-1001</points>
<intersection>231 13</intersection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>231,-869.5,231,-867</points>
<connection>
<GID>5443</GID>
<name>OUT_0</name></connection>
<intersection>-867 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>231,-1003.5,231,-1001</points>
<connection>
<GID>5546</GID>
<name>OUT_0</name></connection>
<intersection>-1001 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>231,-985,231,-982.5</points>
<connection>
<GID>5564</GID>
<name>OUT_0</name></connection>
<intersection>-982.5 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>231,-966,231,-963.5</points>
<connection>
<GID>5575</GID>
<name>OUT_0</name></connection>
<intersection>-963.5 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>231,-947.5,231,-945</points>
<connection>
<GID>5596</GID>
<name>OUT_0</name></connection>
<intersection>-945 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>231,-925.5,231,-923</points>
<connection>
<GID>5698</GID>
<name>OUT_0</name></connection>
<intersection>-923 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>231,-907,231,-904.5</points>
<connection>
<GID>5734</GID>
<name>OUT_0</name></connection>
<intersection>-904.5 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>231,-888,231,-885.5</points>
<connection>
<GID>5407</GID>
<name>OUT_0</name></connection>
<intersection>-885.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,6,220,6</points>
<connection>
<GID>1476</GID>
<name>OUT</name></connection>
<connection>
<GID>1478</GID>
<name>clock</name></connection>
<connection>
<GID>1480</GID>
<name>clock</name></connection>
<connection>
<GID>1482</GID>
<name>clock</name></connection>
<connection>
<GID>1484</GID>
<name>clock</name></connection>
<connection>
<GID>1486</GID>
<name>clock</name></connection>
<connection>
<GID>1488</GID>
<name>clock</name></connection>
<connection>
<GID>1490</GID>
<name>clock</name></connection>
<connection>
<GID>1492</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4108</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-114,-861.5,25.5,-861.5</points>
<connection>
<GID>5409</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114,-871,-114,-845.5</points>
<intersection>-871 4</intersection>
<intersection>-861.5 2</intersection>
<intersection>-845.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-114,-871,37,-871</points>
<connection>
<GID>5411</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-121,-845.5,-114,-845.5</points>
<connection>
<GID>5542</GID>
<name>OUT_7</name></connection>
<intersection>-114 3</intersection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-3.5,231,-3.5</points>
<connection>
<GID>1493</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1491</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1489</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1487</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1485</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1483</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1481</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1479</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1477</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4109</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-115,-880,25.5,-880</points>
<connection>
<GID>5736</GID>
<name>IN_0</name></connection>
<intersection>-115 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-115,-889.5,-115,-846.5</points>
<intersection>-889.5 5</intersection>
<intersection>-880 2</intersection>
<intersection>-846.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-115,-889.5,37,-889.5</points>
<connection>
<GID>5738</GID>
<name>IN_0</name></connection>
<intersection>-115 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-121,-846.5,-115,-846.5</points>
<connection>
<GID>5542</GID>
<name>OUT_6</name></connection>
<intersection>-115 4</intersection></hsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,12.5,68,12.5</points>
<connection>
<GID>1497</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,12.5,62,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,28,62,28</points>
<connection>
<GID>1496</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4110</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-116,-899,25.5,-899</points>
<connection>
<GID>5700</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-116,-908.5,-116,-847.5</points>
<intersection>-908.5 4</intersection>
<intersection>-899 2</intersection>
<intersection>-847.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-116,-908.5,37,-908.5</points>
<connection>
<GID>5702</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-121,-847.5,-116,-847.5</points>
<connection>
<GID>5542</GID>
<name>OUT_5</name></connection>
<intersection>-116 3</intersection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,12.5,91,12.5</points>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,12.5,85,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,28,85,28</points>
<connection>
<GID>1498</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4111</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-117,-917.5,25.5,-917.5</points>
<connection>
<GID>5620</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-927,-117,-848.5</points>
<intersection>-927 4</intersection>
<intersection>-917.5 2</intersection>
<intersection>-848.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-927,37,-927</points>
<connection>
<GID>5622</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-848.5,-117,-848.5</points>
<connection>
<GID>5542</GID>
<name>OUT_4</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,12.5,116,12.5</points>
<connection>
<GID>1501</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,12.5,110,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,28,110,28</points>
<connection>
<GID>1500</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118,-939.5,25.5,-939.5</points>
<connection>
<GID>5576</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118,-949,-118,-849.5</points>
<intersection>-949 4</intersection>
<intersection>-939.5 1</intersection>
<intersection>-849.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118,-949,36.5,-949</points>
<connection>
<GID>5577</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-849.5,-118,-849.5</points>
<connection>
<GID>5542</GID>
<name>OUT_3</name></connection>
<intersection>-118 3</intersection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,12.5,139,12.5</points>
<connection>
<GID>1503</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,12.5,133,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,28,133,28</points>
<connection>
<GID>1502</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,-958,25.5,-958</points>
<connection>
<GID>5565</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-967.5,-119,-850.5</points>
<intersection>-967.5 4</intersection>
<intersection>-958 1</intersection>
<intersection>-850.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-967.5,36.5,-967.5</points>
<connection>
<GID>5450</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-850.5,-119,-850.5</points>
<connection>
<GID>5542</GID>
<name>OUT_2</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,12.5,162,12.5</points>
<connection>
<GID>1505</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,12.5,156,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,28,156,28</points>
<connection>
<GID>1504</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-977,25.5,-977</points>
<connection>
<GID>5547</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-986.5,-120,-851.5</points>
<intersection>-986.5 4</intersection>
<intersection>-977 1</intersection>
<intersection>-851.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-120,-986.5,36.5,-986.5</points>
<connection>
<GID>5548</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-121,-851.5,-120,-851.5</points>
<connection>
<GID>5542</GID>
<name>OUT_1</name></connection>
<intersection>-120 3</intersection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,12.5,185,12.5</points>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,12.5,179,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,28,179,28</points>
<connection>
<GID>1506</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-995.5,25.5,-995.5</points>
<connection>
<GID>5445</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-1005,-121,-852.5</points>
<connection>
<GID>5542</GID>
<name>OUT_0</name></connection>
<intersection>-1005 4</intersection>
<intersection>-995.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-1005,36.5,-1005</points>
<connection>
<GID>5447</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,12.5,210,12.5</points>
<connection>
<GID>1509</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,12.5,204,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,28,204,28</points>
<connection>
<GID>1508</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-1019,24.5,-854</points>
<connection>
<GID>5678</GID>
<name>N_in1</name></connection>
<connection>
<GID>5670</GID>
<name>N_in0</name></connection>
<intersection>-997.5 10</intersection>
<intersection>-979 9</intersection>
<intersection>-960 8</intersection>
<intersection>-941.5 7</intersection>
<intersection>-919.5 6</intersection>
<intersection>-901 5</intersection>
<intersection>-882 4</intersection>
<intersection>-863.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-863.5,25.5,-863.5</points>
<connection>
<GID>5409</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-882,25.5,-882</points>
<connection>
<GID>5736</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>24.5,-901,25.5,-901</points>
<connection>
<GID>5700</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>24.5,-919.5,25.5,-919.5</points>
<connection>
<GID>5620</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>24.5,-941.5,25.5,-941.5</points>
<connection>
<GID>5576</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>24.5,-960,25.5,-960</points>
<connection>
<GID>5565</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>24.5,-979,25.5,-979</points>
<connection>
<GID>5547</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>24.5,-997.5,25.5,-997.5</points>
<connection>
<GID>5445</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,12.5,233,12.5</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,12.5,227,28</points>
<intersection>12.5 1</intersection>
<intersection>28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,28,227,28</points>
<connection>
<GID>1510</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-1019,34.5,-854</points>
<connection>
<GID>5674</GID>
<name>N_in1</name></connection>
<connection>
<GID>5666</GID>
<name>N_in0</name></connection>
<intersection>-1007 3</intersection>
<intersection>-988.5 5</intersection>
<intersection>-969.5 7</intersection>
<intersection>-951 9</intersection>
<intersection>-929 11</intersection>
<intersection>-910.5 13</intersection>
<intersection>-891.5 15</intersection>
<intersection>-873 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34.5,-1007,36.5,-1007</points>
<connection>
<GID>5447</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>34.5,-988.5,36.5,-988.5</points>
<connection>
<GID>5548</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>34.5,-969.5,36.5,-969.5</points>
<connection>
<GID>5450</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>34.5,-951,36.5,-951</points>
<connection>
<GID>5577</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>34.5,-929,37,-929</points>
<connection>
<GID>5622</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>34.5,-910.5,37,-910.5</points>
<connection>
<GID>5702</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>34.5,-891.5,37,-891.5</points>
<connection>
<GID>5738</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>34.5,-873,37,-873</points>
<connection>
<GID>5411</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,25,220,25</points>
<connection>
<GID>1510</GID>
<name>clock</name></connection>
<connection>
<GID>1508</GID>
<name>clock</name></connection>
<connection>
<GID>1506</GID>
<name>clock</name></connection>
<connection>
<GID>1504</GID>
<name>clock</name></connection>
<connection>
<GID>1502</GID>
<name>clock</name></connection>
<connection>
<GID>1500</GID>
<name>clock</name></connection>
<connection>
<GID>1498</GID>
<name>clock</name></connection>
<connection>
<GID>1496</GID>
<name>clock</name></connection>
<connection>
<GID>1494</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-852,24.5,-845.5</points>
<connection>
<GID>5670</GID>
<name>N_in1</name></connection>
<connection>
<GID>5540</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,15.5,231,15.5</points>
<connection>
<GID>1497</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1499</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1501</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1503</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1505</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1507</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1509</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1511</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1495</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-852,34.5,-845.5</points>
<connection>
<GID>5666</GID>
<name>N_in1</name></connection>
<connection>
<GID>5539</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,31,68,31</points>
<connection>
<GID>1515</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,31,62,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,46.5,62,46.5</points>
<connection>
<GID>1514</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-852,47.5,-845.5</points>
<connection>
<GID>5597</GID>
<name>N_in1</name></connection>
<connection>
<GID>5520</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,31,91,31</points>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,31,85,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,46.5,85,46.5</points>
<connection>
<GID>1516</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-851.5,70.5,-845</points>
<connection>
<GID>5598</GID>
<name>N_in1</name></connection>
<connection>
<GID>5521</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,31,116,31</points>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,31,110,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,46.5,110,46.5</points>
<connection>
<GID>1518</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-852,73.5,-845</points>
<connection>
<GID>5599</GID>
<name>N_in1</name></connection>
<connection>
<GID>5522</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,31,139,31</points>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,31,133,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,46.5,133,46.5</points>
<connection>
<GID>1520</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-851.5,93,-845</points>
<connection>
<GID>5600</GID>
<name>N_in1</name></connection>
<connection>
<GID>5523</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,31,162,31</points>
<connection>
<GID>1523</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,31,156,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,46.5,156,46.5</points>
<connection>
<GID>1522</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-851.5,96.5,-845</points>
<connection>
<GID>5601</GID>
<name>N_in1</name></connection>
<connection>
<GID>5524</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,31,185,31</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,31,179,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,46.5,179,46.5</points>
<connection>
<GID>1524</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-852,117.5,-845</points>
<connection>
<GID>5602</GID>
<name>N_in1</name></connection>
<connection>
<GID>5525</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,31,210,31</points>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,31,204,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,46.5,204,46.5</points>
<connection>
<GID>1526</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-851.5,121.5,-845</points>
<connection>
<GID>5603</GID>
<name>N_in1</name></connection>
<connection>
<GID>5526</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,31,233,31</points>
<connection>
<GID>1529</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,31,227,46.5</points>
<intersection>31 1</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,46.5,227,46.5</points>
<connection>
<GID>1528</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-851.5,140,-845</points>
<connection>
<GID>5604</GID>
<name>N_in1</name></connection>
<connection>
<GID>5527</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,43.5,220,43.5</points>
<connection>
<GID>1528</GID>
<name>clock</name></connection>
<connection>
<GID>1526</GID>
<name>clock</name></connection>
<connection>
<GID>1524</GID>
<name>clock</name></connection>
<connection>
<GID>1522</GID>
<name>clock</name></connection>
<connection>
<GID>1520</GID>
<name>clock</name></connection>
<connection>
<GID>1518</GID>
<name>clock</name></connection>
<connection>
<GID>1516</GID>
<name>clock</name></connection>
<connection>
<GID>1514</GID>
<name>clock</name></connection>
<connection>
<GID>1512</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-851.5,144,-845</points>
<connection>
<GID>5606</GID>
<name>N_in1</name></connection>
<connection>
<GID>5528</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,34,231,34</points>
<connection>
<GID>1515</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1517</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1519</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1521</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1523</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1525</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1527</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1529</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1513</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-851.5,163,-844.5</points>
<connection>
<GID>5608</GID>
<name>N_in1</name></connection>
<connection>
<GID>5529</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-103,68,-103</points>
<connection>
<GID>1533</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-103,62,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-87.5,62,-87.5</points>
<connection>
<GID>1532</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-851.5,168,-844.5</points>
<connection>
<GID>5610</GID>
<name>N_in1</name></connection>
<connection>
<GID>5530</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-103,91,-103</points>
<connection>
<GID>1535</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-103,85,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-87.5,85,-87.5</points>
<connection>
<GID>1534</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-851.5,186,-844</points>
<connection>
<GID>5614</GID>
<name>N_in1</name></connection>
<connection>
<GID>5531</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-103,116,-103</points>
<connection>
<GID>1537</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-103,110,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-87.5,110,-87.5</points>
<connection>
<GID>1536</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-851.5,190.5,-844</points>
<connection>
<GID>5612</GID>
<name>N_in1</name></connection>
<connection>
<GID>5532</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-103,139,-103</points>
<connection>
<GID>1539</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-103,133,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-87.5,133,-87.5</points>
<connection>
<GID>1538</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,-852,211.5,-843.5</points>
<connection>
<GID>5616</GID>
<name>N_in1</name></connection>
<connection>
<GID>5533</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-103,162,-103</points>
<connection>
<GID>1541</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-103,156,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-87.5,156,-87.5</points>
<connection>
<GID>1540</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215,-852,215,-843.5</points>
<connection>
<GID>5658</GID>
<name>N_in1</name></connection>
<connection>
<GID>5534</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-103,185,-103</points>
<connection>
<GID>1543</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-103,179,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-87.5,179,-87.5</points>
<connection>
<GID>1542</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-853,236,-843.5</points>
<connection>
<GID>5618</GID>
<name>N_in1</name></connection>
<connection>
<GID>5536</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-103,210,-103</points>
<connection>
<GID>1545</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-103,204,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-87.5,204,-87.5</points>
<connection>
<GID>1544</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1138,63,-1138</points>
<connection>
<GID>5954</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1138,57,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1122.5,57,-1122.5</points>
<connection>
<GID>5948</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-103,233,-103</points>
<connection>
<GID>1547</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-103,227,-87.5</points>
<intersection>-103 1</intersection>
<intersection>-87.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-87.5,227,-87.5</points>
<connection>
<GID>1546</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1138,86,-1138</points>
<connection>
<GID>5972</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1138,80,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1122.5,80,-1122.5</points>
<connection>
<GID>5970</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-90.5,220,-90.5</points>
<connection>
<GID>1542</GID>
<name>clock</name></connection>
<connection>
<GID>1540</GID>
<name>clock</name></connection>
<connection>
<GID>1538</GID>
<name>clock</name></connection>
<connection>
<GID>1536</GID>
<name>clock</name></connection>
<connection>
<GID>1534</GID>
<name>clock</name></connection>
<connection>
<GID>1532</GID>
<name>clock</name></connection>
<connection>
<GID>1530</GID>
<name>OUT</name></connection>
<connection>
<GID>1546</GID>
<name>clock</name></connection>
<connection>
<GID>1544</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1138,111,-1138</points>
<connection>
<GID>5976</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1138,105,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1122.5,105,-1122.5</points>
<connection>
<GID>5974</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-100,231,-100</points>
<connection>
<GID>1545</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1547</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1533</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1535</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1537</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1539</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1541</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1543</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1531</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1138,134,-1138</points>
<connection>
<GID>5980</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1138,128,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1122.5,128,-1122.5</points>
<connection>
<GID>5978</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-84.5,68,-84.5</points>
<connection>
<GID>1551</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-84.5,62,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-69,62,-69</points>
<connection>
<GID>1550</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1138,157,-1138</points>
<connection>
<GID>5984</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1138,151,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1122.5,151,-1122.5</points>
<connection>
<GID>5982</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-84.5,91,-84.5</points>
<connection>
<GID>1553</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-84.5,85,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-69,85,-69</points>
<connection>
<GID>1552</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1138,180,-1138</points>
<connection>
<GID>5988</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1138,174,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1122.5,174,-1122.5</points>
<connection>
<GID>5986</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-84.5,116,-84.5</points>
<connection>
<GID>1555</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-84.5,110,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-69,110,-69</points>
<connection>
<GID>1554</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1138,205,-1138</points>
<connection>
<GID>5992</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1138,199,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1122.5,199,-1122.5</points>
<connection>
<GID>5990</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-84.5,139,-84.5</points>
<connection>
<GID>1557</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-84.5,133,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-69,133,-69</points>
<connection>
<GID>1556</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1138,228,-1138</points>
<connection>
<GID>5996</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1138,222,-1122.5</points>
<intersection>-1138 1</intersection>
<intersection>-1122.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1122.5,222,-1122.5</points>
<connection>
<GID>5994</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-84.5,162,-84.5</points>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-84.5,156,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-69,156,-69</points>
<connection>
<GID>1558</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1125.5,215,-1125.5</points>
<connection>
<GID>5994</GID>
<name>clock</name></connection>
<connection>
<GID>5990</GID>
<name>clock</name></connection>
<connection>
<GID>5986</GID>
<name>clock</name></connection>
<connection>
<GID>5982</GID>
<name>clock</name></connection>
<connection>
<GID>5978</GID>
<name>clock</name></connection>
<connection>
<GID>5974</GID>
<name>clock</name></connection>
<connection>
<GID>5970</GID>
<name>clock</name></connection>
<connection>
<GID>5948</GID>
<name>clock</name></connection>
<connection>
<GID>5938</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-84.5,185,-84.5</points>
<connection>
<GID>1561</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-84.5,179,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-69,179,-69</points>
<connection>
<GID>1560</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1135,226,-1135</points>
<connection>
<GID>5996</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5992</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5988</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5984</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5980</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5976</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5972</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5954</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5943</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-84.5,210,-84.5</points>
<connection>
<GID>1563</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-84.5,204,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-69,204,-69</points>
<connection>
<GID>1562</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1119.5,63,-1119.5</points>
<connection>
<GID>6004</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1119.5,57,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1104,57,-1104</points>
<connection>
<GID>6002</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-84.5,233,-84.5</points>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-84.5,227,-69</points>
<intersection>-84.5 1</intersection>
<intersection>-69 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-69,227,-69</points>
<connection>
<GID>1564</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1119.5,86,-1119.5</points>
<connection>
<GID>6008</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1119.5,80,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1104,80,-1104</points>
<connection>
<GID>6006</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-72,220,-72</points>
<connection>
<GID>1548</GID>
<name>OUT</name></connection>
<connection>
<GID>1550</GID>
<name>clock</name></connection>
<connection>
<GID>1552</GID>
<name>clock</name></connection>
<connection>
<GID>1554</GID>
<name>clock</name></connection>
<connection>
<GID>1556</GID>
<name>clock</name></connection>
<connection>
<GID>1558</GID>
<name>clock</name></connection>
<connection>
<GID>1560</GID>
<name>clock</name></connection>
<connection>
<GID>1562</GID>
<name>clock</name></connection>
<connection>
<GID>1564</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1119.5,111,-1119.5</points>
<connection>
<GID>6012</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1119.5,105,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1104,105,-1104</points>
<connection>
<GID>6010</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-81.5,231,-81.5</points>
<connection>
<GID>1551</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1553</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1555</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1557</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1559</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1561</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1563</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1565</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1549</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1119.5,134,-1119.5</points>
<connection>
<GID>6016</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1119.5,128,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1104,128,-1104</points>
<connection>
<GID>6014</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-65.5,68,-65.5</points>
<connection>
<GID>1569</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-65.5,62,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-50,62,-50</points>
<connection>
<GID>1568</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1119.5,157,-1119.5</points>
<connection>
<GID>6020</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1119.5,151,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1104,151,-1104</points>
<connection>
<GID>6018</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-65.5,91,-65.5</points>
<connection>
<GID>1571</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-65.5,85,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-50,85,-50</points>
<connection>
<GID>1570</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1119.5,180,-1119.5</points>
<connection>
<GID>6024</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1119.5,174,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1104,174,-1104</points>
<connection>
<GID>6022</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-65.5,116,-65.5</points>
<connection>
<GID>1573</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-65.5,110,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-50,110,-50</points>
<connection>
<GID>1572</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1119.5,205,-1119.5</points>
<connection>
<GID>6028</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1119.5,199,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1104,199,-1104</points>
<connection>
<GID>6026</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-65.5,139,-65.5</points>
<connection>
<GID>1575</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-65.5,133,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-50,133,-50</points>
<connection>
<GID>1574</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1119.5,228,-1119.5</points>
<connection>
<GID>6032</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1119.5,222,-1104</points>
<intersection>-1119.5 1</intersection>
<intersection>-1104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1104,222,-1104</points>
<connection>
<GID>6030</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-65.5,162,-65.5</points>
<connection>
<GID>1577</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-65.5,156,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-50,156,-50</points>
<connection>
<GID>1576</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1107,215,-1107</points>
<connection>
<GID>6030</GID>
<name>clock</name></connection>
<connection>
<GID>6026</GID>
<name>clock</name></connection>
<connection>
<GID>6022</GID>
<name>clock</name></connection>
<connection>
<GID>6018</GID>
<name>clock</name></connection>
<connection>
<GID>6014</GID>
<name>clock</name></connection>
<connection>
<GID>6010</GID>
<name>clock</name></connection>
<connection>
<GID>6006</GID>
<name>clock</name></connection>
<connection>
<GID>6002</GID>
<name>clock</name></connection>
<connection>
<GID>5998</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-65.5,185,-65.5</points>
<connection>
<GID>1579</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-65.5,179,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-50,179,-50</points>
<connection>
<GID>1578</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1116.5,226,-1116.5</points>
<connection>
<GID>6032</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6028</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6024</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6020</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6016</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6012</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6008</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6004</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6000</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-65.5,210,-65.5</points>
<connection>
<GID>1581</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-65.5,204,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-50,204,-50</points>
<connection>
<GID>1580</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1100.5,63,-1100.5</points>
<connection>
<GID>6040</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1100.5,57,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1085,57,-1085</points>
<connection>
<GID>6038</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-65.5,233,-65.5</points>
<connection>
<GID>1583</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-65.5,227,-50</points>
<intersection>-65.5 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-50,227,-50</points>
<connection>
<GID>1582</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1100.5,86,-1100.5</points>
<connection>
<GID>6044</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1100.5,80,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1085,80,-1085</points>
<connection>
<GID>6042</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-53,220,-53</points>
<connection>
<GID>1566</GID>
<name>OUT</name></connection>
<connection>
<GID>1568</GID>
<name>clock</name></connection>
<connection>
<GID>1570</GID>
<name>clock</name></connection>
<connection>
<GID>1572</GID>
<name>clock</name></connection>
<connection>
<GID>1574</GID>
<name>clock</name></connection>
<connection>
<GID>1576</GID>
<name>clock</name></connection>
<connection>
<GID>1578</GID>
<name>clock</name></connection>
<connection>
<GID>1580</GID>
<name>clock</name></connection>
<connection>
<GID>1582</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1100.5,111,-1100.5</points>
<connection>
<GID>6048</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1100.5,105,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1085,105,-1085</points>
<connection>
<GID>6046</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-62.5,231,-62.5</points>
<connection>
<GID>1569</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1571</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1573</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1575</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1577</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1579</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1581</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1583</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1567</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1100.5,134,-1100.5</points>
<connection>
<GID>6052</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1100.5,128,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1085,128,-1085</points>
<connection>
<GID>6050</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-47,68,-47</points>
<connection>
<GID>1587</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-47,62,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-31.5,62,-31.5</points>
<connection>
<GID>1586</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1100.5,157,-1100.5</points>
<connection>
<GID>6056</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1100.5,151,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1085,151,-1085</points>
<connection>
<GID>6054</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-47,91,-47</points>
<connection>
<GID>1589</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-47,85,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-31.5,85,-31.5</points>
<connection>
<GID>1588</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1100.5,180,-1100.5</points>
<connection>
<GID>6060</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1100.5,174,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1085,174,-1085</points>
<connection>
<GID>6058</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-47,116,-47</points>
<connection>
<GID>1591</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-47,110,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-31.5,110,-31.5</points>
<connection>
<GID>1590</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1100.5,205,-1100.5</points>
<connection>
<GID>6064</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1100.5,199,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1085,199,-1085</points>
<connection>
<GID>6062</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-47,139,-47</points>
<connection>
<GID>1593</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-47,133,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-31.5,133,-31.5</points>
<connection>
<GID>1592</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1100.5,228,-1100.5</points>
<connection>
<GID>6068</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1100.5,222,-1085</points>
<intersection>-1100.5 1</intersection>
<intersection>-1085 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1085,222,-1085</points>
<connection>
<GID>6066</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-47,162,-47</points>
<connection>
<GID>1595</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-47,156,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-31.5,156,-31.5</points>
<connection>
<GID>1594</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1088,215,-1088</points>
<connection>
<GID>6066</GID>
<name>clock</name></connection>
<connection>
<GID>6062</GID>
<name>clock</name></connection>
<connection>
<GID>6058</GID>
<name>clock</name></connection>
<connection>
<GID>6054</GID>
<name>clock</name></connection>
<connection>
<GID>6050</GID>
<name>clock</name></connection>
<connection>
<GID>6046</GID>
<name>clock</name></connection>
<connection>
<GID>6042</GID>
<name>clock</name></connection>
<connection>
<GID>6038</GID>
<name>clock</name></connection>
<connection>
<GID>6034</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-47,185,-47</points>
<connection>
<GID>1597</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-47,179,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-31.5,179,-31.5</points>
<connection>
<GID>1596</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1097.5,226,-1097.5</points>
<connection>
<GID>6068</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6064</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6060</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6056</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6052</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6048</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6044</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6040</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6036</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-47,210,-47</points>
<connection>
<GID>1599</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-47,204,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-31.5,204,-31.5</points>
<connection>
<GID>1598</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1082,63,-1082</points>
<connection>
<GID>6076</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1082,57,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1066.5,57,-1066.5</points>
<connection>
<GID>6074</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-47,233,-47</points>
<connection>
<GID>1601</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-47,227,-31.5</points>
<intersection>-47 1</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-31.5,227,-31.5</points>
<connection>
<GID>1600</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1082,86,-1082</points>
<connection>
<GID>6080</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1082,80,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1066.5,80,-1066.5</points>
<connection>
<GID>6078</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-34.5,220,-34.5</points>
<connection>
<GID>1584</GID>
<name>OUT</name></connection>
<connection>
<GID>1586</GID>
<name>clock</name></connection>
<connection>
<GID>1588</GID>
<name>clock</name></connection>
<connection>
<GID>1590</GID>
<name>clock</name></connection>
<connection>
<GID>1592</GID>
<name>clock</name></connection>
<connection>
<GID>1594</GID>
<name>clock</name></connection>
<connection>
<GID>1596</GID>
<name>clock</name></connection>
<connection>
<GID>1598</GID>
<name>clock</name></connection>
<connection>
<GID>1600</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1082,111,-1082</points>
<connection>
<GID>6084</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1082,105,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1066.5,105,-1066.5</points>
<connection>
<GID>6082</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-44,231,-44</points>
<connection>
<GID>1601</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1599</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1597</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1595</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1593</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1591</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1589</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1587</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1585</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1082,134,-1082</points>
<connection>
<GID>6088</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1082,128,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1066.5,128,-1066.5</points>
<connection>
<GID>6086</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-113,49.5,52</points>
<connection>
<GID>1603</GID>
<name>N_in0</name></connection>
<connection>
<GID>1635</GID>
<name>N_in1</name></connection>
<intersection>-87.5 12</intersection>
<intersection>-69 11</intersection>
<intersection>-50 10</intersection>
<intersection>-31.5 9</intersection>
<intersection>-9.5 8</intersection>
<intersection>9 7</intersection>
<intersection>28 6</intersection>
<intersection>46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,46.5,55,46.5</points>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>49.5,28,55,28</points>
<connection>
<GID>1496</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>49.5,9,55,9</points>
<connection>
<GID>1478</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>49.5,-9.5,55,-9.5</points>
<connection>
<GID>1442</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>49.5,-31.5,55,-31.5</points>
<connection>
<GID>1586</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>49.5,-50,55,-50</points>
<connection>
<GID>1568</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>49.5,-69,55,-69</points>
<connection>
<GID>1550</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>49.5,-87.5,55,-87.5</points>
<connection>
<GID>1532</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1082,157,-1082</points>
<connection>
<GID>6092</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1082,151,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1066.5,151,-1066.5</points>
<connection>
<GID>6090</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-112.5,72.5,52.5</points>
<connection>
<GID>1636</GID>
<name>N_in1</name></connection>
<connection>
<GID>1605</GID>
<name>N_in0</name></connection>
<intersection>-97.5 4</intersection>
<intersection>-79 5</intersection>
<intersection>-60 6</intersection>
<intersection>-41.5 7</intersection>
<intersection>-19.5 8</intersection>
<intersection>-1 9</intersection>
<intersection>18 10</intersection>
<intersection>36.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68,-97.5,72.5,-97.5</points>
<connection>
<GID>1533</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68,-79,72.5,-79</points>
<connection>
<GID>1551</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68,-60,72.5,-60</points>
<connection>
<GID>1569</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68,-41.5,72.5,-41.5</points>
<connection>
<GID>1587</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68,-19.5,72.5,-19.5</points>
<connection>
<GID>1447</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68,-1,72.5,-1</points>
<connection>
<GID>1479</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68,18,72.5,18</points>
<connection>
<GID>1497</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>68,36.5,72.5,36.5</points>
<connection>
<GID>1515</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1082,180,-1082</points>
<connection>
<GID>6096</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1082,174,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1066.5,174,-1066.5</points>
<connection>
<GID>6094</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-112.5,75.5,52</points>
<connection>
<GID>1606</GID>
<name>N_in0</name></connection>
<connection>
<GID>1637</GID>
<name>N_in1</name></connection>
<intersection>-87.5 10</intersection>
<intersection>-69 9</intersection>
<intersection>-50 8</intersection>
<intersection>-31.5 7</intersection>
<intersection>-9.5 6</intersection>
<intersection>9 5</intersection>
<intersection>28 4</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75.5,46.5,78,46.5</points>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>75.5,28,78,28</points>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>75.5,9,78,9</points>
<connection>
<GID>1480</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>75.5,-9.5,78,-9.5</points>
<connection>
<GID>1462</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>75.5,-31.5,78,-31.5</points>
<connection>
<GID>1588</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>75.5,-50,78,-50</points>
<connection>
<GID>1570</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>75.5,-69,78,-69</points>
<connection>
<GID>1552</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>75.5,-87.5,78,-87.5</points>
<connection>
<GID>1534</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1082,205,-1082</points>
<connection>
<GID>6100</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1082,199,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1066.5,199,-1066.5</points>
<connection>
<GID>6098</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-112.5,95,52.5</points>
<connection>
<GID>1607</GID>
<name>N_in0</name></connection>
<connection>
<GID>1638</GID>
<name>N_in1</name></connection>
<intersection>-97.5 6</intersection>
<intersection>-79 7</intersection>
<intersection>-60 8</intersection>
<intersection>-41.5 9</intersection>
<intersection>-19.5 10</intersection>
<intersection>-1 11</intersection>
<intersection>18 12</intersection>
<intersection>36.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91,-97.5,95,-97.5</points>
<connection>
<GID>1535</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>91,-79,95,-79</points>
<connection>
<GID>1553</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>91,-60,95,-60</points>
<connection>
<GID>1571</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>91,-41.5,95,-41.5</points>
<connection>
<GID>1589</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>91,-19.5,95,-19.5</points>
<connection>
<GID>1463</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>91,-1,95,-1</points>
<connection>
<GID>1481</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>91,18,95,18</points>
<connection>
<GID>1499</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>91,36.5,95,36.5</points>
<connection>
<GID>1517</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>4173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1082,228,-1082</points>
<connection>
<GID>6104</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1082,222,-1066.5</points>
<intersection>-1082 1</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1066.5,222,-1066.5</points>
<connection>
<GID>6102</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-112.5,98.5,52.5</points>
<connection>
<GID>1639</GID>
<name>N_in1</name></connection>
<connection>
<GID>1608</GID>
<name>N_in0</name></connection>
<intersection>-87.5 13</intersection>
<intersection>-69 12</intersection>
<intersection>-50 11</intersection>
<intersection>-31.5 10</intersection>
<intersection>-9.5 9</intersection>
<intersection>9 8</intersection>
<intersection>28 7</intersection>
<intersection>46.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>98.5,46.5,103,46.5</points>
<connection>
<GID>1518</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>98.5,28,103,28</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>98.5,9,103,9</points>
<connection>
<GID>1482</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>98.5,-9.5,103,-9.5</points>
<connection>
<GID>1464</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>98.5,-31.5,103,-31.5</points>
<connection>
<GID>1590</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>98.5,-50,103,-50</points>
<connection>
<GID>1572</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>98.5,-69,103,-69</points>
<connection>
<GID>1554</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>98.5,-87.5,103,-87.5</points>
<connection>
<GID>1536</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1069.5,215,-1069.5</points>
<connection>
<GID>6102</GID>
<name>clock</name></connection>
<connection>
<GID>6098</GID>
<name>clock</name></connection>
<connection>
<GID>6094</GID>
<name>clock</name></connection>
<connection>
<GID>6090</GID>
<name>clock</name></connection>
<connection>
<GID>6086</GID>
<name>clock</name></connection>
<connection>
<GID>6082</GID>
<name>clock</name></connection>
<connection>
<GID>6078</GID>
<name>clock</name></connection>
<connection>
<GID>6074</GID>
<name>clock</name></connection>
<connection>
<GID>6070</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-112.5,119.5,52</points>
<connection>
<GID>1609</GID>
<name>N_in0</name></connection>
<connection>
<GID>1640</GID>
<name>N_in1</name></connection>
<intersection>-97.5 6</intersection>
<intersection>-79 7</intersection>
<intersection>-60 8</intersection>
<intersection>-41.5 9</intersection>
<intersection>-19.5 10</intersection>
<intersection>-1 11</intersection>
<intersection>18 12</intersection>
<intersection>36.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116,-97.5,119.5,-97.5</points>
<connection>
<GID>1537</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116,-79,119.5,-79</points>
<connection>
<GID>1555</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>116,-60,119.5,-60</points>
<connection>
<GID>1573</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116,-41.5,119.5,-41.5</points>
<connection>
<GID>1591</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116,-19.5,119.5,-19.5</points>
<connection>
<GID>1465</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>116,-1,119.5,-1</points>
<connection>
<GID>1483</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>116,18,119.5,18</points>
<connection>
<GID>1501</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>116,36.5,119.5,36.5</points>
<connection>
<GID>1519</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1079,226,-1079</points>
<connection>
<GID>6104</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6100</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6096</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6092</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6088</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6084</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6080</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6076</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6072</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-112.5,123.5,52.5</points>
<connection>
<GID>1641</GID>
<name>N_in1</name></connection>
<connection>
<GID>1610</GID>
<name>N_in0</name></connection>
<intersection>-87.5 13</intersection>
<intersection>-69 12</intersection>
<intersection>-50 11</intersection>
<intersection>-31.5 10</intersection>
<intersection>-9.5 9</intersection>
<intersection>9 8</intersection>
<intersection>28 7</intersection>
<intersection>46.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>123.5,46.5,126,46.5</points>
<connection>
<GID>1520</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>123.5,28,126,28</points>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>123.5,9,126,9</points>
<connection>
<GID>1484</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>123.5,-9.5,126,-9.5</points>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>123.5,-31.5,126,-31.5</points>
<connection>
<GID>1592</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>123.5,-50,126,-50</points>
<connection>
<GID>1574</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>123.5,-69,126,-69</points>
<connection>
<GID>1556</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>123.5,-87.5,126,-87.5</points>
<connection>
<GID>1538</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1216,63,-1216</points>
<connection>
<GID>6112</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1216,57,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1200.5,57,-1200.5</points>
<connection>
<GID>6110</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-112.5,142,52.5</points>
<connection>
<GID>1611</GID>
<name>N_in0</name></connection>
<connection>
<GID>1642</GID>
<name>N_in1</name></connection>
<intersection>-97.5 6</intersection>
<intersection>-79 7</intersection>
<intersection>-60 8</intersection>
<intersection>-41.5 9</intersection>
<intersection>-19.5 10</intersection>
<intersection>-1 11</intersection>
<intersection>18 12</intersection>
<intersection>36.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-97.5,142,-97.5</points>
<connection>
<GID>1539</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,-79,142,-79</points>
<connection>
<GID>1557</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>139,-60,142,-60</points>
<connection>
<GID>1575</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>139,-41.5,142,-41.5</points>
<connection>
<GID>1593</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>139,-19.5,142,-19.5</points>
<connection>
<GID>1467</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139,-1,142,-1</points>
<connection>
<GID>1485</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>139,18,142,18</points>
<connection>
<GID>1503</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>139,36.5,142,36.5</points>
<connection>
<GID>1521</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>4177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1216,86,-1216</points>
<connection>
<GID>6116</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1216,80,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1200.5,80,-1200.5</points>
<connection>
<GID>6114</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-112.5,146,52.5</points>
<connection>
<GID>1643</GID>
<name>N_in1</name></connection>
<connection>
<GID>1612</GID>
<name>N_in0</name></connection>
<intersection>-87.5 13</intersection>
<intersection>-69 12</intersection>
<intersection>-50 11</intersection>
<intersection>-31.5 10</intersection>
<intersection>-9.5 9</intersection>
<intersection>9 8</intersection>
<intersection>28 7</intersection>
<intersection>46.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>146,46.5,149,46.5</points>
<connection>
<GID>1522</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>146,28,149,28</points>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>146,9,149,9</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>146,-9.5,149,-9.5</points>
<connection>
<GID>1468</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>146,-31.5,149,-31.5</points>
<connection>
<GID>1594</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>146,-50,149,-50</points>
<connection>
<GID>1576</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>146,-69,149,-69</points>
<connection>
<GID>1558</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>146,-87.5,149,-87.5</points>
<connection>
<GID>1540</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment></shape></wire>
<wire>
<ID>4178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1216,111,-1216</points>
<connection>
<GID>6120</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1216,105,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1200.5,105,-1200.5</points>
<connection>
<GID>6118</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-112,165,52.5</points>
<connection>
<GID>1613</GID>
<name>N_in0</name></connection>
<connection>
<GID>1644</GID>
<name>N_in1</name></connection>
<intersection>-97.5 6</intersection>
<intersection>-79 7</intersection>
<intersection>-60 8</intersection>
<intersection>-41.5 9</intersection>
<intersection>-19.5 10</intersection>
<intersection>-1 11</intersection>
<intersection>18 12</intersection>
<intersection>36.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>162,-97.5,165,-97.5</points>
<connection>
<GID>1541</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162,-79,165,-79</points>
<connection>
<GID>1559</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>162,-60,165,-60</points>
<connection>
<GID>1577</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162,-41.5,165,-41.5</points>
<connection>
<GID>1595</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>162,-19.5,165,-19.5</points>
<connection>
<GID>1469</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>162,-1,165,-1</points>
<connection>
<GID>1487</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>162,18,165,18</points>
<connection>
<GID>1505</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>162,36.5,165,36.5</points>
<connection>
<GID>1523</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>4179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1216,134,-1216</points>
<connection>
<GID>5761</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1216,128,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1200.5,128,-1200.5</points>
<connection>
<GID>5759</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-112,170,52.5</points>
<connection>
<GID>1645</GID>
<name>N_in1</name></connection>
<connection>
<GID>1614</GID>
<name>N_in0</name></connection>
<intersection>-87.5 13</intersection>
<intersection>-69 12</intersection>
<intersection>-50 11</intersection>
<intersection>-31.5 10</intersection>
<intersection>-9.5 9</intersection>
<intersection>9 8</intersection>
<intersection>28 7</intersection>
<intersection>46.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>170,46.5,172,46.5</points>
<connection>
<GID>1524</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>170,28,172,28</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>170,9,172,9</points>
<connection>
<GID>1488</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>170,-9.5,172,-9.5</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>170,-31.5,172,-31.5</points>
<connection>
<GID>1596</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>170,-50,172,-50</points>
<connection>
<GID>1578</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>170,-69,172,-69</points>
<connection>
<GID>1560</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>170,-87.5,172,-87.5</points>
<connection>
<GID>1542</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>4180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1216,157,-1216</points>
<connection>
<GID>5765</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1216,151,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1200.5,151,-1200.5</points>
<connection>
<GID>5763</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-111.5,188,52.5</points>
<connection>
<GID>1616</GID>
<name>N_in0</name></connection>
<connection>
<GID>1646</GID>
<name>N_in1</name></connection>
<intersection>-97.5 16</intersection>
<intersection>-79 15</intersection>
<intersection>-60 14</intersection>
<intersection>-41.5 13</intersection>
<intersection>-19.5 12</intersection>
<intersection>-1 11</intersection>
<intersection>18 10</intersection>
<intersection>36.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>185,36.5,188,36.5</points>
<connection>
<GID>1525</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>185,18,188,18</points>
<connection>
<GID>1507</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>185,-1,188,-1</points>
<connection>
<GID>1489</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185,-19.5,188,-19.5</points>
<connection>
<GID>1471</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>185,-41.5,188,-41.5</points>
<connection>
<GID>1597</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>185,-60,188,-60</points>
<connection>
<GID>1579</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>185,-79,188,-79</points>
<connection>
<GID>1561</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>185,-97.5,188,-97.5</points>
<connection>
<GID>1543</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment></shape></wire>
<wire>
<ID>4181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1216,180,-1216</points>
<connection>
<GID>5769</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1216,174,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1200.5,174,-1200.5</points>
<connection>
<GID>5767</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-111.5,192.5,52.5</points>
<connection>
<GID>1647</GID>
<name>N_in1</name></connection>
<connection>
<GID>1615</GID>
<name>N_in0</name></connection>
<intersection>-87.5 13</intersection>
<intersection>-69 12</intersection>
<intersection>-50 11</intersection>
<intersection>-31.5 10</intersection>
<intersection>-9.5 9</intersection>
<intersection>9 8</intersection>
<intersection>28 7</intersection>
<intersection>46.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>192.5,46.5,197,46.5</points>
<connection>
<GID>1526</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>192.5,28,197,28</points>
<connection>
<GID>1508</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>192.5,9,197,9</points>
<connection>
<GID>1490</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>192.5,-9.5,197,-9.5</points>
<connection>
<GID>1472</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>192.5,-31.5,197,-31.5</points>
<connection>
<GID>1598</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>192.5,-50,197,-50</points>
<connection>
<GID>1580</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>192.5,-69,197,-69</points>
<connection>
<GID>1562</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>192.5,-87.5,197,-87.5</points>
<connection>
<GID>1544</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1216,205,-1216</points>
<connection>
<GID>5773</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1216,199,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1200.5,199,-1200.5</points>
<connection>
<GID>5771</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-111,213.5,52</points>
<connection>
<GID>1648</GID>
<name>N_in1</name></connection>
<connection>
<GID>1617</GID>
<name>N_in0</name></connection>
<intersection>-97.5 6</intersection>
<intersection>-79 7</intersection>
<intersection>-60 8</intersection>
<intersection>-41.5 9</intersection>
<intersection>-19.5 10</intersection>
<intersection>-1 11</intersection>
<intersection>18 12</intersection>
<intersection>36.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>210,-97.5,213.5,-97.5</points>
<connection>
<GID>1545</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>210,-79,213.5,-79</points>
<connection>
<GID>1563</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>210,-60,213.5,-60</points>
<connection>
<GID>1581</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>210,-41.5,213.5,-41.5</points>
<connection>
<GID>1599</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210,-19.5,213.5,-19.5</points>
<connection>
<GID>1473</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>210,-1,213.5,-1</points>
<connection>
<GID>1491</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>210,18,213.5,18</points>
<connection>
<GID>1509</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>210,36.5,213.5,36.5</points>
<connection>
<GID>1527</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1216,228,-1216</points>
<connection>
<GID>5777</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1216,222,-1200.5</points>
<intersection>-1216 1</intersection>
<intersection>-1200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1200.5,222,-1200.5</points>
<connection>
<GID>5775</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-111,217,52</points>
<connection>
<GID>1651</GID>
<name>N_in0</name></connection>
<connection>
<GID>1649</GID>
<name>N_in1</name></connection>
<intersection>-87.5 11</intersection>
<intersection>-69 10</intersection>
<intersection>-50 9</intersection>
<intersection>-31.5 7</intersection>
<intersection>-9.5 6</intersection>
<intersection>9 5</intersection>
<intersection>28 4</intersection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,46.5,220,46.5</points>
<connection>
<GID>1528</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>217,28,220,28</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>217,9,220,9</points>
<connection>
<GID>1492</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>217,-9.5,220,-9.5</points>
<connection>
<GID>1474</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>217,-31.5,220,-31.5</points>
<connection>
<GID>1600</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>217,-50,220,-50</points>
<connection>
<GID>1582</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>217,-69,220,-69</points>
<connection>
<GID>1564</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>217,-87.5,220,-87.5</points>
<connection>
<GID>1546</GID>
<name>IN_0</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>4184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1203.5,215,-1203.5</points>
<connection>
<GID>6118</GID>
<name>clock</name></connection>
<connection>
<GID>6114</GID>
<name>clock</name></connection>
<connection>
<GID>6110</GID>
<name>clock</name></connection>
<connection>
<GID>6106</GID>
<name>OUT</name></connection>
<connection>
<GID>5775</GID>
<name>clock</name></connection>
<connection>
<GID>5771</GID>
<name>clock</name></connection>
<connection>
<GID>5767</GID>
<name>clock</name></connection>
<connection>
<GID>5763</GID>
<name>clock</name></connection>
<connection>
<GID>5759</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-111,238,51</points>
<connection>
<GID>1653</GID>
<name>N_in1</name></connection>
<connection>
<GID>1618</GID>
<name>N_in0</name></connection>
<intersection>-97.5 11</intersection>
<intersection>-79 10</intersection>
<intersection>-60 9</intersection>
<intersection>-41.5 8</intersection>
<intersection>-19.5 7</intersection>
<intersection>-1 6</intersection>
<intersection>18 5</intersection>
<intersection>36.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>233,36.5,238,36.5</points>
<connection>
<GID>1529</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>233,18,238,18</points>
<connection>
<GID>1511</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>233,-1,238,-1</points>
<connection>
<GID>1493</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>233,-19.5,238,-19.5</points>
<connection>
<GID>1475</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>233,-41.5,238,-41.5</points>
<connection>
<GID>1601</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>233,-60,238,-60</points>
<connection>
<GID>1583</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>233,-79,238,-79</points>
<connection>
<GID>1565</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>233,-97.5,238,-97.5</points>
<connection>
<GID>1547</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>4185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1213,226,-1213</points>
<connection>
<GID>6120</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6116</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6112</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6108</GID>
<name>OUT</name></connection>
<connection>
<GID>5777</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5773</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5769</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5765</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5761</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-119,44.5,27.5,44.5</points>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-107,-119,44.5</points>
<connection>
<GID>1664</GID>
<name>OUT_15</name></connection>
<intersection>35 4</intersection>
<intersection>44.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,35,39,35</points>
<connection>
<GID>1513</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>4186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1197.5,63,-1197.5</points>
<connection>
<GID>5785</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1197.5,57,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1182,57,-1182</points>
<connection>
<GID>5783</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-118,26,27.5,26</points>
<connection>
<GID>1494</GID>
<name>IN_0</name></connection>
<intersection>-118 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-118,-108,-118,26</points>
<intersection>-108 6</intersection>
<intersection>16.5 5</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-118,16.5,39,16.5</points>
<connection>
<GID>1495</GID>
<name>IN_0</name></connection>
<intersection>-118 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119,-108,-118,-108</points>
<connection>
<GID>1664</GID>
<name>OUT_14</name></connection>
<intersection>-118 4</intersection></hsegment></shape></wire>
<wire>
<ID>4187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1197.5,86,-1197.5</points>
<connection>
<GID>5789</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1197.5,80,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1182,80,-1182</points>
<connection>
<GID>5787</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-117,7,27.5,7</points>
<connection>
<GID>1476</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-109,-117,7</points>
<intersection>-109 6</intersection>
<intersection>-2.5 4</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-2.5,39,-2.5</points>
<connection>
<GID>1477</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119,-109,-117,-109</points>
<connection>
<GID>1664</GID>
<name>OUT_13</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>4188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1197.5,111,-1197.5</points>
<connection>
<GID>5793</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1197.5,105,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1182,105,-1182</points>
<connection>
<GID>5791</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-116,-11.5,27.5,-11.5</points>
<connection>
<GID>1434</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-116,-110,-116,-11.5</points>
<intersection>-110 5</intersection>
<intersection>-21 4</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-116,-21,39,-21</points>
<connection>
<GID>1438</GID>
<name>IN_0</name></connection>
<intersection>-116 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-110,-116,-110</points>
<connection>
<GID>1664</GID>
<name>OUT_12</name></connection>
<intersection>-116 3</intersection></hsegment></shape></wire>
<wire>
<ID>4189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1197.5,134,-1197.5</points>
<connection>
<GID>5797</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1197.5,128,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1182,128,-1182</points>
<connection>
<GID>5795</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1197.5,157,-1197.5</points>
<connection>
<GID>5801</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1197.5,151,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1182,151,-1182</points>
<connection>
<GID>5799</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115,-33.5,27.5,-33.5</points>
<connection>
<GID>1584</GID>
<name>IN_0</name></connection>
<intersection>-115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-115,-111,-115,-33.5</points>
<intersection>-111 6</intersection>
<intersection>-43 4</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-115,-43,38.5,-43</points>
<connection>
<GID>1585</GID>
<name>IN_0</name></connection>
<intersection>-115 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119,-111,-115,-111</points>
<connection>
<GID>1664</GID>
<name>OUT_11</name></connection>
<intersection>-115 3</intersection></hsegment></shape></wire>
<wire>
<ID>4191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1197.5,180,-1197.5</points>
<connection>
<GID>5805</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1197.5,174,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1182,174,-1182</points>
<connection>
<GID>5803</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-52,27.5,-52</points>
<connection>
<GID>1566</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114,-112,-114,-52</points>
<intersection>-112 5</intersection>
<intersection>-61.5 4</intersection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-114,-61.5,38.5,-61.5</points>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection>
<intersection>-114 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-112,-114,-112</points>
<connection>
<GID>1664</GID>
<name>OUT_10</name></connection>
<intersection>-114 3</intersection></hsegment></shape></wire>
<wire>
<ID>4192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1197.5,205,-1197.5</points>
<connection>
<GID>5809</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1197.5,199,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1182,199,-1182</points>
<connection>
<GID>5807</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,-71,27.5,-71</points>
<connection>
<GID>1548</GID>
<name>IN_0</name></connection>
<intersection>-113 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-113,-113,-113,-71</points>
<intersection>-113 5</intersection>
<intersection>-80.5 4</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-113,-80.5,38.5,-80.5</points>
<connection>
<GID>1549</GID>
<name>IN_0</name></connection>
<intersection>-113 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-113,-113,-113</points>
<connection>
<GID>1664</GID>
<name>OUT_9</name></connection>
<intersection>-113 3</intersection></hsegment></shape></wire>
<wire>
<ID>4193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1197.5,228,-1197.5</points>
<connection>
<GID>5813</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1197.5,222,-1182</points>
<intersection>-1197.5 1</intersection>
<intersection>-1182 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1182,222,-1182</points>
<connection>
<GID>5811</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-112,-89.5,27.5,-89.5</points>
<connection>
<GID>1530</GID>
<name>IN_0</name></connection>
<intersection>-112 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-112,-114,-112,-89.5</points>
<intersection>-114 5</intersection>
<intersection>-99 4</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-112,-99,38.5,-99</points>
<connection>
<GID>1531</GID>
<name>IN_0</name></connection>
<intersection>-112 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119,-114,-112,-114</points>
<connection>
<GID>1664</GID>
<name>OUT_8</name></connection>
<intersection>-112 3</intersection></hsegment></shape></wire>
<wire>
<ID>4194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1185,215,-1185</points>
<connection>
<GID>5811</GID>
<name>clock</name></connection>
<connection>
<GID>5807</GID>
<name>clock</name></connection>
<connection>
<GID>5803</GID>
<name>clock</name></connection>
<connection>
<GID>5799</GID>
<name>clock</name></connection>
<connection>
<GID>5795</GID>
<name>clock</name></connection>
<connection>
<GID>5791</GID>
<name>clock</name></connection>
<connection>
<GID>5787</GID>
<name>clock</name></connection>
<connection>
<GID>5783</GID>
<name>clock</name></connection>
<connection>
<GID>5779</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1194.5,226,-1194.5</points>
<connection>
<GID>5813</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5809</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5805</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5801</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5797</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5793</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5789</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5785</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5781</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1178.5,63,-1178.5</points>
<connection>
<GID>5823</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1178.5,57,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1163,57,-1163</points>
<connection>
<GID>5821</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-113,26.5,52</points>
<connection>
<GID>1658</GID>
<name>N_in0</name></connection>
<connection>
<GID>1660</GID>
<name>N_in1</name></connection>
<intersection>-91.5 10</intersection>
<intersection>-73 9</intersection>
<intersection>-54 8</intersection>
<intersection>-35.5 7</intersection>
<intersection>-13.5 6</intersection>
<intersection>5 5</intersection>
<intersection>24 4</intersection>
<intersection>42.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,42.5,27.5,42.5</points>
<connection>
<GID>1512</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26.5,24,27.5,24</points>
<connection>
<GID>1494</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26.5,5,27.5,5</points>
<connection>
<GID>1476</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>26.5,-13.5,27.5,-13.5</points>
<connection>
<GID>1434</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>26.5,-35.5,27.5,-35.5</points>
<connection>
<GID>1584</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>26.5,-54,27.5,-54</points>
<connection>
<GID>1566</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>26.5,-73,27.5,-73</points>
<connection>
<GID>1548</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>26.5,-91.5,27.5,-91.5</points>
<connection>
<GID>1530</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1178.5,86,-1178.5</points>
<connection>
<GID>5828</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1178.5,80,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1163,80,-1163</points>
<connection>
<GID>5826</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-113,36.5,52</points>
<connection>
<GID>1657</GID>
<name>N_in0</name></connection>
<connection>
<GID>1659</GID>
<name>N_in1</name></connection>
<intersection>-101 3</intersection>
<intersection>-82.5 5</intersection>
<intersection>-63.5 7</intersection>
<intersection>-45 9</intersection>
<intersection>-23 11</intersection>
<intersection>-4.5 13</intersection>
<intersection>14.5 15</intersection>
<intersection>33 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-101,38.5,-101</points>
<connection>
<GID>1531</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>36.5,-82.5,38.5,-82.5</points>
<connection>
<GID>1549</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>36.5,-63.5,38.5,-63.5</points>
<connection>
<GID>1567</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>36.5,-45,38.5,-45</points>
<connection>
<GID>1585</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>36.5,-23,39,-23</points>
<connection>
<GID>1438</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>36.5,-4.5,39,-4.5</points>
<connection>
<GID>1477</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>36.5,14.5,39,14.5</points>
<connection>
<GID>1495</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>36.5,33,39,33</points>
<connection>
<GID>1513</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1178.5,111,-1178.5</points>
<connection>
<GID>5833</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1178.5,105,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1163,105,-1163</points>
<connection>
<GID>5831</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-200.5,68,-200.5</points>
<connection>
<GID>4202</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-200.5,62,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-185,62,-185</points>
<connection>
<GID>4196</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1178.5,134,-1178.5</points>
<connection>
<GID>5838</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1178.5,128,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1163,128,-1163</points>
<connection>
<GID>5836</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-200.5,91,-200.5</points>
<connection>
<GID>4215</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-200.5,85,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-185,85,-185</points>
<connection>
<GID>4214</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1178.5,157,-1178.5</points>
<connection>
<GID>5843</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1178.5,151,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1163,151,-1163</points>
<connection>
<GID>5841</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-200.5,116,-200.5</points>
<connection>
<GID>4219</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-200.5,110,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-185,110,-185</points>
<connection>
<GID>4217</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1178.5,180,-1178.5</points>
<connection>
<GID>5846</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1178.5,174,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1163,174,-1163</points>
<connection>
<GID>5845</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-200.5,139,-200.5</points>
<connection>
<GID>4223</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-200.5,133,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-185,133,-185</points>
<connection>
<GID>4221</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1178.5,205,-1178.5</points>
<connection>
<GID>5849</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1178.5,199,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1163,199,-1163</points>
<connection>
<GID>5848</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-200.5,162,-200.5</points>
<connection>
<GID>4226</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-200.5,156,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-185,156,-185</points>
<connection>
<GID>4224</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1178.5,228,-1178.5</points>
<connection>
<GID>5851</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1178.5,222,-1163</points>
<intersection>-1178.5 1</intersection>
<intersection>-1163 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1163,222,-1163</points>
<connection>
<GID>5850</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-200.5,185,-200.5</points>
<connection>
<GID>4228</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-200.5,179,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-185,179,-185</points>
<connection>
<GID>4227</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1166,215,-1166</points>
<connection>
<GID>5850</GID>
<name>clock</name></connection>
<connection>
<GID>5848</GID>
<name>clock</name></connection>
<connection>
<GID>5845</GID>
<name>clock</name></connection>
<connection>
<GID>5841</GID>
<name>clock</name></connection>
<connection>
<GID>5836</GID>
<name>clock</name></connection>
<connection>
<GID>5831</GID>
<name>clock</name></connection>
<connection>
<GID>5826</GID>
<name>clock</name></connection>
<connection>
<GID>5821</GID>
<name>clock</name></connection>
<connection>
<GID>5816</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-200.5,210,-200.5</points>
<connection>
<GID>4230</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-200.5,204,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-185,204,-185</points>
<connection>
<GID>4229</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1175.5,226,-1175.5</points>
<connection>
<GID>5851</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5849</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5846</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5843</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5838</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5833</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5828</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5823</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5818</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-200.5,233,-200.5</points>
<connection>
<GID>4232</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-200.5,227,-185</points>
<intersection>-200.5 1</intersection>
<intersection>-185 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-185,227,-185</points>
<connection>
<GID>4231</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1160,63,-1160</points>
<connection>
<GID>5855</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1160,57,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1144.5,57,-1144.5</points>
<connection>
<GID>5854</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-188,220,-188</points>
<connection>
<GID>4231</GID>
<name>clock</name></connection>
<connection>
<GID>4229</GID>
<name>clock</name></connection>
<connection>
<GID>4227</GID>
<name>clock</name></connection>
<connection>
<GID>4224</GID>
<name>clock</name></connection>
<connection>
<GID>4221</GID>
<name>clock</name></connection>
<connection>
<GID>4217</GID>
<name>clock</name></connection>
<connection>
<GID>4214</GID>
<name>clock</name></connection>
<connection>
<GID>4196</GID>
<name>clock</name></connection>
<connection>
<GID>4193</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1160,86,-1160</points>
<connection>
<GID>5857</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1160,80,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1144.5,80,-1144.5</points>
<connection>
<GID>5856</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-197.5,231,-197.5</points>
<connection>
<GID>4232</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4230</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4228</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4226</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4223</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4219</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4215</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4202</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4194</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1160,111,-1160</points>
<connection>
<GID>5859</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1160,105,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1144.5,105,-1144.5</points>
<connection>
<GID>5858</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-182,68,-182</points>
<connection>
<GID>4236</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-182,62,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-166.5,62,-166.5</points>
<connection>
<GID>4235</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1160,134,-1160</points>
<connection>
<GID>5861</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1160,128,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1144.5,128,-1144.5</points>
<connection>
<GID>5860</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-182,91,-182</points>
<connection>
<GID>4238</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-182,85,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-166.5,85,-166.5</points>
<connection>
<GID>4237</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1160,157,-1160</points>
<connection>
<GID>5863</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1160,151,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1144.5,151,-1144.5</points>
<connection>
<GID>5862</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-182,116,-182</points>
<connection>
<GID>4240</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-182,110,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-166.5,110,-166.5</points>
<connection>
<GID>4239</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1160,180,-1160</points>
<connection>
<GID>5865</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1160,174,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1144.5,174,-1144.5</points>
<connection>
<GID>5864</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-182,139,-182</points>
<connection>
<GID>4242</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-182,133,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-166.5,133,-166.5</points>
<connection>
<GID>4241</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1160,205,-1160</points>
<connection>
<GID>5867</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1160,199,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1144.5,199,-1144.5</points>
<connection>
<GID>5866</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-182,162,-182</points>
<connection>
<GID>4244</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-182,156,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-166.5,156,-166.5</points>
<connection>
<GID>4243</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1160,228,-1160</points>
<connection>
<GID>5869</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1160,222,-1144.5</points>
<intersection>-1160 1</intersection>
<intersection>-1144.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1144.5,222,-1144.5</points>
<connection>
<GID>5868</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-182,185,-182</points>
<connection>
<GID>4246</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-182,179,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-166.5,179,-166.5</points>
<connection>
<GID>4245</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1147.5,215,-1147.5</points>
<connection>
<GID>5868</GID>
<name>clock</name></connection>
<connection>
<GID>5866</GID>
<name>clock</name></connection>
<connection>
<GID>5864</GID>
<name>clock</name></connection>
<connection>
<GID>5862</GID>
<name>clock</name></connection>
<connection>
<GID>5860</GID>
<name>clock</name></connection>
<connection>
<GID>5858</GID>
<name>clock</name></connection>
<connection>
<GID>5856</GID>
<name>clock</name></connection>
<connection>
<GID>5854</GID>
<name>clock</name></connection>
<connection>
<GID>5852</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-182,210,-182</points>
<connection>
<GID>4248</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-182,204,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-166.5,204,-166.5</points>
<connection>
<GID>4247</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1157,226,-1157</points>
<connection>
<GID>5869</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5867</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5865</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5863</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5861</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5859</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5857</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5855</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5853</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-182,233,-182</points>
<connection>
<GID>4250</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-182,227,-166.5</points>
<intersection>-182 1</intersection>
<intersection>-166.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-166.5,227,-166.5</points>
<connection>
<GID>4249</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-1226,44.5,-1061</points>
<connection>
<GID>5885</GID>
<name>N_in1</name></connection>
<connection>
<GID>5870</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 12</intersection>
<intersection>-1182 11</intersection>
<intersection>-1163 10</intersection>
<intersection>-1144.5 9</intersection>
<intersection>-1122.5 8</intersection>
<intersection>-1104 7</intersection>
<intersection>-1085 6</intersection>
<intersection>-1066.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-1066.5,50,-1066.5</points>
<connection>
<GID>6074</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>44.5,-1085,50,-1085</points>
<connection>
<GID>6038</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-1104,50,-1104</points>
<connection>
<GID>6002</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>44.5,-1122.5,50,-1122.5</points>
<connection>
<GID>5948</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>44.5,-1144.5,50,-1144.5</points>
<connection>
<GID>5854</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>44.5,-1163,50,-1163</points>
<connection>
<GID>5821</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>44.5,-1182,50,-1182</points>
<connection>
<GID>5783</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>44.5,-1200.5,50,-1200.5</points>
<connection>
<GID>6110</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-169.5,220,-169.5</points>
<connection>
<GID>4249</GID>
<name>clock</name></connection>
<connection>
<GID>4247</GID>
<name>clock</name></connection>
<connection>
<GID>4245</GID>
<name>clock</name></connection>
<connection>
<GID>4243</GID>
<name>clock</name></connection>
<connection>
<GID>4241</GID>
<name>clock</name></connection>
<connection>
<GID>4239</GID>
<name>clock</name></connection>
<connection>
<GID>4237</GID>
<name>clock</name></connection>
<connection>
<GID>4235</GID>
<name>clock</name></connection>
<connection>
<GID>4233</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-1225.5,67.5,-1060.5</points>
<connection>
<GID>5886</GID>
<name>N_in1</name></connection>
<connection>
<GID>5871</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 4</intersection>
<intersection>-1190 5</intersection>
<intersection>-1171 6</intersection>
<intersection>-1152.5 7</intersection>
<intersection>-1130.5 8</intersection>
<intersection>-1112 9</intersection>
<intersection>-1093 10</intersection>
<intersection>-1074.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63,-1208.5,67.5,-1208.5</points>
<intersection>63 12</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-1190,67.5,-1190</points>
<intersection>63 13</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>63,-1171,67.5,-1171</points>
<intersection>63 14</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>63,-1152.5,67.5,-1152.5</points>
<intersection>63 15</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>63,-1130.5,67.5,-1130.5</points>
<intersection>63 18</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-1112,67.5,-1112</points>
<intersection>63 19</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>63,-1093,67.5,-1093</points>
<intersection>63 20</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>63,-1074.5,67.5,-1074.5</points>
<intersection>63 21</intersection>
<intersection>67.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>63,-1210.5,63,-1208.5</points>
<connection>
<GID>6112</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>63,-1192,63,-1190</points>
<connection>
<GID>5785</GID>
<name>OUT_0</name></connection>
<intersection>-1190 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>63,-1173,63,-1171</points>
<connection>
<GID>5823</GID>
<name>OUT_0</name></connection>
<intersection>-1171 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>63,-1154.5,63,-1152.5</points>
<connection>
<GID>5855</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>63,-1132.5,63,-1130.5</points>
<connection>
<GID>5954</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>63,-1114,63,-1112</points>
<connection>
<GID>6004</GID>
<name>OUT_0</name></connection>
<intersection>-1112 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>63,-1095,63,-1093</points>
<connection>
<GID>6040</GID>
<name>OUT_0</name></connection>
<intersection>-1093 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>63,-1076.5,63,-1074.5</points>
<connection>
<GID>6076</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-179,231,-179</points>
<connection>
<GID>4250</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4248</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4246</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4244</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4242</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4240</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4238</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4236</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4234</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-1225.5,70.5,-1061</points>
<connection>
<GID>5887</GID>
<name>N_in1</name></connection>
<connection>
<GID>5872</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 10</intersection>
<intersection>-1182 9</intersection>
<intersection>-1163 8</intersection>
<intersection>-1144.5 7</intersection>
<intersection>-1122.5 6</intersection>
<intersection>-1104 5</intersection>
<intersection>-1085 4</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70.5,-1066.5,73,-1066.5</points>
<connection>
<GID>6078</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-1085,73,-1085</points>
<connection>
<GID>6042</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-1104,73,-1104</points>
<connection>
<GID>6006</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>70.5,-1122.5,73,-1122.5</points>
<connection>
<GID>5970</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>70.5,-1144.5,73,-1144.5</points>
<connection>
<GID>5856</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>70.5,-1163,73,-1163</points>
<connection>
<GID>5826</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>70.5,-1182,73,-1182</points>
<connection>
<GID>5787</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>70.5,-1200.5,73,-1200.5</points>
<connection>
<GID>6114</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-163,68,-163</points>
<connection>
<GID>4254</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-163,62,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-147.5,62,-147.5</points>
<connection>
<GID>4253</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-1225.5,90,-1060.5</points>
<connection>
<GID>5888</GID>
<name>N_in1</name></connection>
<connection>
<GID>5873</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 6</intersection>
<intersection>-1190 7</intersection>
<intersection>-1171 8</intersection>
<intersection>-1152.5 9</intersection>
<intersection>-1130.5 10</intersection>
<intersection>-1112 11</intersection>
<intersection>-1093 12</intersection>
<intersection>-1074.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-1208.5,90,-1208.5</points>
<intersection>86 14</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>86,-1190,90,-1190</points>
<intersection>86 15</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>86,-1171,90,-1171</points>
<intersection>86 16</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>86,-1152.5,90,-1152.5</points>
<intersection>86 17</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>86,-1130.5,90,-1130.5</points>
<intersection>86 20</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>86,-1112,90,-1112</points>
<intersection>86 21</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>86,-1093,90,-1093</points>
<intersection>86 22</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>86,-1074.5,90,-1074.5</points>
<intersection>86 23</intersection>
<intersection>90 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>86,-1210.5,86,-1208.5</points>
<connection>
<GID>6116</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>86,-1192,86,-1190</points>
<connection>
<GID>5789</GID>
<name>OUT_0</name></connection>
<intersection>-1190 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>86,-1173,86,-1171</points>
<connection>
<GID>5828</GID>
<name>OUT_0</name></connection>
<intersection>-1171 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>86,-1154.5,86,-1152.5</points>
<connection>
<GID>5857</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>86,-1132.5,86,-1130.5</points>
<connection>
<GID>5972</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>86,-1114,86,-1112</points>
<connection>
<GID>6008</GID>
<name>OUT_0</name></connection>
<intersection>-1112 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>86,-1095,86,-1093</points>
<connection>
<GID>6044</GID>
<name>OUT_0</name></connection>
<intersection>-1093 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>86,-1076.5,86,-1074.5</points>
<connection>
<GID>6080</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-163,91,-163</points>
<connection>
<GID>4256</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-163,85,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-147.5,85,-147.5</points>
<connection>
<GID>4255</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-1225.5,93.5,-1060.5</points>
<connection>
<GID>5889</GID>
<name>N_in1</name></connection>
<connection>
<GID>5874</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 13</intersection>
<intersection>-1182 12</intersection>
<intersection>-1163 11</intersection>
<intersection>-1144.5 10</intersection>
<intersection>-1122.5 9</intersection>
<intersection>-1104 8</intersection>
<intersection>-1085 7</intersection>
<intersection>-1066.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>93.5,-1066.5,98,-1066.5</points>
<connection>
<GID>6082</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>93.5,-1085,98,-1085</points>
<connection>
<GID>6046</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>93.5,-1104,98,-1104</points>
<connection>
<GID>6010</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-1122.5,98,-1122.5</points>
<connection>
<GID>5974</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>93.5,-1144.5,98,-1144.5</points>
<connection>
<GID>5858</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>93.5,-1163,98,-1163</points>
<connection>
<GID>5831</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>93.5,-1182,98,-1182</points>
<connection>
<GID>5791</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>93.5,-1200.5,98,-1200.5</points>
<connection>
<GID>6118</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-163,116,-163</points>
<connection>
<GID>4258</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-163,110,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-147.5,110,-147.5</points>
<connection>
<GID>4257</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-1225.5,114.5,-1061</points>
<connection>
<GID>5890</GID>
<name>N_in1</name></connection>
<connection>
<GID>5875</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 6</intersection>
<intersection>-1190 7</intersection>
<intersection>-1171 8</intersection>
<intersection>-1152.5 9</intersection>
<intersection>-1130.5 10</intersection>
<intersection>-1112 11</intersection>
<intersection>-1093 12</intersection>
<intersection>-1074.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>111,-1208.5,114.5,-1208.5</points>
<intersection>111 14</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111,-1190,114.5,-1190</points>
<intersection>111 15</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111,-1171,114.5,-1171</points>
<intersection>111 16</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111,-1152.5,114.5,-1152.5</points>
<intersection>111 17</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,-1130.5,114.5,-1130.5</points>
<intersection>111 20</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>111,-1112,114.5,-1112</points>
<intersection>111 21</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>111,-1093,114.5,-1093</points>
<intersection>111 22</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111,-1074.5,114.5,-1074.5</points>
<intersection>111 23</intersection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>111,-1210.5,111,-1208.5</points>
<connection>
<GID>6120</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>111,-1192,111,-1190</points>
<connection>
<GID>5793</GID>
<name>OUT_0</name></connection>
<intersection>-1190 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>111,-1173,111,-1171</points>
<connection>
<GID>5833</GID>
<name>OUT_0</name></connection>
<intersection>-1171 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>111,-1154.5,111,-1152.5</points>
<connection>
<GID>5859</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>111,-1132.5,111,-1130.5</points>
<connection>
<GID>5976</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>111,-1114,111,-1112</points>
<connection>
<GID>6012</GID>
<name>OUT_0</name></connection>
<intersection>-1112 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>111,-1095,111,-1093</points>
<connection>
<GID>6048</GID>
<name>OUT_0</name></connection>
<intersection>-1093 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>111,-1076.5,111,-1074.5</points>
<connection>
<GID>6084</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-163,139,-163</points>
<connection>
<GID>4260</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-163,133,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-147.5,133,-147.5</points>
<connection>
<GID>4259</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-1225.5,118.5,-1060.5</points>
<connection>
<GID>5891</GID>
<name>N_in1</name></connection>
<connection>
<GID>5876</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 13</intersection>
<intersection>-1182 12</intersection>
<intersection>-1163 11</intersection>
<intersection>-1144.5 10</intersection>
<intersection>-1122.5 9</intersection>
<intersection>-1104 8</intersection>
<intersection>-1085 7</intersection>
<intersection>-1066.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>118.5,-1066.5,121,-1066.5</points>
<connection>
<GID>6086</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>118.5,-1085,121,-1085</points>
<connection>
<GID>6050</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118.5,-1104,121,-1104</points>
<connection>
<GID>6014</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>118.5,-1122.5,121,-1122.5</points>
<connection>
<GID>5978</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>118.5,-1144.5,121,-1144.5</points>
<connection>
<GID>5860</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>118.5,-1163,121,-1163</points>
<connection>
<GID>5836</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>118.5,-1182,121,-1182</points>
<connection>
<GID>5795</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>118.5,-1200.5,121,-1200.5</points>
<connection>
<GID>5759</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-163,162,-163</points>
<connection>
<GID>4262</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-163,156,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-147.5,156,-147.5</points>
<connection>
<GID>4261</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-1225.5,137,-1060.5</points>
<connection>
<GID>5892</GID>
<name>N_in1</name></connection>
<connection>
<GID>5877</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 6</intersection>
<intersection>-1190 7</intersection>
<intersection>-1171 8</intersection>
<intersection>-1152.5 9</intersection>
<intersection>-1130.5 10</intersection>
<intersection>-1112 11</intersection>
<intersection>-1093 12</intersection>
<intersection>-1074.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>134,-1208.5,137,-1208.5</points>
<intersection>134 14</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>134,-1190,137,-1190</points>
<intersection>134 15</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>134,-1171,137,-1171</points>
<intersection>134 16</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>134,-1152.5,137,-1152.5</points>
<intersection>134 17</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>134,-1130.5,137,-1130.5</points>
<intersection>134 20</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>134,-1112,137,-1112</points>
<intersection>134 21</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>134,-1093,137,-1093</points>
<intersection>134 22</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>134,-1074.5,137,-1074.5</points>
<intersection>134 23</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>134,-1210.5,134,-1208.5</points>
<connection>
<GID>5761</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>134,-1192,134,-1190</points>
<connection>
<GID>5797</GID>
<name>OUT_0</name></connection>
<intersection>-1190 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>134,-1173,134,-1171</points>
<connection>
<GID>5838</GID>
<name>OUT_0</name></connection>
<intersection>-1171 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>134,-1154.5,134,-1152.5</points>
<connection>
<GID>5861</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>134,-1132.5,134,-1130.5</points>
<connection>
<GID>5980</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>134,-1114,134,-1112</points>
<connection>
<GID>6016</GID>
<name>OUT_0</name></connection>
<intersection>-1112 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>134,-1095,134,-1093</points>
<connection>
<GID>6052</GID>
<name>OUT_0</name></connection>
<intersection>-1093 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>134,-1076.5,134,-1074.5</points>
<connection>
<GID>6088</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-163,185,-163</points>
<connection>
<GID>4264</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-163,179,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-147.5,179,-147.5</points>
<connection>
<GID>4263</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-1225.5,141,-1060.5</points>
<connection>
<GID>5893</GID>
<name>N_in1</name></connection>
<connection>
<GID>5878</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 13</intersection>
<intersection>-1182 12</intersection>
<intersection>-1163 11</intersection>
<intersection>-1144.5 10</intersection>
<intersection>-1122.5 9</intersection>
<intersection>-1104 8</intersection>
<intersection>-1085 7</intersection>
<intersection>-1066.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>141,-1066.5,144,-1066.5</points>
<connection>
<GID>6090</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>141,-1085,144,-1085</points>
<connection>
<GID>6054</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>141,-1104,144,-1104</points>
<connection>
<GID>6018</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>141,-1122.5,144,-1122.5</points>
<connection>
<GID>5982</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>141,-1144.5,144,-1144.5</points>
<connection>
<GID>5862</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>141,-1163,144,-1163</points>
<connection>
<GID>5841</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>141,-1182,144,-1182</points>
<connection>
<GID>5799</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>141,-1200.5,144,-1200.5</points>
<connection>
<GID>5763</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>1145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-163,210,-163</points>
<connection>
<GID>4266</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-163,204,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-147.5,204,-147.5</points>
<connection>
<GID>4265</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-1225,160,-1060.5</points>
<connection>
<GID>5894</GID>
<name>N_in1</name></connection>
<connection>
<GID>5879</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 6</intersection>
<intersection>-1190 7</intersection>
<intersection>-1171 8</intersection>
<intersection>-1152.5 9</intersection>
<intersection>-1130.5 10</intersection>
<intersection>-1112 11</intersection>
<intersection>-1093 12</intersection>
<intersection>-1074.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>157,-1208.5,160,-1208.5</points>
<intersection>157 14</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>157,-1190,160,-1190</points>
<intersection>157 15</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>157,-1171,160,-1171</points>
<intersection>157 16</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,-1152.5,160,-1152.5</points>
<intersection>157 17</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>157,-1130.5,160,-1130.5</points>
<intersection>157 20</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>157,-1112,160,-1112</points>
<intersection>157 21</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>157,-1093,160,-1093</points>
<intersection>157 22</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>157,-1074.5,160,-1074.5</points>
<intersection>157 23</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>157,-1210.5,157,-1208.5</points>
<connection>
<GID>5765</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>157,-1192,157,-1190</points>
<connection>
<GID>5801</GID>
<name>OUT_0</name></connection>
<intersection>-1190 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>157,-1173,157,-1171</points>
<connection>
<GID>5843</GID>
<name>OUT_0</name></connection>
<intersection>-1171 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>157,-1154.5,157,-1152.5</points>
<connection>
<GID>5863</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>157,-1132.5,157,-1130.5</points>
<connection>
<GID>5984</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>157,-1114,157,-1112</points>
<connection>
<GID>6020</GID>
<name>OUT_0</name></connection>
<intersection>-1112 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>157,-1095,157,-1093</points>
<connection>
<GID>6056</GID>
<name>OUT_0</name></connection>
<intersection>-1093 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>157,-1076.5,157,-1074.5</points>
<connection>
<GID>6092</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-163,233,-163</points>
<connection>
<GID>4268</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-163,227,-147.5</points>
<intersection>-163 1</intersection>
<intersection>-147.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-147.5,227,-147.5</points>
<connection>
<GID>4267</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-1225,165,-1060.5</points>
<connection>
<GID>5895</GID>
<name>N_in1</name></connection>
<connection>
<GID>5880</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 13</intersection>
<intersection>-1182 12</intersection>
<intersection>-1163 11</intersection>
<intersection>-1144.5 10</intersection>
<intersection>-1122.5 9</intersection>
<intersection>-1104 8</intersection>
<intersection>-1085 7</intersection>
<intersection>-1066.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>165,-1066.5,167,-1066.5</points>
<connection>
<GID>6094</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>165,-1085,167,-1085</points>
<connection>
<GID>6058</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>165,-1104,167,-1104</points>
<connection>
<GID>6022</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>165,-1122.5,167,-1122.5</points>
<connection>
<GID>5986</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>165,-1144.5,167,-1144.5</points>
<connection>
<GID>5864</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>165,-1163,167,-1163</points>
<connection>
<GID>5845</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>165,-1182,167,-1182</points>
<connection>
<GID>5803</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>165,-1200.5,167,-1200.5</points>
<connection>
<GID>5767</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>1147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-150.5,220,-150.5</points>
<connection>
<GID>4267</GID>
<name>clock</name></connection>
<connection>
<GID>4265</GID>
<name>clock</name></connection>
<connection>
<GID>4263</GID>
<name>clock</name></connection>
<connection>
<GID>4261</GID>
<name>clock</name></connection>
<connection>
<GID>4259</GID>
<name>clock</name></connection>
<connection>
<GID>4257</GID>
<name>clock</name></connection>
<connection>
<GID>4255</GID>
<name>clock</name></connection>
<connection>
<GID>4253</GID>
<name>clock</name></connection>
<connection>
<GID>4251</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-1224.5,183,-1060.5</points>
<connection>
<GID>5896</GID>
<name>N_in1</name></connection>
<connection>
<GID>5882</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 16</intersection>
<intersection>-1190 15</intersection>
<intersection>-1171 14</intersection>
<intersection>-1152.5 13</intersection>
<intersection>-1130.5 12</intersection>
<intersection>-1112 11</intersection>
<intersection>-1093 10</intersection>
<intersection>-1074.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>180,-1074.5,183,-1074.5</points>
<intersection>180 26</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>180,-1093,183,-1093</points>
<intersection>180 25</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>180,-1112,183,-1112</points>
<intersection>180 24</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>180,-1130.5,183,-1130.5</points>
<intersection>180 23</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>180,-1152.5,183,-1152.5</points>
<intersection>180 20</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>180,-1171,183,-1171</points>
<intersection>180 19</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>180,-1190,183,-1190</points>
<intersection>180 18</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>180,-1208.5,183,-1208.5</points>
<intersection>180 17</intersection>
<intersection>183 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>180,-1210.5,180,-1208.5</points>
<connection>
<GID>5769</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>180,-1192,180,-1190</points>
<connection>
<GID>5805</GID>
<name>OUT_0</name></connection>
<intersection>-1190 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>180,-1173,180,-1171</points>
<connection>
<GID>5846</GID>
<name>OUT_0</name></connection>
<intersection>-1171 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>180,-1154.5,180,-1152.5</points>
<connection>
<GID>5865</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>180,-1132.5,180,-1130.5</points>
<connection>
<GID>5988</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>180,-1114,180,-1112</points>
<connection>
<GID>6024</GID>
<name>OUT_0</name></connection>
<intersection>-1112 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>180,-1095,180,-1093</points>
<connection>
<GID>6060</GID>
<name>OUT_0</name></connection>
<intersection>-1093 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>180,-1076.5,180,-1074.5</points>
<connection>
<GID>6096</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>1148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-160,231,-160</points>
<connection>
<GID>4268</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4266</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4264</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4262</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4260</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4258</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4256</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4254</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4252</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-1224.5,187.5,-1060.5</points>
<connection>
<GID>5897</GID>
<name>N_in1</name></connection>
<connection>
<GID>5881</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 13</intersection>
<intersection>-1182 12</intersection>
<intersection>-1163 11</intersection>
<intersection>-1144.5 10</intersection>
<intersection>-1122.5 9</intersection>
<intersection>-1104 8</intersection>
<intersection>-1085 7</intersection>
<intersection>-1066.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>187.5,-1066.5,192,-1066.5</points>
<connection>
<GID>6098</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>187.5,-1085,192,-1085</points>
<connection>
<GID>6062</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187.5,-1104,192,-1104</points>
<connection>
<GID>6026</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>187.5,-1122.5,192,-1122.5</points>
<connection>
<GID>5990</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>187.5,-1144.5,192,-1144.5</points>
<connection>
<GID>5866</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>187.5,-1163,192,-1163</points>
<connection>
<GID>5848</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>187.5,-1182,192,-1182</points>
<connection>
<GID>5807</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>187.5,-1200.5,192,-1200.5</points>
<connection>
<GID>5771</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-144.5,68,-144.5</points>
<connection>
<GID>4272</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-144.5,62,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-129,62,-129</points>
<connection>
<GID>4271</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-1224,208.5,-1061</points>
<connection>
<GID>5898</GID>
<name>N_in1</name></connection>
<connection>
<GID>5883</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 6</intersection>
<intersection>-1190 7</intersection>
<intersection>-1171 8</intersection>
<intersection>-1152.5 9</intersection>
<intersection>-1130.5 10</intersection>
<intersection>-1112 11</intersection>
<intersection>-1093 12</intersection>
<intersection>-1074.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>205,-1208.5,208.5,-1208.5</points>
<intersection>205 14</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205,-1190,208.5,-1190</points>
<intersection>205 15</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>205,-1171,208.5,-1171</points>
<intersection>205 16</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>205,-1152.5,208.5,-1152.5</points>
<intersection>205 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>205,-1130.5,208.5,-1130.5</points>
<intersection>205 20</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205,-1112,208.5,-1112</points>
<intersection>205 21</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>205,-1093,208.5,-1093</points>
<intersection>205 22</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>205,-1074.5,208.5,-1074.5</points>
<intersection>205 23</intersection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>205,-1210.5,205,-1208.5</points>
<connection>
<GID>5773</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>205,-1192,205,-1190</points>
<connection>
<GID>5809</GID>
<name>OUT_0</name></connection>
<intersection>-1190 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>205,-1173,205,-1171</points>
<connection>
<GID>5849</GID>
<name>OUT_0</name></connection>
<intersection>-1171 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>205,-1154.5,205,-1152.5</points>
<connection>
<GID>5867</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>205,-1132.5,205,-1130.5</points>
<connection>
<GID>5992</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>205,-1114,205,-1112</points>
<connection>
<GID>6028</GID>
<name>OUT_0</name></connection>
<intersection>-1112 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>205,-1095,205,-1093</points>
<connection>
<GID>6064</GID>
<name>OUT_0</name></connection>
<intersection>-1093 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>205,-1076.5,205,-1074.5</points>
<connection>
<GID>6100</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-144.5,91,-144.5</points>
<connection>
<GID>4274</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-144.5,85,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-129,85,-129</points>
<connection>
<GID>4273</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-1224,212,-1061</points>
<connection>
<GID>5899</GID>
<name>N_in1</name></connection>
<connection>
<GID>5900</GID>
<name>N_in0</name></connection>
<intersection>-1200.5 11</intersection>
<intersection>-1182 10</intersection>
<intersection>-1163 9</intersection>
<intersection>-1144.5 7</intersection>
<intersection>-1122.5 6</intersection>
<intersection>-1104 5</intersection>
<intersection>-1085 4</intersection>
<intersection>-1066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-1066.5,215,-1066.5</points>
<connection>
<GID>6102</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>212,-1085,215,-1085</points>
<connection>
<GID>6066</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>212,-1104,215,-1104</points>
<connection>
<GID>6030</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>212,-1122.5,215,-1122.5</points>
<connection>
<GID>5994</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>212,-1144.5,215,-1144.5</points>
<connection>
<GID>5868</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>212,-1163,215,-1163</points>
<connection>
<GID>5850</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>212,-1182,215,-1182</points>
<connection>
<GID>5811</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>212,-1200.5,215,-1200.5</points>
<connection>
<GID>5775</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>1151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-144.5,116,-144.5</points>
<connection>
<GID>4276</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-144.5,110,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-129,110,-129</points>
<connection>
<GID>4275</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-1224,233,-1062</points>
<connection>
<GID>5901</GID>
<name>N_in1</name></connection>
<connection>
<GID>5884</GID>
<name>N_in0</name></connection>
<intersection>-1208.5 11</intersection>
<intersection>-1190 10</intersection>
<intersection>-1171 9</intersection>
<intersection>-1152.5 8</intersection>
<intersection>-1130.5 7</intersection>
<intersection>-1112 6</intersection>
<intersection>-1093 5</intersection>
<intersection>-1074.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>228,-1074.5,233,-1074.5</points>
<intersection>228 21</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-1093,233,-1093</points>
<intersection>228 20</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>228,-1112,233,-1112</points>
<intersection>228 19</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>228,-1130.5,233,-1130.5</points>
<intersection>228 18</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>228,-1152.5,233,-1152.5</points>
<intersection>228 15</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>228,-1171,233,-1171</points>
<intersection>228 14</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>228,-1190,233,-1190</points>
<intersection>228 13</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>228,-1208.5,233,-1208.5</points>
<intersection>228 12</intersection>
<intersection>233 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>228,-1210.5,228,-1208.5</points>
<connection>
<GID>5777</GID>
<name>OUT_0</name></connection>
<intersection>-1208.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>228,-1192,228,-1190</points>
<connection>
<GID>5813</GID>
<name>OUT_0</name></connection>
<intersection>-1190 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>228,-1173,228,-1171</points>
<connection>
<GID>5851</GID>
<name>OUT_0</name></connection>
<intersection>-1171 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>228,-1154.5,228,-1152.5</points>
<connection>
<GID>5869</GID>
<name>OUT_0</name></connection>
<intersection>-1152.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>228,-1132.5,228,-1130.5</points>
<connection>
<GID>5996</GID>
<name>OUT_0</name></connection>
<intersection>-1130.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>228,-1114,228,-1112</points>
<connection>
<GID>6032</GID>
<name>OUT_0</name></connection>
<intersection>-1112 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>228,-1095,228,-1093</points>
<connection>
<GID>6068</GID>
<name>OUT_0</name></connection>
<intersection>-1093 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>228,-1076.5,228,-1074.5</points>
<connection>
<GID>6104</GID>
<name>OUT_0</name></connection>
<intersection>-1074.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>1152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-144.5,139,-144.5</points>
<connection>
<GID>4278</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-144.5,133,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-129,133,-129</points>
<connection>
<GID>4277</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4232</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-124,-1068.5,22.5,-1068.5</points>
<connection>
<GID>6070</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-1220,-124,-1068.5</points>
<connection>
<GID>5907</GID>
<name>OUT_15</name></connection>
<intersection>-1078 4</intersection>
<intersection>-1068.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-1078,34,-1078</points>
<connection>
<GID>6072</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>1153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-144.5,162,-144.5</points>
<connection>
<GID>4280</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-144.5,156,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-129,156,-129</points>
<connection>
<GID>4279</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4233</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-123,-1087,22.5,-1087</points>
<connection>
<GID>6034</GID>
<name>IN_0</name></connection>
<intersection>-123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-123,-1221,-123,-1087</points>
<intersection>-1221 6</intersection>
<intersection>-1096.5 5</intersection>
<intersection>-1087 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-123,-1096.5,34,-1096.5</points>
<connection>
<GID>6036</GID>
<name>IN_0</name></connection>
<intersection>-123 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-1221,-123,-1221</points>
<connection>
<GID>5907</GID>
<name>OUT_14</name></connection>
<intersection>-123 4</intersection></hsegment></shape></wire>
<wire>
<ID>1154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-144.5,185,-144.5</points>
<connection>
<GID>4282</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-144.5,179,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-129,179,-129</points>
<connection>
<GID>4281</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4234</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-122,-1106,22.5,-1106</points>
<connection>
<GID>5998</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-1222,-122,-1106</points>
<intersection>-1222 6</intersection>
<intersection>-1115.5 4</intersection>
<intersection>-1106 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-1115.5,34,-1115.5</points>
<connection>
<GID>6000</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-1222,-122,-1222</points>
<connection>
<GID>5907</GID>
<name>OUT_13</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>1155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-144.5,210,-144.5</points>
<connection>
<GID>4284</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-144.5,204,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-129,204,-129</points>
<connection>
<GID>4283</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4235</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-121,-1124.5,22.5,-1124.5</points>
<connection>
<GID>5938</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-1223,-121,-1124.5</points>
<intersection>-1223 5</intersection>
<intersection>-1134 4</intersection>
<intersection>-1124.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-1134,34,-1134</points>
<connection>
<GID>5943</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1223,-121,-1223</points>
<connection>
<GID>5907</GID>
<name>OUT_12</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>1156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-144.5,233,-144.5</points>
<connection>
<GID>4286</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-144.5,227,-129</points>
<intersection>-144.5 1</intersection>
<intersection>-129 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-129,227,-129</points>
<connection>
<GID>4285</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-1146.5,22.5,-1146.5</points>
<connection>
<GID>5852</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-1224,-120,-1146.5</points>
<intersection>-1224 6</intersection>
<intersection>-1156 4</intersection>
<intersection>-1146.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-120,-1156,33.5,-1156</points>
<connection>
<GID>5853</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-1224,-120,-1224</points>
<connection>
<GID>5907</GID>
<name>OUT_11</name></connection>
<intersection>-120 3</intersection></hsegment></shape></wire>
<wire>
<ID>1157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-132,220,-132</points>
<connection>
<GID>4277</GID>
<name>clock</name></connection>
<connection>
<GID>4275</GID>
<name>clock</name></connection>
<connection>
<GID>4273</GID>
<name>clock</name></connection>
<connection>
<GID>4271</GID>
<name>clock</name></connection>
<connection>
<GID>4269</GID>
<name>OUT</name></connection>
<connection>
<GID>4285</GID>
<name>clock</name></connection>
<connection>
<GID>4283</GID>
<name>clock</name></connection>
<connection>
<GID>4281</GID>
<name>clock</name></connection>
<connection>
<GID>4279</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,-1165,22.5,-1165</points>
<connection>
<GID>5816</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-1225,-119,-1165</points>
<intersection>-1225 5</intersection>
<intersection>-1174.5 4</intersection>
<intersection>-1165 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-1174.5,33.5,-1174.5</points>
<connection>
<GID>5818</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1225,-119,-1225</points>
<connection>
<GID>5907</GID>
<name>OUT_10</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>1158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-141.5,231,-141.5</points>
<connection>
<GID>4278</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4276</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4274</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4272</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4270</GID>
<name>OUT</name></connection>
<connection>
<GID>4286</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4284</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4282</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4280</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118,-1184,22.5,-1184</points>
<connection>
<GID>5779</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118,-1226,-118,-1184</points>
<intersection>-1226 5</intersection>
<intersection>-1193.5 4</intersection>
<intersection>-1184 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118,-1193.5,33.5,-1193.5</points>
<connection>
<GID>5781</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1226,-118,-1226</points>
<connection>
<GID>5907</GID>
<name>OUT_9</name></connection>
<intersection>-118 3</intersection></hsegment></shape></wire>
<wire>
<ID>1159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-278.5,68,-278.5</points>
<connection>
<GID>4290</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-278.5,62,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-263,62,-263</points>
<connection>
<GID>4289</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-117,-1202.5,22.5,-1202.5</points>
<connection>
<GID>6106</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-1227,-117,-1202.5</points>
<intersection>-1227 5</intersection>
<intersection>-1212 4</intersection>
<intersection>-1202.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-1212,33.5,-1212</points>
<connection>
<GID>6108</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1227,-117,-1227</points>
<connection>
<GID>5907</GID>
<name>OUT_8</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>1160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-278.5,91,-278.5</points>
<connection>
<GID>4292</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-278.5,85,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-263,85,-263</points>
<connection>
<GID>4291</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-1226,21.5,-1061</points>
<connection>
<GID>5905</GID>
<name>N_in1</name></connection>
<connection>
<GID>5903</GID>
<name>N_in0</name></connection>
<intersection>-1204.5 10</intersection>
<intersection>-1186 9</intersection>
<intersection>-1167 8</intersection>
<intersection>-1148.5 7</intersection>
<intersection>-1126.5 6</intersection>
<intersection>-1108 5</intersection>
<intersection>-1089 4</intersection>
<intersection>-1070.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-1070.5,22.5,-1070.5</points>
<connection>
<GID>6070</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-1089,22.5,-1089</points>
<connection>
<GID>6034</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>21.5,-1108,22.5,-1108</points>
<connection>
<GID>5998</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-1126.5,22.5,-1126.5</points>
<connection>
<GID>5938</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21.5,-1148.5,22.5,-1148.5</points>
<connection>
<GID>5852</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>21.5,-1167,22.5,-1167</points>
<connection>
<GID>5816</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>21.5,-1186,22.5,-1186</points>
<connection>
<GID>5779</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>21.5,-1204.5,22.5,-1204.5</points>
<connection>
<GID>6106</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-278.5,116,-278.5</points>
<connection>
<GID>4294</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-278.5,110,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-263,110,-263</points>
<connection>
<GID>4293</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-1226,31.5,-1061</points>
<connection>
<GID>5904</GID>
<name>N_in1</name></connection>
<connection>
<GID>5902</GID>
<name>N_in0</name></connection>
<intersection>-1214 3</intersection>
<intersection>-1195.5 5</intersection>
<intersection>-1176.5 7</intersection>
<intersection>-1158 9</intersection>
<intersection>-1136 11</intersection>
<intersection>-1117.5 13</intersection>
<intersection>-1098.5 15</intersection>
<intersection>-1080 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-1214,33.5,-1214</points>
<connection>
<GID>6108</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-1195.5,33.5,-1195.5</points>
<connection>
<GID>5781</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31.5,-1176.5,33.5,-1176.5</points>
<connection>
<GID>5818</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>31.5,-1158,33.5,-1158</points>
<connection>
<GID>5853</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>31.5,-1136,34,-1136</points>
<connection>
<GID>5943</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>31.5,-1117.5,34,-1117.5</points>
<connection>
<GID>6000</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>31.5,-1098.5,34,-1098.5</points>
<connection>
<GID>6036</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>31.5,-1080,34,-1080</points>
<connection>
<GID>6072</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-278.5,139,-278.5</points>
<connection>
<GID>4296</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-278.5,133,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-263,133,-263</points>
<connection>
<GID>4295</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1313.5,63,-1313.5</points>
<connection>
<GID>6003</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1313.5,57,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1298,57,-1298</points>
<connection>
<GID>5991</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-278.5,162,-278.5</points>
<connection>
<GID>4298</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-278.5,156,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-263,156,-263</points>
<connection>
<GID>4297</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1313.5,86,-1313.5</points>
<connection>
<GID>6029</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1313.5,80,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1298,80,-1298</points>
<connection>
<GID>6027</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-278.5,185,-278.5</points>
<connection>
<GID>4300</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-278.5,179,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-263,179,-263</points>
<connection>
<GID>4299</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1313.5,111,-1313.5</points>
<connection>
<GID>6037</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1313.5,105,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1298,105,-1298</points>
<connection>
<GID>6033</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-278.5,210,-278.5</points>
<connection>
<GID>1666</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-278.5,204,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-263,204,-263</points>
<connection>
<GID>1665</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1313.5,134,-1313.5</points>
<connection>
<GID>6045</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1313.5,128,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1298,128,-1298</points>
<connection>
<GID>6041</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-278.5,233,-278.5</points>
<connection>
<GID>1668</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-278.5,227,-263</points>
<intersection>-278.5 1</intersection>
<intersection>-263 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-263,227,-263</points>
<connection>
<GID>1667</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1313.5,157,-1313.5</points>
<connection>
<GID>6051</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1313.5,151,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1298,151,-1298</points>
<connection>
<GID>6047</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>1167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-266,220,-266</points>
<connection>
<GID>1667</GID>
<name>clock</name></connection>
<connection>
<GID>1665</GID>
<name>clock</name></connection>
<connection>
<GID>4299</GID>
<name>clock</name></connection>
<connection>
<GID>4297</GID>
<name>clock</name></connection>
<connection>
<GID>4295</GID>
<name>clock</name></connection>
<connection>
<GID>4293</GID>
<name>clock</name></connection>
<connection>
<GID>4291</GID>
<name>clock</name></connection>
<connection>
<GID>4289</GID>
<name>clock</name></connection>
<connection>
<GID>4287</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1313.5,180,-1313.5</points>
<connection>
<GID>6055</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1313.5,174,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1298,174,-1298</points>
<connection>
<GID>6053</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>1168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-275.5,231,-275.5</points>
<connection>
<GID>1668</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1666</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4300</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4298</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4296</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4294</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4292</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4290</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>4288</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1313.5,205,-1313.5</points>
<connection>
<GID>6059</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1313.5,199,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1298,199,-1298</points>
<connection>
<GID>6057</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>1169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-260,68,-260</points>
<connection>
<GID>1672</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-260,62,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-244.5,62,-244.5</points>
<connection>
<GID>1671</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1313.5,228,-1313.5</points>
<connection>
<GID>6063</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1313.5,222,-1298</points>
<intersection>-1313.5 1</intersection>
<intersection>-1298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1298,222,-1298</points>
<connection>
<GID>6061</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>1170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-260,91,-260</points>
<connection>
<GID>1674</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-260,85,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-244.5,85,-244.5</points>
<connection>
<GID>1673</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1301,215,-1301</points>
<connection>
<GID>6061</GID>
<name>clock</name></connection>
<connection>
<GID>6057</GID>
<name>clock</name></connection>
<connection>
<GID>6053</GID>
<name>clock</name></connection>
<connection>
<GID>6047</GID>
<name>clock</name></connection>
<connection>
<GID>6041</GID>
<name>clock</name></connection>
<connection>
<GID>6033</GID>
<name>clock</name></connection>
<connection>
<GID>6027</GID>
<name>clock</name></connection>
<connection>
<GID>5991</GID>
<name>clock</name></connection>
<connection>
<GID>5985</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-260,116,-260</points>
<connection>
<GID>1676</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-260,110,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-244.5,110,-244.5</points>
<connection>
<GID>1675</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1310.5,226,-1310.5</points>
<connection>
<GID>6063</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6059</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6055</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6051</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6045</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6037</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6029</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6003</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5987</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-260,139,-260</points>
<connection>
<GID>1678</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-260,133,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-244.5,133,-244.5</points>
<connection>
<GID>1677</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1295,63,-1295</points>
<connection>
<GID>6071</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1295,57,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1279.5,57,-1279.5</points>
<connection>
<GID>6069</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>1173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-260,162,-260</points>
<connection>
<GID>1680</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-260,156,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-244.5,156,-244.5</points>
<connection>
<GID>1679</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1295,86,-1295</points>
<connection>
<GID>6075</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1295,80,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1279.5,80,-1279.5</points>
<connection>
<GID>6073</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>1174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-260,185,-260</points>
<connection>
<GID>1682</GID>
<name>IN_0</name></connection>
<intersection>179 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>179,-260,179,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>178,-244.5,179,-244.5</points>
<connection>
<GID>1681</GID>
<name>OUT_0</name></connection>
<intersection>179 2</intersection></hsegment></shape></wire>
<wire>
<ID>4254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1295,111,-1295</points>
<connection>
<GID>6079</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1295,105,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1279.5,105,-1279.5</points>
<connection>
<GID>6077</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>1175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-260,210,-260</points>
<connection>
<GID>1684</GID>
<name>IN_0</name></connection>
<intersection>204 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204,-260,204,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-244.5,204,-244.5</points>
<connection>
<GID>1683</GID>
<name>OUT_0</name></connection>
<intersection>204 2</intersection></hsegment></shape></wire>
<wire>
<ID>4255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1295,134,-1295</points>
<connection>
<GID>6083</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1295,128,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1279.5,128,-1279.5</points>
<connection>
<GID>6081</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>1176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227,-260,233,-260</points>
<connection>
<GID>1686</GID>
<name>IN_0</name></connection>
<intersection>227 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227,-260,227,-244.5</points>
<intersection>-260 1</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>226,-244.5,227,-244.5</points>
<connection>
<GID>1685</GID>
<name>OUT_0</name></connection>
<intersection>227 2</intersection></hsegment></shape></wire>
<wire>
<ID>4256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1295,157,-1295</points>
<connection>
<GID>6087</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1295,151,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1279.5,151,-1279.5</points>
<connection>
<GID>6085</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1295,180,-1295</points>
<connection>
<GID>6091</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1295,174,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1279.5,174,-1279.5</points>
<connection>
<GID>6089</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1295,205,-1295</points>
<connection>
<GID>6095</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1295,199,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1279.5,199,-1279.5</points>
<connection>
<GID>6093</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1295,228,-1295</points>
<connection>
<GID>6099</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1295,222,-1279.5</points>
<intersection>-1295 1</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1279.5,222,-1279.5</points>
<connection>
<GID>6097</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1282.5,215,-1282.5</points>
<connection>
<GID>6097</GID>
<name>clock</name></connection>
<connection>
<GID>6093</GID>
<name>clock</name></connection>
<connection>
<GID>6089</GID>
<name>clock</name></connection>
<connection>
<GID>6085</GID>
<name>clock</name></connection>
<connection>
<GID>6081</GID>
<name>clock</name></connection>
<connection>
<GID>6077</GID>
<name>clock</name></connection>
<connection>
<GID>6073</GID>
<name>clock</name></connection>
<connection>
<GID>6069</GID>
<name>clock</name></connection>
<connection>
<GID>6065</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1292,226,-1292</points>
<connection>
<GID>6099</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6095</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6091</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6087</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6083</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6079</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6075</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6071</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6067</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1276,63,-1276</points>
<connection>
<GID>6107</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1276,57,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1260.5,57,-1260.5</points>
<connection>
<GID>6105</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>4263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1276,86,-1276</points>
<connection>
<GID>6111</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1276,80,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1260.5,80,-1260.5</points>
<connection>
<GID>6109</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>4264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1276,111,-1276</points>
<connection>
<GID>6115</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1276,105,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1260.5,105,-1260.5</points>
<connection>
<GID>6113</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>4265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1276,134,-1276</points>
<connection>
<GID>6119</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1276,128,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1260.5,128,-1260.5</points>
<connection>
<GID>6117</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1276,157,-1276</points>
<connection>
<GID>5760</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1276,151,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1260.5,151,-1260.5</points>
<connection>
<GID>6121</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4267</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1276,180,-1276</points>
<connection>
<GID>5764</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1276,174,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1260.5,174,-1260.5</points>
<connection>
<GID>5762</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1276,205,-1276</points>
<connection>
<GID>5768</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1276,199,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1260.5,199,-1260.5</points>
<connection>
<GID>5766</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1276,228,-1276</points>
<connection>
<GID>5772</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1276,222,-1260.5</points>
<intersection>-1276 1</intersection>
<intersection>-1260.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1260.5,222,-1260.5</points>
<connection>
<GID>5770</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1263.5,215,-1263.5</points>
<connection>
<GID>6121</GID>
<name>clock</name></connection>
<connection>
<GID>6117</GID>
<name>clock</name></connection>
<connection>
<GID>6113</GID>
<name>clock</name></connection>
<connection>
<GID>6109</GID>
<name>clock</name></connection>
<connection>
<GID>6105</GID>
<name>clock</name></connection>
<connection>
<GID>6101</GID>
<name>OUT</name></connection>
<connection>
<GID>5770</GID>
<name>clock</name></connection>
<connection>
<GID>5766</GID>
<name>clock</name></connection>
<connection>
<GID>5762</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1273,226,-1273</points>
<connection>
<GID>6119</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6115</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6111</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6107</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6103</GID>
<name>OUT</name></connection>
<connection>
<GID>5772</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5768</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5764</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5760</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4272</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1257.5,63,-1257.5</points>
<connection>
<GID>5780</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1257.5,57,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1242,57,-1242</points>
<connection>
<GID>5778</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>4273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1257.5,86,-1257.5</points>
<connection>
<GID>5784</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1257.5,80,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1242,80,-1242</points>
<connection>
<GID>5782</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>4274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1257.5,111,-1257.5</points>
<connection>
<GID>5788</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1257.5,105,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1242,105,-1242</points>
<connection>
<GID>5786</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>4275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1257.5,134,-1257.5</points>
<connection>
<GID>5792</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1257.5,128,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1242,128,-1242</points>
<connection>
<GID>5790</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1257.5,157,-1257.5</points>
<connection>
<GID>5796</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1257.5,151,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1242,151,-1242</points>
<connection>
<GID>5794</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1257.5,180,-1257.5</points>
<connection>
<GID>5800</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1257.5,174,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1242,174,-1242</points>
<connection>
<GID>5798</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1257.5,205,-1257.5</points>
<connection>
<GID>5804</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1257.5,199,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1242,199,-1242</points>
<connection>
<GID>5802</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4279</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1257.5,228,-1257.5</points>
<connection>
<GID>5808</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1257.5,222,-1242</points>
<intersection>-1257.5 1</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1242,222,-1242</points>
<connection>
<GID>5806</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4280</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1245,215,-1245</points>
<connection>
<GID>5806</GID>
<name>clock</name></connection>
<connection>
<GID>5802</GID>
<name>clock</name></connection>
<connection>
<GID>5798</GID>
<name>clock</name></connection>
<connection>
<GID>5794</GID>
<name>clock</name></connection>
<connection>
<GID>5790</GID>
<name>clock</name></connection>
<connection>
<GID>5786</GID>
<name>clock</name></connection>
<connection>
<GID>5782</GID>
<name>clock</name></connection>
<connection>
<GID>5778</GID>
<name>clock</name></connection>
<connection>
<GID>5774</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-1254.5,226,-1254.5</points>
<connection>
<GID>5808</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5804</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5800</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5796</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5792</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5788</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5784</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5780</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5776</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1391.5,63,-1391.5</points>
<connection>
<GID>5817</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1391.5,57,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1376,57,-1376</points>
<connection>
<GID>5814</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>4283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1391.5,86,-1391.5</points>
<connection>
<GID>5822</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1391.5,80,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1376,80,-1376</points>
<connection>
<GID>5819</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>4284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1391.5,111,-1391.5</points>
<connection>
<GID>5827</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1391.5,105,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1376,105,-1376</points>
<connection>
<GID>5824</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>4285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1391.5,134,-1391.5</points>
<connection>
<GID>5832</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1391.5,128,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1376,128,-1376</points>
<connection>
<GID>5829</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1391.5,157,-1391.5</points>
<connection>
<GID>5837</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1391.5,151,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1376,151,-1376</points>
<connection>
<GID>5834</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1391.5,180,-1391.5</points>
<connection>
<GID>5842</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1391.5,174,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1376,174,-1376</points>
<connection>
<GID>5839</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1391.5,205,-1391.5</points>
<connection>
<GID>5909</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1391.5,199,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1376,199,-1376</points>
<connection>
<GID>5908</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1391.5,228,-1391.5</points>
<connection>
<GID>5911</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1391.5,222,-1376</points>
<intersection>-1391.5 1</intersection>
<intersection>-1376 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1376,222,-1376</points>
<connection>
<GID>5910</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1379,215,-1379</points>
<connection>
<GID>5910</GID>
<name>clock</name></connection>
<connection>
<GID>5908</GID>
<name>clock</name></connection>
<connection>
<GID>5839</GID>
<name>clock</name></connection>
<connection>
<GID>5834</GID>
<name>clock</name></connection>
<connection>
<GID>5829</GID>
<name>clock</name></connection>
<connection>
<GID>5824</GID>
<name>clock</name></connection>
<connection>
<GID>5819</GID>
<name>clock</name></connection>
<connection>
<GID>5814</GID>
<name>clock</name></connection>
<connection>
<GID>5810</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1388.5,226,-1388.5</points>
<connection>
<GID>5911</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5909</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5842</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5837</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5832</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5827</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5822</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5817</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5812</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1373,63,-1373</points>
<connection>
<GID>5915</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1373,57,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1357.5,57,-1357.5</points>
<connection>
<GID>5914</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>4293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1373,86,-1373</points>
<connection>
<GID>5917</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1373,80,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1357.5,80,-1357.5</points>
<connection>
<GID>5916</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>4294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1373,111,-1373</points>
<connection>
<GID>5919</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1373,105,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1357.5,105,-1357.5</points>
<connection>
<GID>5918</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>4295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1373,134,-1373</points>
<connection>
<GID>5921</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1373,128,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1357.5,128,-1357.5</points>
<connection>
<GID>5920</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1373,157,-1373</points>
<connection>
<GID>5923</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1373,151,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1357.5,151,-1357.5</points>
<connection>
<GID>5922</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1373,180,-1373</points>
<connection>
<GID>5925</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1373,174,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1357.5,174,-1357.5</points>
<connection>
<GID>5924</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1373,205,-1373</points>
<connection>
<GID>5927</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1373,199,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1357.5,199,-1357.5</points>
<connection>
<GID>5926</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1373,228,-1373</points>
<connection>
<GID>5929</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1373,222,-1357.5</points>
<intersection>-1373 1</intersection>
<intersection>-1357.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1357.5,222,-1357.5</points>
<connection>
<GID>5928</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1360.5,215,-1360.5</points>
<connection>
<GID>5928</GID>
<name>clock</name></connection>
<connection>
<GID>5926</GID>
<name>clock</name></connection>
<connection>
<GID>5924</GID>
<name>clock</name></connection>
<connection>
<GID>5922</GID>
<name>clock</name></connection>
<connection>
<GID>5920</GID>
<name>clock</name></connection>
<connection>
<GID>5918</GID>
<name>clock</name></connection>
<connection>
<GID>5916</GID>
<name>clock</name></connection>
<connection>
<GID>5914</GID>
<name>clock</name></connection>
<connection>
<GID>5912</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1370,226,-1370</points>
<connection>
<GID>5929</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5927</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5925</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5923</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5921</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5919</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5917</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5915</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5913</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1354,63,-1354</points>
<connection>
<GID>5825</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1354,57,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1338.5,57,-1338.5</points>
<connection>
<GID>5820</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>4303</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1354,86,-1354</points>
<connection>
<GID>5835</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1354,80,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1338.5,80,-1338.5</points>
<connection>
<GID>5830</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>4304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1354,111,-1354</points>
<connection>
<GID>5844</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1354,105,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1338.5,105,-1338.5</points>
<connection>
<GID>5840</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>4305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1354,134,-1354</points>
<connection>
<GID>5931</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1354,128,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1338.5,128,-1338.5</points>
<connection>
<GID>5847</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1354,157,-1354</points>
<connection>
<GID>5933</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1354,151,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1338.5,151,-1338.5</points>
<connection>
<GID>5932</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1354,180,-1354</points>
<connection>
<GID>5935</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1354,174,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1338.5,174,-1338.5</points>
<connection>
<GID>5934</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1354,205,-1354</points>
<connection>
<GID>5937</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1354,199,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1338.5,199,-1338.5</points>
<connection>
<GID>5936</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4309</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1354,228,-1354</points>
<connection>
<GID>5940</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1354,222,-1338.5</points>
<intersection>-1354 1</intersection>
<intersection>-1338.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1338.5,222,-1338.5</points>
<connection>
<GID>5939</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1341.5,215,-1341.5</points>
<connection>
<GID>5939</GID>
<name>clock</name></connection>
<connection>
<GID>5936</GID>
<name>clock</name></connection>
<connection>
<GID>5934</GID>
<name>clock</name></connection>
<connection>
<GID>5932</GID>
<name>clock</name></connection>
<connection>
<GID>5930</GID>
<name>OUT</name></connection>
<connection>
<GID>5847</GID>
<name>clock</name></connection>
<connection>
<GID>5840</GID>
<name>clock</name></connection>
<connection>
<GID>5830</GID>
<name>clock</name></connection>
<connection>
<GID>5820</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1351,226,-1351</points>
<connection>
<GID>5940</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5937</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5935</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5933</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5931</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5844</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5835</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5825</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5815</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-1335.5,63,-1335.5</points>
<connection>
<GID>5945</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-1335.5,57,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-1320,57,-1320</points>
<connection>
<GID>5944</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>4313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-1335.5,86,-1335.5</points>
<connection>
<GID>5947</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-1335.5,80,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1320,80,-1320</points>
<connection>
<GID>5946</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>4314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-1335.5,111,-1335.5</points>
<connection>
<GID>5950</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-1335.5,105,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-1320,105,-1320</points>
<connection>
<GID>5949</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>4315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-1335.5,134,-1335.5</points>
<connection>
<GID>5952</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-1335.5,128,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-1320,128,-1320</points>
<connection>
<GID>5951</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>4316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-1335.5,157,-1335.5</points>
<connection>
<GID>5955</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-1335.5,151,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-1320,151,-1320</points>
<connection>
<GID>5953</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>4317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-1335.5,180,-1335.5</points>
<connection>
<GID>5957</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-1335.5,174,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-1320,174,-1320</points>
<connection>
<GID>5956</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>4318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-1335.5,205,-1335.5</points>
<connection>
<GID>5959</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-1335.5,199,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-1320,199,-1320</points>
<connection>
<GID>5958</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>4319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-1335.5,228,-1335.5</points>
<connection>
<GID>5961</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-1335.5,222,-1320</points>
<intersection>-1335.5 1</intersection>
<intersection>-1320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-1320,222,-1320</points>
<connection>
<GID>5960</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>4320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-1323,215,-1323</points>
<connection>
<GID>5960</GID>
<name>clock</name></connection>
<connection>
<GID>5958</GID>
<name>clock</name></connection>
<connection>
<GID>5956</GID>
<name>clock</name></connection>
<connection>
<GID>5953</GID>
<name>clock</name></connection>
<connection>
<GID>5951</GID>
<name>clock</name></connection>
<connection>
<GID>5949</GID>
<name>clock</name></connection>
<connection>
<GID>5946</GID>
<name>clock</name></connection>
<connection>
<GID>5944</GID>
<name>clock</name></connection>
<connection>
<GID>5941</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1332.5,226,-1332.5</points>
<connection>
<GID>5961</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5959</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5957</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5955</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5952</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5950</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5947</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5945</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5942</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-1401.5,44.5,-1236.5</points>
<connection>
<GID>5989</GID>
<name>N_in1</name></connection>
<connection>
<GID>5962</GID>
<name>N_in0</name></connection>
<intersection>-1376 12</intersection>
<intersection>-1357.5 11</intersection>
<intersection>-1338.5 10</intersection>
<intersection>-1320 9</intersection>
<intersection>-1298 8</intersection>
<intersection>-1279.5 7</intersection>
<intersection>-1260.5 6</intersection>
<intersection>-1242 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-1242,50,-1242</points>
<connection>
<GID>5778</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>44.5,-1260.5,50,-1260.5</points>
<connection>
<GID>6105</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-1279.5,50,-1279.5</points>
<connection>
<GID>6069</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>44.5,-1298,50,-1298</points>
<connection>
<GID>5991</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>44.5,-1320,50,-1320</points>
<connection>
<GID>5944</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>44.5,-1338.5,50,-1338.5</points>
<connection>
<GID>5820</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>44.5,-1357.5,50,-1357.5</points>
<connection>
<GID>5914</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>44.5,-1376,50,-1376</points>
<connection>
<GID>5814</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-1401,67.5,-1236</points>
<connection>
<GID>5993</GID>
<name>N_in1</name></connection>
<connection>
<GID>5963</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 4</intersection>
<intersection>-1365 5</intersection>
<intersection>-1346 6</intersection>
<intersection>-1327.5 7</intersection>
<intersection>-1305.5 8</intersection>
<intersection>-1287 9</intersection>
<intersection>-1268 10</intersection>
<intersection>-1249.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63,-1383.5,67.5,-1383.5</points>
<intersection>63 12</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-1365,67.5,-1365</points>
<intersection>63 14</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>63,-1346,67.5,-1346</points>
<intersection>63 13</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>63,-1327.5,67.5,-1327.5</points>
<intersection>63 15</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>63,-1305.5,67.5,-1305.5</points>
<intersection>63 18</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-1287,67.5,-1287</points>
<intersection>63 19</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>63,-1268,67.5,-1268</points>
<intersection>63 20</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>63,-1249.5,67.5,-1249.5</points>
<intersection>63 21</intersection>
<intersection>67.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>63,-1386,63,-1383.5</points>
<connection>
<GID>5817</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>63,-1348.5,63,-1346</points>
<connection>
<GID>5825</GID>
<name>OUT_0</name></connection>
<intersection>-1346 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>63,-1367.5,63,-1365</points>
<connection>
<GID>5915</GID>
<name>OUT_0</name></connection>
<intersection>-1365 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>63,-1330,63,-1327.5</points>
<connection>
<GID>5945</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>63,-1308,63,-1305.5</points>
<connection>
<GID>6003</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>63,-1289.5,63,-1287</points>
<connection>
<GID>6071</GID>
<name>OUT_0</name></connection>
<intersection>-1287 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>63,-1270.5,63,-1268</points>
<connection>
<GID>6107</GID>
<name>OUT_0</name></connection>
<intersection>-1268 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>63,-1252,63,-1249.5</points>
<connection>
<GID>5780</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>4324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-1401,70.5,-1236.5</points>
<connection>
<GID>5995</GID>
<name>N_in1</name></connection>
<connection>
<GID>5964</GID>
<name>N_in0</name></connection>
<intersection>-1376 10</intersection>
<intersection>-1357.5 9</intersection>
<intersection>-1338.5 8</intersection>
<intersection>-1320 7</intersection>
<intersection>-1298 6</intersection>
<intersection>-1279.5 5</intersection>
<intersection>-1260.5 4</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70.5,-1242,73,-1242</points>
<connection>
<GID>5782</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-1260.5,73,-1260.5</points>
<connection>
<GID>6109</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-1279.5,73,-1279.5</points>
<connection>
<GID>6073</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>70.5,-1298,73,-1298</points>
<connection>
<GID>6027</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>70.5,-1320,73,-1320</points>
<connection>
<GID>5946</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>70.5,-1338.5,73,-1338.5</points>
<connection>
<GID>5830</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>70.5,-1357.5,73,-1357.5</points>
<connection>
<GID>5916</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>70.5,-1376,73,-1376</points>
<connection>
<GID>5819</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-1401,90,-1236</points>
<connection>
<GID>5997</GID>
<name>N_in1</name></connection>
<connection>
<GID>5965</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 6</intersection>
<intersection>-1365 7</intersection>
<intersection>-1346 8</intersection>
<intersection>-1327.5 9</intersection>
<intersection>-1305.5 10</intersection>
<intersection>-1287 11</intersection>
<intersection>-1268 12</intersection>
<intersection>-1249.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-1383.5,90,-1383.5</points>
<intersection>86 14</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>86,-1365,90,-1365</points>
<intersection>86 16</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>86,-1346,90,-1346</points>
<intersection>86 15</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>86,-1327.5,90,-1327.5</points>
<intersection>86 17</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>86,-1305.5,90,-1305.5</points>
<intersection>86 20</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>86,-1287,90,-1287</points>
<intersection>86 21</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>86,-1268,90,-1268</points>
<intersection>86 22</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>86,-1249.5,90,-1249.5</points>
<intersection>86 23</intersection>
<intersection>90 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>86,-1386,86,-1383.5</points>
<connection>
<GID>5822</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>86,-1348.5,86,-1346</points>
<connection>
<GID>5835</GID>
<name>OUT_0</name></connection>
<intersection>-1346 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>86,-1367.5,86,-1365</points>
<connection>
<GID>5917</GID>
<name>OUT_0</name></connection>
<intersection>-1365 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>86,-1330,86,-1327.5</points>
<connection>
<GID>5947</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>86,-1308,86,-1305.5</points>
<connection>
<GID>6029</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>86,-1289.5,86,-1287</points>
<connection>
<GID>6075</GID>
<name>OUT_0</name></connection>
<intersection>-1287 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>86,-1270.5,86,-1268</points>
<connection>
<GID>6111</GID>
<name>OUT_0</name></connection>
<intersection>-1268 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>86,-1252,86,-1249.5</points>
<connection>
<GID>5784</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-1401,93.5,-1236</points>
<connection>
<GID>5999</GID>
<name>N_in1</name></connection>
<connection>
<GID>5966</GID>
<name>N_in0</name></connection>
<intersection>-1376 13</intersection>
<intersection>-1357.5 12</intersection>
<intersection>-1338.5 11</intersection>
<intersection>-1320 10</intersection>
<intersection>-1298 9</intersection>
<intersection>-1279.5 8</intersection>
<intersection>-1260.5 7</intersection>
<intersection>-1242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>93.5,-1242,98,-1242</points>
<connection>
<GID>5786</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>93.5,-1260.5,98,-1260.5</points>
<connection>
<GID>6113</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>93.5,-1279.5,98,-1279.5</points>
<connection>
<GID>6077</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-1298,98,-1298</points>
<connection>
<GID>6033</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>93.5,-1320,98,-1320</points>
<connection>
<GID>5949</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>93.5,-1338.5,98,-1338.5</points>
<connection>
<GID>5840</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>93.5,-1357.5,98,-1357.5</points>
<connection>
<GID>5918</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>93.5,-1376,98,-1376</points>
<connection>
<GID>5824</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-1401,114.5,-1236.5</points>
<connection>
<GID>6001</GID>
<name>N_in1</name></connection>
<connection>
<GID>5967</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 6</intersection>
<intersection>-1365 7</intersection>
<intersection>-1346 8</intersection>
<intersection>-1327.5 9</intersection>
<intersection>-1305.5 10</intersection>
<intersection>-1287 11</intersection>
<intersection>-1268 12</intersection>
<intersection>-1249.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>111,-1383.5,114.5,-1383.5</points>
<intersection>111 14</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111,-1365,114.5,-1365</points>
<intersection>111 16</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111,-1346,114.5,-1346</points>
<intersection>111 15</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111,-1327.5,114.5,-1327.5</points>
<intersection>111 17</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,-1305.5,114.5,-1305.5</points>
<intersection>111 20</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>111,-1287,114.5,-1287</points>
<intersection>111 21</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>111,-1268,114.5,-1268</points>
<intersection>111 22</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111,-1249.5,114.5,-1249.5</points>
<intersection>111 23</intersection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>111,-1386,111,-1383.5</points>
<connection>
<GID>5827</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>111,-1348.5,111,-1346</points>
<connection>
<GID>5844</GID>
<name>OUT_0</name></connection>
<intersection>-1346 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>111,-1367.5,111,-1365</points>
<connection>
<GID>5919</GID>
<name>OUT_0</name></connection>
<intersection>-1365 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>111,-1330,111,-1327.5</points>
<connection>
<GID>5950</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>111,-1308,111,-1305.5</points>
<connection>
<GID>6037</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>111,-1289.5,111,-1287</points>
<connection>
<GID>6079</GID>
<name>OUT_0</name></connection>
<intersection>-1287 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>111,-1270.5,111,-1268</points>
<connection>
<GID>6115</GID>
<name>OUT_0</name></connection>
<intersection>-1268 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>111,-1252,111,-1249.5</points>
<connection>
<GID>5788</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-1401,118.5,-1236</points>
<connection>
<GID>6005</GID>
<name>N_in1</name></connection>
<connection>
<GID>5968</GID>
<name>N_in0</name></connection>
<intersection>-1376 13</intersection>
<intersection>-1357.5 12</intersection>
<intersection>-1338.5 11</intersection>
<intersection>-1320 10</intersection>
<intersection>-1298 9</intersection>
<intersection>-1279.5 8</intersection>
<intersection>-1260.5 7</intersection>
<intersection>-1242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>118.5,-1242,121,-1242</points>
<connection>
<GID>5790</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>118.5,-1260.5,121,-1260.5</points>
<connection>
<GID>6117</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118.5,-1279.5,121,-1279.5</points>
<connection>
<GID>6081</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>118.5,-1298,121,-1298</points>
<connection>
<GID>6041</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>118.5,-1320,121,-1320</points>
<connection>
<GID>5951</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>118.5,-1338.5,121,-1338.5</points>
<connection>
<GID>5847</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>118.5,-1357.5,121,-1357.5</points>
<connection>
<GID>5920</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>118.5,-1376,121,-1376</points>
<connection>
<GID>5829</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-1401,137,-1236</points>
<connection>
<GID>6007</GID>
<name>N_in1</name></connection>
<connection>
<GID>5969</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 6</intersection>
<intersection>-1365 7</intersection>
<intersection>-1346 8</intersection>
<intersection>-1327.5 9</intersection>
<intersection>-1305.5 10</intersection>
<intersection>-1287 11</intersection>
<intersection>-1268 12</intersection>
<intersection>-1249.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>134,-1383.5,137,-1383.5</points>
<intersection>134 14</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>134,-1365,137,-1365</points>
<intersection>134 15</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>134,-1346,137,-1346</points>
<intersection>134 16</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>134,-1327.5,137,-1327.5</points>
<intersection>134 17</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>134,-1305.5,137,-1305.5</points>
<intersection>134 20</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>134,-1287,137,-1287</points>
<intersection>134 21</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>134,-1268,137,-1268</points>
<intersection>134 22</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>134,-1249.5,137,-1249.5</points>
<intersection>134 23</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>134,-1386,134,-1383.5</points>
<connection>
<GID>5832</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>134,-1367.5,134,-1365</points>
<connection>
<GID>5921</GID>
<name>OUT_0</name></connection>
<intersection>-1365 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>134,-1348.5,134,-1346</points>
<connection>
<GID>5931</GID>
<name>OUT_0</name></connection>
<intersection>-1346 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>134,-1330,134,-1327.5</points>
<connection>
<GID>5952</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>134,-1308,134,-1305.5</points>
<connection>
<GID>6045</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>134,-1289.5,134,-1287</points>
<connection>
<GID>6083</GID>
<name>OUT_0</name></connection>
<intersection>-1287 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>134,-1270.5,134,-1268</points>
<connection>
<GID>6119</GID>
<name>OUT_0</name></connection>
<intersection>-1268 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>134,-1252,134,-1249.5</points>
<connection>
<GID>5792</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-1401,141,-1236</points>
<connection>
<GID>6009</GID>
<name>N_in1</name></connection>
<connection>
<GID>5971</GID>
<name>N_in0</name></connection>
<intersection>-1376 13</intersection>
<intersection>-1357.5 12</intersection>
<intersection>-1338.5 11</intersection>
<intersection>-1320 10</intersection>
<intersection>-1298 9</intersection>
<intersection>-1279.5 8</intersection>
<intersection>-1260.5 7</intersection>
<intersection>-1242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>141,-1242,144,-1242</points>
<connection>
<GID>5794</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>141,-1260.5,144,-1260.5</points>
<connection>
<GID>6121</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>141,-1279.5,144,-1279.5</points>
<connection>
<GID>6085</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>141,-1298,144,-1298</points>
<connection>
<GID>6047</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>141,-1320,144,-1320</points>
<connection>
<GID>5953</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>141,-1338.5,144,-1338.5</points>
<connection>
<GID>5932</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>141,-1357.5,144,-1357.5</points>
<connection>
<GID>5922</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>141,-1376,144,-1376</points>
<connection>
<GID>5834</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>4331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-1400.5,160,-1236</points>
<connection>
<GID>6011</GID>
<name>N_in1</name></connection>
<connection>
<GID>5973</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 6</intersection>
<intersection>-1365 7</intersection>
<intersection>-1346 8</intersection>
<intersection>-1327.5 9</intersection>
<intersection>-1305.5 10</intersection>
<intersection>-1287 11</intersection>
<intersection>-1268 12</intersection>
<intersection>-1249.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>157,-1383.5,160,-1383.5</points>
<intersection>157 15</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>157,-1365,160,-1365</points>
<intersection>157 16</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>157,-1346,160,-1346</points>
<intersection>157 17</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,-1327.5,160,-1327.5</points>
<intersection>157 18</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>157,-1305.5,160,-1305.5</points>
<intersection>157 21</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>157,-1287,160,-1287</points>
<intersection>157 22</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>157,-1268,160,-1268</points>
<intersection>157 23</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>157,-1249.5,160,-1249.5</points>
<intersection>157 14</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>157,-1252,157,-1249.5</points>
<connection>
<GID>5796</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>157,-1386,157,-1383.5</points>
<connection>
<GID>5837</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>157,-1367.5,157,-1365</points>
<connection>
<GID>5923</GID>
<name>OUT_0</name></connection>
<intersection>-1365 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>157,-1348.5,157,-1346</points>
<connection>
<GID>5933</GID>
<name>OUT_0</name></connection>
<intersection>-1346 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>157,-1330,157,-1327.5</points>
<connection>
<GID>5955</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>157,-1308,157,-1305.5</points>
<connection>
<GID>6051</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>157,-1289.5,157,-1287</points>
<connection>
<GID>6087</GID>
<name>OUT_0</name></connection>
<intersection>-1287 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>157,-1270.5,157,-1268</points>
<connection>
<GID>5760</GID>
<name>OUT_0</name></connection>
<intersection>-1268 12</intersection></vsegment></shape></wire>
<wire>
<ID>4332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-1400.5,165,-1236</points>
<connection>
<GID>6013</GID>
<name>N_in1</name></connection>
<connection>
<GID>5975</GID>
<name>N_in0</name></connection>
<intersection>-1376 13</intersection>
<intersection>-1357.5 12</intersection>
<intersection>-1338.5 11</intersection>
<intersection>-1320 10</intersection>
<intersection>-1298 9</intersection>
<intersection>-1279.5 8</intersection>
<intersection>-1260.5 7</intersection>
<intersection>-1242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>165,-1242,167,-1242</points>
<connection>
<GID>5798</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>165,-1260.5,167,-1260.5</points>
<connection>
<GID>5762</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>165,-1279.5,167,-1279.5</points>
<connection>
<GID>6089</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>165,-1298,167,-1298</points>
<connection>
<GID>6053</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>165,-1320,167,-1320</points>
<connection>
<GID>5956</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>165,-1338.5,167,-1338.5</points>
<connection>
<GID>5934</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>165,-1357.5,167,-1357.5</points>
<connection>
<GID>5924</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>165,-1376,167,-1376</points>
<connection>
<GID>5839</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>4333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-1400,183,-1236</points>
<connection>
<GID>6015</GID>
<name>N_in1</name></connection>
<connection>
<GID>5979</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 16</intersection>
<intersection>-1365 15</intersection>
<intersection>-1346 14</intersection>
<intersection>-1327.5 13</intersection>
<intersection>-1305.5 12</intersection>
<intersection>-1287 11</intersection>
<intersection>-1268 10</intersection>
<intersection>-1249.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>180,-1249.5,183,-1249.5</points>
<intersection>180 17</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>180,-1268,183,-1268</points>
<intersection>180 26</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>180,-1287,183,-1287</points>
<intersection>180 25</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>180,-1305.5,183,-1305.5</points>
<intersection>180 24</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>180,-1327.5,183,-1327.5</points>
<intersection>180 21</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>180,-1346,183,-1346</points>
<intersection>180 20</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>180,-1365,183,-1365</points>
<intersection>180 19</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>180,-1383.5,183,-1383.5</points>
<intersection>180 18</intersection>
<intersection>183 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>180,-1252,180,-1249.5</points>
<connection>
<GID>5800</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>180,-1386,180,-1383.5</points>
<connection>
<GID>5842</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>180,-1367.5,180,-1365</points>
<connection>
<GID>5925</GID>
<name>OUT_0</name></connection>
<intersection>-1365 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>180,-1348.5,180,-1346</points>
<connection>
<GID>5935</GID>
<name>OUT_0</name></connection>
<intersection>-1346 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>180,-1330,180,-1327.5</points>
<connection>
<GID>5957</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>180,-1308,180,-1305.5</points>
<connection>
<GID>6055</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>180,-1289.5,180,-1287</points>
<connection>
<GID>6091</GID>
<name>OUT_0</name></connection>
<intersection>-1287 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>180,-1270.5,180,-1268</points>
<connection>
<GID>5764</GID>
<name>OUT_0</name></connection>
<intersection>-1268 10</intersection></vsegment></shape></wire>
<wire>
<ID>4334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-1400,187.5,-1236</points>
<connection>
<GID>6017</GID>
<name>N_in1</name></connection>
<connection>
<GID>5977</GID>
<name>N_in0</name></connection>
<intersection>-1376 13</intersection>
<intersection>-1357.5 12</intersection>
<intersection>-1338.5 11</intersection>
<intersection>-1320 10</intersection>
<intersection>-1298 9</intersection>
<intersection>-1279.5 8</intersection>
<intersection>-1260.5 7</intersection>
<intersection>-1242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>187.5,-1242,192,-1242</points>
<connection>
<GID>5802</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>187.5,-1260.5,192,-1260.5</points>
<connection>
<GID>5766</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187.5,-1279.5,192,-1279.5</points>
<connection>
<GID>6093</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>187.5,-1298,192,-1298</points>
<connection>
<GID>6057</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>187.5,-1320,192,-1320</points>
<connection>
<GID>5958</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>187.5,-1338.5,192,-1338.5</points>
<connection>
<GID>5936</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>187.5,-1357.5,192,-1357.5</points>
<connection>
<GID>5926</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>187.5,-1376,192,-1376</points>
<connection>
<GID>5908</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-1399.5,208.5,-1236.5</points>
<connection>
<GID>6019</GID>
<name>N_in1</name></connection>
<connection>
<GID>5981</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 6</intersection>
<intersection>-1365 7</intersection>
<intersection>-1346 8</intersection>
<intersection>-1327.5 9</intersection>
<intersection>-1305.5 10</intersection>
<intersection>-1287 11</intersection>
<intersection>-1268 12</intersection>
<intersection>-1249.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>205,-1383.5,208.5,-1383.5</points>
<intersection>205 15</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205,-1365,208.5,-1365</points>
<intersection>205 16</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>205,-1346,208.5,-1346</points>
<intersection>205 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>205,-1327.5,208.5,-1327.5</points>
<intersection>205 18</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>205,-1305.5,208.5,-1305.5</points>
<intersection>205 21</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205,-1287,208.5,-1287</points>
<intersection>205 22</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>205,-1268,208.5,-1268</points>
<intersection>205 23</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>205,-1249.5,208.5,-1249.5</points>
<intersection>205 14</intersection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>205,-1252,205,-1249.5</points>
<connection>
<GID>5804</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>205,-1386,205,-1383.5</points>
<connection>
<GID>5909</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>205,-1367.5,205,-1365</points>
<connection>
<GID>5927</GID>
<name>OUT_0</name></connection>
<intersection>-1365 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>205,-1348.5,205,-1346</points>
<connection>
<GID>5937</GID>
<name>OUT_0</name></connection>
<intersection>-1346 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>205,-1330,205,-1327.5</points>
<connection>
<GID>5959</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>205,-1308,205,-1305.5</points>
<connection>
<GID>6059</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>205,-1289.5,205,-1287</points>
<connection>
<GID>6095</GID>
<name>OUT_0</name></connection>
<intersection>-1287 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>205,-1270.5,205,-1268</points>
<connection>
<GID>5768</GID>
<name>OUT_0</name></connection>
<intersection>-1268 12</intersection></vsegment></shape></wire>
<wire>
<ID>4336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-1399.5,212,-1236.5</points>
<connection>
<GID>6021</GID>
<name>N_in1</name></connection>
<connection>
<GID>6023</GID>
<name>N_in0</name></connection>
<intersection>-1376 11</intersection>
<intersection>-1357.5 10</intersection>
<intersection>-1338.5 9</intersection>
<intersection>-1320 7</intersection>
<intersection>-1298 6</intersection>
<intersection>-1279.5 5</intersection>
<intersection>-1260.5 4</intersection>
<intersection>-1242 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-1242,215,-1242</points>
<connection>
<GID>5806</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>212,-1260.5,215,-1260.5</points>
<connection>
<GID>5770</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>212,-1279.5,215,-1279.5</points>
<connection>
<GID>6097</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>212,-1298,215,-1298</points>
<connection>
<GID>6061</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>212,-1320,215,-1320</points>
<connection>
<GID>5960</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>212,-1338.5,215,-1338.5</points>
<connection>
<GID>5939</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>212,-1357.5,215,-1357.5</points>
<connection>
<GID>5928</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>212,-1376,215,-1376</points>
<connection>
<GID>5910</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>4337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-1399.5,233,-1237.5</points>
<connection>
<GID>6025</GID>
<name>N_in1</name></connection>
<connection>
<GID>5983</GID>
<name>N_in0</name></connection>
<intersection>-1383.5 11</intersection>
<intersection>-1365 10</intersection>
<intersection>-1346 9</intersection>
<intersection>-1327.5 8</intersection>
<intersection>-1305.5 7</intersection>
<intersection>-1287 6</intersection>
<intersection>-1268 5</intersection>
<intersection>-1249.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>228,-1249.5,233,-1249.5</points>
<intersection>228 12</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-1268,233,-1268</points>
<intersection>228 21</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>228,-1287,233,-1287</points>
<intersection>228 20</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>228,-1305.5,233,-1305.5</points>
<intersection>228 19</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>228,-1327.5,233,-1327.5</points>
<intersection>228 16</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>228,-1346,233,-1346</points>
<intersection>228 15</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>228,-1365,233,-1365</points>
<intersection>228 14</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>228,-1383.5,233,-1383.5</points>
<intersection>228 13</intersection>
<intersection>233 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>228,-1252,228,-1249.5</points>
<connection>
<GID>5808</GID>
<name>OUT_0</name></connection>
<intersection>-1249.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>228,-1386,228,-1383.5</points>
<connection>
<GID>5911</GID>
<name>OUT_0</name></connection>
<intersection>-1383.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>228,-1367.5,228,-1365</points>
<connection>
<GID>5929</GID>
<name>OUT_0</name></connection>
<intersection>-1365 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>228,-1348.5,228,-1346</points>
<connection>
<GID>5940</GID>
<name>OUT_0</name></connection>
<intersection>-1346 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>228,-1330,228,-1327.5</points>
<connection>
<GID>5961</GID>
<name>OUT_0</name></connection>
<intersection>-1327.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>228,-1308,228,-1305.5</points>
<connection>
<GID>6063</GID>
<name>OUT_0</name></connection>
<intersection>-1305.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>228,-1289.5,228,-1287</points>
<connection>
<GID>6099</GID>
<name>OUT_0</name></connection>
<intersection>-1287 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>228,-1270.5,228,-1268</points>
<connection>
<GID>5772</GID>
<name>OUT_0</name></connection>
<intersection>-1268 5</intersection></vsegment></shape></wire>
<wire>
<ID>4338</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-117,-1244,22.5,-1244</points>
<connection>
<GID>5774</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-1253.5,-117,-1228</points>
<intersection>-1253.5 4</intersection>
<intersection>-1244 2</intersection>
<intersection>-1228 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-1253.5,34,-1253.5</points>
<connection>
<GID>5776</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-1228,-117,-1228</points>
<connection>
<GID>5907</GID>
<name>OUT_7</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>4339</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-118,-1262.5,22.5,-1262.5</points>
<connection>
<GID>6101</GID>
<name>IN_0</name></connection>
<intersection>-118 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-118,-1272,-118,-1229</points>
<intersection>-1272 5</intersection>
<intersection>-1262.5 2</intersection>
<intersection>-1229 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-118,-1272,34,-1272</points>
<connection>
<GID>6103</GID>
<name>IN_0</name></connection>
<intersection>-118 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-1229,-118,-1229</points>
<connection>
<GID>5907</GID>
<name>OUT_6</name></connection>
<intersection>-118 4</intersection></hsegment></shape></wire>
<wire>
<ID>4340</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-119,-1281.5,22.5,-1281.5</points>
<connection>
<GID>6065</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-1291,-119,-1230</points>
<intersection>-1291 4</intersection>
<intersection>-1281.5 2</intersection>
<intersection>-1230 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-1291,34,-1291</points>
<connection>
<GID>6067</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-1230,-119,-1230</points>
<connection>
<GID>5907</GID>
<name>OUT_5</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>4341</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-120,-1300,22.5,-1300</points>
<connection>
<GID>5985</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-1309.5,-120,-1231</points>
<intersection>-1309.5 4</intersection>
<intersection>-1300 2</intersection>
<intersection>-1231 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-120,-1309.5,34,-1309.5</points>
<connection>
<GID>5987</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1231,-120,-1231</points>
<connection>
<GID>5907</GID>
<name>OUT_4</name></connection>
<intersection>-120 3</intersection></hsegment></shape></wire>
<wire>
<ID>4342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-1322,22.5,-1322</points>
<connection>
<GID>5941</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-1331.5,-121,-1232</points>
<intersection>-1331.5 4</intersection>
<intersection>-1322 1</intersection>
<intersection>-1232 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-1331.5,33.5,-1331.5</points>
<connection>
<GID>5942</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1232,-121,-1232</points>
<connection>
<GID>5907</GID>
<name>OUT_3</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-1340.5,22.5,-1340.5</points>
<connection>
<GID>5930</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-1350,-122,-1233</points>
<intersection>-1350 4</intersection>
<intersection>-1340.5 1</intersection>
<intersection>-1233 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-1350,33.5,-1350</points>
<connection>
<GID>5815</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1233,-122,-1233</points>
<connection>
<GID>5907</GID>
<name>OUT_2</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>4344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123,-1359.5,22.5,-1359.5</points>
<connection>
<GID>5912</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-1369,-123,-1234</points>
<intersection>-1369 4</intersection>
<intersection>-1359.5 1</intersection>
<intersection>-1234 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-1369,33.5,-1369</points>
<connection>
<GID>5913</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-1234,-123,-1234</points>
<connection>
<GID>5907</GID>
<name>OUT_1</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>4345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,-1378,22.5,-1378</points>
<connection>
<GID>5810</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-1387.5,-124,-1235</points>
<connection>
<GID>5907</GID>
<name>OUT_0</name></connection>
<intersection>-1387.5 4</intersection>
<intersection>-1378 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-1387.5,33.5,-1387.5</points>
<connection>
<GID>5812</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>4346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-1401.5,21.5,-1236.5</points>
<connection>
<GID>6043</GID>
<name>N_in1</name></connection>
<connection>
<GID>6035</GID>
<name>N_in0</name></connection>
<intersection>-1380 10</intersection>
<intersection>-1361.5 9</intersection>
<intersection>-1342.5 8</intersection>
<intersection>-1324 7</intersection>
<intersection>-1302 6</intersection>
<intersection>-1283.5 5</intersection>
<intersection>-1264.5 4</intersection>
<intersection>-1246 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-1246,22.5,-1246</points>
<connection>
<GID>5774</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-1264.5,22.5,-1264.5</points>
<connection>
<GID>6101</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>21.5,-1283.5,22.5,-1283.5</points>
<connection>
<GID>6065</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-1302,22.5,-1302</points>
<connection>
<GID>5985</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21.5,-1324,22.5,-1324</points>
<connection>
<GID>5941</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>21.5,-1342.5,22.5,-1342.5</points>
<connection>
<GID>5930</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>21.5,-1361.5,22.5,-1361.5</points>
<connection>
<GID>5912</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>21.5,-1380,22.5,-1380</points>
<connection>
<GID>5810</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-1401.5,31.5,-1236.5</points>
<connection>
<GID>6039</GID>
<name>N_in1</name></connection>
<connection>
<GID>6031</GID>
<name>N_in0</name></connection>
<intersection>-1389.5 3</intersection>
<intersection>-1371 5</intersection>
<intersection>-1352 7</intersection>
<intersection>-1333.5 9</intersection>
<intersection>-1311.5 11</intersection>
<intersection>-1293 13</intersection>
<intersection>-1274 15</intersection>
<intersection>-1255.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-1389.5,33.5,-1389.5</points>
<connection>
<GID>5812</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-1371,33.5,-1371</points>
<connection>
<GID>5913</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31.5,-1352,33.5,-1352</points>
<connection>
<GID>5815</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>31.5,-1333.5,33.5,-1333.5</points>
<connection>
<GID>5942</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>31.5,-1311.5,34,-1311.5</points>
<connection>
<GID>5987</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>31.5,-1293,34,-1293</points>
<connection>
<GID>6067</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>31.5,-1274,34,-1274</points>
<connection>
<GID>6103</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>31.5,-1255.5,34,-1255.5</points>
<connection>
<GID>5776</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-1234.5,21.5,-1228</points>
<connection>
<GID>6035</GID>
<name>N_in1</name></connection>
<connection>
<GID>5905</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-1234.5,31.5,-1228</points>
<connection>
<GID>6031</GID>
<name>N_in1</name></connection>
<connection>
<GID>5904</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-1234.5,44.5,-1228</points>
<connection>
<GID>5962</GID>
<name>N_in1</name></connection>
<connection>
<GID>5885</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-1234,67.5,-1227.5</points>
<connection>
<GID>5963</GID>
<name>N_in1</name></connection>
<connection>
<GID>5886</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-1234.5,70.5,-1227.5</points>
<connection>
<GID>5964</GID>
<name>N_in1</name></connection>
<connection>
<GID>5887</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-1234,90,-1227.5</points>
<connection>
<GID>5965</GID>
<name>N_in1</name></connection>
<connection>
<GID>5888</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-1234,93.5,-1227.5</points>
<connection>
<GID>5966</GID>
<name>N_in1</name></connection>
<connection>
<GID>5889</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-1234.5,114.5,-1227.5</points>
<connection>
<GID>5967</GID>
<name>N_in1</name></connection>
<connection>
<GID>5890</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-1234,118.5,-1227.5</points>
<connection>
<GID>5968</GID>
<name>N_in1</name></connection>
<connection>
<GID>5891</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-1234,137,-1227.5</points>
<connection>
<GID>5969</GID>
<name>N_in1</name></connection>
<connection>
<GID>5892</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-1234,141,-1227.5</points>
<connection>
<GID>5971</GID>
<name>N_in1</name></connection>
<connection>
<GID>5893</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-1234,160,-1227</points>
<connection>
<GID>5973</GID>
<name>N_in1</name></connection>
<connection>
<GID>5894</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-1234,165,-1227</points>
<connection>
<GID>5975</GID>
<name>N_in1</name></connection>
<connection>
<GID>5895</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-1234,183,-1226.5</points>
<connection>
<GID>5979</GID>
<name>N_in1</name></connection>
<connection>
<GID>5896</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-1234,187.5,-1226.5</points>
<connection>
<GID>5977</GID>
<name>N_in1</name></connection>
<connection>
<GID>5897</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-1234.5,208.5,-1226</points>
<connection>
<GID>5981</GID>
<name>N_in1</name></connection>
<connection>
<GID>5898</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-1234.5,212,-1226</points>
<connection>
<GID>6023</GID>
<name>N_in1</name></connection>
<connection>
<GID>5899</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-1235.5,233,-1226</points>
<connection>
<GID>5983</GID>
<name>N_in1</name></connection>
<connection>
<GID>5901</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4366</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1525,61,-1525</points>
<connection>
<GID>6319</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1525,55,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1509.5,55,-1509.5</points>
<connection>
<GID>6313</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4367</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1525,84,-1525</points>
<connection>
<GID>6337</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1525,78,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1509.5,78,-1509.5</points>
<connection>
<GID>6335</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1525,109,-1525</points>
<connection>
<GID>6341</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1525,103,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1509.5,103,-1509.5</points>
<connection>
<GID>6339</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1525,132,-1525</points>
<connection>
<GID>6345</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1525,126,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1509.5,126,-1509.5</points>
<connection>
<GID>6343</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4370</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1525,155,-1525</points>
<connection>
<GID>6349</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1525,149,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1509.5,149,-1509.5</points>
<connection>
<GID>6347</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1525,178,-1525</points>
<connection>
<GID>6353</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1525,172,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1509.5,172,-1509.5</points>
<connection>
<GID>6351</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1525,203,-1525</points>
<connection>
<GID>6357</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1525,197,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1509.5,197,-1509.5</points>
<connection>
<GID>6355</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1525,226,-1525</points>
<connection>
<GID>6361</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1525,220,-1509.5</points>
<intersection>-1525 1</intersection>
<intersection>-1509.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1509.5,220,-1509.5</points>
<connection>
<GID>6359</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1512.5,213,-1512.5</points>
<connection>
<GID>6359</GID>
<name>clock</name></connection>
<connection>
<GID>6355</GID>
<name>clock</name></connection>
<connection>
<GID>6351</GID>
<name>clock</name></connection>
<connection>
<GID>6347</GID>
<name>clock</name></connection>
<connection>
<GID>6343</GID>
<name>clock</name></connection>
<connection>
<GID>6339</GID>
<name>clock</name></connection>
<connection>
<GID>6335</GID>
<name>clock</name></connection>
<connection>
<GID>6313</GID>
<name>clock</name></connection>
<connection>
<GID>6303</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4375</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1522,224,-1522</points>
<connection>
<GID>6361</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6357</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6353</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6349</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6345</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6341</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6337</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6319</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6308</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1506.5,61,-1506.5</points>
<connection>
<GID>6369</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1506.5,55,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1491,55,-1491</points>
<connection>
<GID>6367</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1506.5,84,-1506.5</points>
<connection>
<GID>6373</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1506.5,78,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1491,78,-1491</points>
<connection>
<GID>6371</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4378</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1506.5,109,-1506.5</points>
<connection>
<GID>6377</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1506.5,103,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1491,103,-1491</points>
<connection>
<GID>6375</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4379</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1506.5,132,-1506.5</points>
<connection>
<GID>6381</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1506.5,126,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1491,126,-1491</points>
<connection>
<GID>6379</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1506.5,155,-1506.5</points>
<connection>
<GID>6385</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1506.5,149,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1491,149,-1491</points>
<connection>
<GID>6383</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4381</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1506.5,178,-1506.5</points>
<connection>
<GID>6389</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1506.5,172,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1491,172,-1491</points>
<connection>
<GID>6387</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4382</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1506.5,203,-1506.5</points>
<connection>
<GID>6393</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1506.5,197,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1491,197,-1491</points>
<connection>
<GID>6391</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4383</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1506.5,226,-1506.5</points>
<connection>
<GID>6397</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1506.5,220,-1491</points>
<intersection>-1506.5 1</intersection>
<intersection>-1491 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1491,220,-1491</points>
<connection>
<GID>6395</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4384</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1494,213,-1494</points>
<connection>
<GID>6395</GID>
<name>clock</name></connection>
<connection>
<GID>6391</GID>
<name>clock</name></connection>
<connection>
<GID>6387</GID>
<name>clock</name></connection>
<connection>
<GID>6383</GID>
<name>clock</name></connection>
<connection>
<GID>6379</GID>
<name>clock</name></connection>
<connection>
<GID>6375</GID>
<name>clock</name></connection>
<connection>
<GID>6371</GID>
<name>clock</name></connection>
<connection>
<GID>6367</GID>
<name>clock</name></connection>
<connection>
<GID>6363</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1503.5,224,-1503.5</points>
<connection>
<GID>6397</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6393</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6389</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6385</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6381</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6377</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6373</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6369</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6365</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1487.5,61,-1487.5</points>
<connection>
<GID>6405</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1487.5,55,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1472,55,-1472</points>
<connection>
<GID>6403</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4387</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1487.5,84,-1487.5</points>
<connection>
<GID>6409</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1487.5,78,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1472,78,-1472</points>
<connection>
<GID>6407</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1487.5,109,-1487.5</points>
<connection>
<GID>6413</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1487.5,103,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1472,103,-1472</points>
<connection>
<GID>6411</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1487.5,132,-1487.5</points>
<connection>
<GID>6417</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1487.5,126,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1472,126,-1472</points>
<connection>
<GID>6415</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4390</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1487.5,155,-1487.5</points>
<connection>
<GID>6421</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1487.5,149,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1472,149,-1472</points>
<connection>
<GID>6419</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4391</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1487.5,178,-1487.5</points>
<connection>
<GID>6425</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1487.5,172,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1472,172,-1472</points>
<connection>
<GID>6423</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1487.5,203,-1487.5</points>
<connection>
<GID>6429</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1487.5,197,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1472,197,-1472</points>
<connection>
<GID>6427</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4393</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1487.5,226,-1487.5</points>
<connection>
<GID>6433</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1487.5,220,-1472</points>
<intersection>-1487.5 1</intersection>
<intersection>-1472 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1472,220,-1472</points>
<connection>
<GID>6431</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1475,213,-1475</points>
<connection>
<GID>6431</GID>
<name>clock</name></connection>
<connection>
<GID>6427</GID>
<name>clock</name></connection>
<connection>
<GID>6423</GID>
<name>clock</name></connection>
<connection>
<GID>6419</GID>
<name>clock</name></connection>
<connection>
<GID>6415</GID>
<name>clock</name></connection>
<connection>
<GID>6411</GID>
<name>clock</name></connection>
<connection>
<GID>6407</GID>
<name>clock</name></connection>
<connection>
<GID>6403</GID>
<name>clock</name></connection>
<connection>
<GID>6399</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4395</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1484.5,224,-1484.5</points>
<connection>
<GID>6433</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6429</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6425</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6421</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6417</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6413</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6409</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6405</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6401</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1469,61,-1469</points>
<connection>
<GID>6441</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1469,55,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1453.5,55,-1453.5</points>
<connection>
<GID>6439</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1469,84,-1469</points>
<connection>
<GID>6445</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1469,78,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1453.5,78,-1453.5</points>
<connection>
<GID>6443</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4398</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1469,109,-1469</points>
<connection>
<GID>6449</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1469,103,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1453.5,103,-1453.5</points>
<connection>
<GID>6447</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1469,132,-1469</points>
<connection>
<GID>6453</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1469,126,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1453.5,126,-1453.5</points>
<connection>
<GID>6451</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4400</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1469,155,-1469</points>
<connection>
<GID>6457</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1469,149,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1453.5,149,-1453.5</points>
<connection>
<GID>6455</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1469,178,-1469</points>
<connection>
<GID>6461</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1469,172,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1453.5,172,-1453.5</points>
<connection>
<GID>6459</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1469,203,-1469</points>
<connection>
<GID>6465</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1469,197,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1453.5,197,-1453.5</points>
<connection>
<GID>6463</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1469,226,-1469</points>
<connection>
<GID>6469</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1469,220,-1453.5</points>
<intersection>-1469 1</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1453.5,220,-1453.5</points>
<connection>
<GID>6467</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4404</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1456.5,213,-1456.5</points>
<connection>
<GID>6467</GID>
<name>clock</name></connection>
<connection>
<GID>6463</GID>
<name>clock</name></connection>
<connection>
<GID>6459</GID>
<name>clock</name></connection>
<connection>
<GID>6455</GID>
<name>clock</name></connection>
<connection>
<GID>6451</GID>
<name>clock</name></connection>
<connection>
<GID>6447</GID>
<name>clock</name></connection>
<connection>
<GID>6443</GID>
<name>clock</name></connection>
<connection>
<GID>6439</GID>
<name>clock</name></connection>
<connection>
<GID>6435</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1466,224,-1466</points>
<connection>
<GID>6469</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6465</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6461</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6457</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6453</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6449</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6445</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6441</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6437</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1603,61,-1603</points>
<connection>
<GID>6477</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1603,55,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1587.5,55,-1587.5</points>
<connection>
<GID>6475</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4407</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1603,84,-1603</points>
<connection>
<GID>6481</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1603,78,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1587.5,78,-1587.5</points>
<connection>
<GID>6479</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4408</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1603,109,-1603</points>
<connection>
<GID>6485</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1603,103,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1587.5,103,-1587.5</points>
<connection>
<GID>6483</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1603,132,-1603</points>
<connection>
<GID>6126</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1603,126,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1587.5,126,-1587.5</points>
<connection>
<GID>6124</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4410</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1603,155,-1603</points>
<connection>
<GID>6130</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1603,149,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1587.5,149,-1587.5</points>
<connection>
<GID>6128</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1603,178,-1603</points>
<connection>
<GID>6134</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1603,172,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1587.5,172,-1587.5</points>
<connection>
<GID>6132</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1603,203,-1603</points>
<connection>
<GID>6138</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1603,197,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1587.5,197,-1587.5</points>
<connection>
<GID>6136</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1603,226,-1603</points>
<connection>
<GID>6142</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1603,220,-1587.5</points>
<intersection>-1603 1</intersection>
<intersection>-1587.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1587.5,220,-1587.5</points>
<connection>
<GID>6140</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1590.5,213,-1590.5</points>
<connection>
<GID>6140</GID>
<name>clock</name></connection>
<connection>
<GID>6136</GID>
<name>clock</name></connection>
<connection>
<GID>6132</GID>
<name>clock</name></connection>
<connection>
<GID>6128</GID>
<name>clock</name></connection>
<connection>
<GID>6124</GID>
<name>clock</name></connection>
<connection>
<GID>6483</GID>
<name>clock</name></connection>
<connection>
<GID>6479</GID>
<name>clock</name></connection>
<connection>
<GID>6475</GID>
<name>clock</name></connection>
<connection>
<GID>6471</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1600,224,-1600</points>
<connection>
<GID>6142</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6138</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6134</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6130</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6126</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6485</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6481</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6477</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6473</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1584.5,61,-1584.5</points>
<connection>
<GID>6150</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1584.5,55,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1569,55,-1569</points>
<connection>
<GID>6148</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1584.5,84,-1584.5</points>
<connection>
<GID>6154</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1584.5,78,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1569,78,-1569</points>
<connection>
<GID>6152</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4418</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1584.5,109,-1584.5</points>
<connection>
<GID>6158</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1584.5,103,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1569,103,-1569</points>
<connection>
<GID>6156</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1584.5,132,-1584.5</points>
<connection>
<GID>6162</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1584.5,126,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1569,126,-1569</points>
<connection>
<GID>6160</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1584.5,155,-1584.5</points>
<connection>
<GID>6166</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1584.5,149,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1569,149,-1569</points>
<connection>
<GID>6164</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1584.5,178,-1584.5</points>
<connection>
<GID>6170</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1584.5,172,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1569,172,-1569</points>
<connection>
<GID>6168</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1584.5,203,-1584.5</points>
<connection>
<GID>6174</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1584.5,197,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1569,197,-1569</points>
<connection>
<GID>6172</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1584.5,226,-1584.5</points>
<connection>
<GID>6178</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1584.5,220,-1569</points>
<intersection>-1584.5 1</intersection>
<intersection>-1569 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1569,220,-1569</points>
<connection>
<GID>6176</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1572,213,-1572</points>
<connection>
<GID>6156</GID>
<name>clock</name></connection>
<connection>
<GID>6152</GID>
<name>clock</name></connection>
<connection>
<GID>6148</GID>
<name>clock</name></connection>
<connection>
<GID>6144</GID>
<name>OUT</name></connection>
<connection>
<GID>6176</GID>
<name>clock</name></connection>
<connection>
<GID>6172</GID>
<name>clock</name></connection>
<connection>
<GID>6168</GID>
<name>clock</name></connection>
<connection>
<GID>6164</GID>
<name>clock</name></connection>
<connection>
<GID>6160</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1581.5,224,-1581.5</points>
<connection>
<GID>6154</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6150</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6146</GID>
<name>OUT</name></connection>
<connection>
<GID>6178</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6174</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6170</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6166</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6162</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6158</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1565.5,61,-1565.5</points>
<connection>
<GID>6188</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1565.5,55,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1550,55,-1550</points>
<connection>
<GID>6186</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1565.5,84,-1565.5</points>
<connection>
<GID>6193</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1565.5,78,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1550,78,-1550</points>
<connection>
<GID>6191</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1565.5,109,-1565.5</points>
<connection>
<GID>6198</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1565.5,103,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1550,103,-1550</points>
<connection>
<GID>6196</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4429</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1565.5,132,-1565.5</points>
<connection>
<GID>6203</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1565.5,126,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1550,126,-1550</points>
<connection>
<GID>6201</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1565.5,155,-1565.5</points>
<connection>
<GID>6208</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1565.5,149,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1550,149,-1550</points>
<connection>
<GID>6206</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4431</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1565.5,178,-1565.5</points>
<connection>
<GID>6211</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1565.5,172,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1550,172,-1550</points>
<connection>
<GID>6210</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4432</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1565.5,203,-1565.5</points>
<connection>
<GID>6214</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1565.5,197,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1550,197,-1550</points>
<connection>
<GID>6213</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4433</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1565.5,226,-1565.5</points>
<connection>
<GID>6216</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1565.5,220,-1550</points>
<intersection>-1565.5 1</intersection>
<intersection>-1550 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1550,220,-1550</points>
<connection>
<GID>6215</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1553,213,-1553</points>
<connection>
<GID>6215</GID>
<name>clock</name></connection>
<connection>
<GID>6213</GID>
<name>clock</name></connection>
<connection>
<GID>6210</GID>
<name>clock</name></connection>
<connection>
<GID>6206</GID>
<name>clock</name></connection>
<connection>
<GID>6201</GID>
<name>clock</name></connection>
<connection>
<GID>6196</GID>
<name>clock</name></connection>
<connection>
<GID>6191</GID>
<name>clock</name></connection>
<connection>
<GID>6186</GID>
<name>clock</name></connection>
<connection>
<GID>6181</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1562.5,224,-1562.5</points>
<connection>
<GID>6216</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6214</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6211</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6208</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6203</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6198</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6193</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6188</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6183</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1547,61,-1547</points>
<connection>
<GID>6220</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1547,55,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1531.5,55,-1531.5</points>
<connection>
<GID>6219</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4437</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1547,84,-1547</points>
<connection>
<GID>6222</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1547,78,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1531.5,78,-1531.5</points>
<connection>
<GID>6221</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1547,109,-1547</points>
<connection>
<GID>6224</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1547,103,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1531.5,103,-1531.5</points>
<connection>
<GID>6223</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4439</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1547,132,-1547</points>
<connection>
<GID>6226</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1547,126,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1531.5,126,-1531.5</points>
<connection>
<GID>6225</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4440</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1547,155,-1547</points>
<connection>
<GID>6228</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1547,149,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1531.5,149,-1531.5</points>
<connection>
<GID>6227</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4441</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1547,178,-1547</points>
<connection>
<GID>6230</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1547,172,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1531.5,172,-1531.5</points>
<connection>
<GID>6229</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4442</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1547,203,-1547</points>
<connection>
<GID>6232</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1547,197,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1531.5,197,-1531.5</points>
<connection>
<GID>6231</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1547,226,-1547</points>
<connection>
<GID>6234</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1547,220,-1531.5</points>
<intersection>-1547 1</intersection>
<intersection>-1531.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1531.5,220,-1531.5</points>
<connection>
<GID>6233</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4444</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1534.5,213,-1534.5</points>
<connection>
<GID>6233</GID>
<name>clock</name></connection>
<connection>
<GID>6231</GID>
<name>clock</name></connection>
<connection>
<GID>6229</GID>
<name>clock</name></connection>
<connection>
<GID>6227</GID>
<name>clock</name></connection>
<connection>
<GID>6225</GID>
<name>clock</name></connection>
<connection>
<GID>6223</GID>
<name>clock</name></connection>
<connection>
<GID>6221</GID>
<name>clock</name></connection>
<connection>
<GID>6219</GID>
<name>clock</name></connection>
<connection>
<GID>6217</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4445</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1544,224,-1544</points>
<connection>
<GID>6234</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6232</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6230</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6228</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6226</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6224</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6222</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6220</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6218</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-1613,42.5,-1448</points>
<connection>
<GID>6250</GID>
<name>N_in1</name></connection>
<connection>
<GID>6235</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 12</intersection>
<intersection>-1569 11</intersection>
<intersection>-1550 10</intersection>
<intersection>-1531.5 9</intersection>
<intersection>-1509.5 8</intersection>
<intersection>-1491 7</intersection>
<intersection>-1472 6</intersection>
<intersection>-1453.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-1453.5,48,-1453.5</points>
<connection>
<GID>6439</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>42.5,-1472,48,-1472</points>
<connection>
<GID>6403</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>42.5,-1491,48,-1491</points>
<connection>
<GID>6367</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>42.5,-1509.5,48,-1509.5</points>
<connection>
<GID>6313</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42.5,-1531.5,48,-1531.5</points>
<connection>
<GID>6219</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>42.5,-1550,48,-1550</points>
<connection>
<GID>6186</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>42.5,-1569,48,-1569</points>
<connection>
<GID>6148</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>42.5,-1587.5,48,-1587.5</points>
<connection>
<GID>6475</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-1612.5,65.5,-1447.5</points>
<connection>
<GID>6251</GID>
<name>N_in1</name></connection>
<connection>
<GID>6236</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 4</intersection>
<intersection>-1579 5</intersection>
<intersection>-1560 6</intersection>
<intersection>-1541.5 7</intersection>
<intersection>-1519.5 8</intersection>
<intersection>-1501 9</intersection>
<intersection>-1482 10</intersection>
<intersection>-1463.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>61,-1597.5,65.5,-1597.5</points>
<connection>
<GID>6477</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-1579,65.5,-1579</points>
<connection>
<GID>6150</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61,-1560,65.5,-1560</points>
<connection>
<GID>6188</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61,-1541.5,65.5,-1541.5</points>
<connection>
<GID>6220</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61,-1519.5,65.5,-1519.5</points>
<connection>
<GID>6319</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61,-1501,65.5,-1501</points>
<connection>
<GID>6369</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61,-1482,65.5,-1482</points>
<connection>
<GID>6405</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>61,-1463.5,65.5,-1463.5</points>
<connection>
<GID>6441</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-1612.5,68.5,-1448</points>
<connection>
<GID>6252</GID>
<name>N_in1</name></connection>
<connection>
<GID>6237</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 10</intersection>
<intersection>-1569 9</intersection>
<intersection>-1550 8</intersection>
<intersection>-1531.5 7</intersection>
<intersection>-1509.5 6</intersection>
<intersection>-1491 5</intersection>
<intersection>-1472 4</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>68.5,-1453.5,71,-1453.5</points>
<connection>
<GID>6443</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-1472,71,-1472</points>
<connection>
<GID>6407</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68.5,-1491,71,-1491</points>
<connection>
<GID>6371</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68.5,-1509.5,71,-1509.5</points>
<connection>
<GID>6335</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68.5,-1531.5,71,-1531.5</points>
<connection>
<GID>6221</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-1550,71,-1550</points>
<connection>
<GID>6191</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68.5,-1569,71,-1569</points>
<connection>
<GID>6152</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68.5,-1587.5,71,-1587.5</points>
<connection>
<GID>6479</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-1612.5,88,-1447.5</points>
<connection>
<GID>6253</GID>
<name>N_in1</name></connection>
<connection>
<GID>6238</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 6</intersection>
<intersection>-1579 7</intersection>
<intersection>-1560 8</intersection>
<intersection>-1541.5 9</intersection>
<intersection>-1519.5 10</intersection>
<intersection>-1501 11</intersection>
<intersection>-1482 12</intersection>
<intersection>-1463.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84,-1597.5,88,-1597.5</points>
<connection>
<GID>6481</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84,-1579,88,-1579</points>
<connection>
<GID>6154</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>84,-1560,88,-1560</points>
<connection>
<GID>6193</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84,-1541.5,88,-1541.5</points>
<connection>
<GID>6222</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84,-1519.5,88,-1519.5</points>
<connection>
<GID>6337</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84,-1501,88,-1501</points>
<connection>
<GID>6373</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>84,-1482,88,-1482</points>
<connection>
<GID>6409</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>84,-1463.5,88,-1463.5</points>
<connection>
<GID>6445</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>4450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-1612.5,91.5,-1447.5</points>
<connection>
<GID>6254</GID>
<name>N_in1</name></connection>
<connection>
<GID>6239</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 13</intersection>
<intersection>-1569 12</intersection>
<intersection>-1550 11</intersection>
<intersection>-1531.5 10</intersection>
<intersection>-1509.5 9</intersection>
<intersection>-1491 8</intersection>
<intersection>-1472 7</intersection>
<intersection>-1453.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91.5,-1453.5,96,-1453.5</points>
<connection>
<GID>6447</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>91.5,-1472,96,-1472</points>
<connection>
<GID>6411</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>91.5,-1491,96,-1491</points>
<connection>
<GID>6375</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>91.5,-1509.5,96,-1509.5</points>
<connection>
<GID>6339</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>91.5,-1531.5,96,-1531.5</points>
<connection>
<GID>6223</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>91.5,-1550,96,-1550</points>
<connection>
<GID>6196</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>91.5,-1569,96,-1569</points>
<connection>
<GID>6156</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>91.5,-1587.5,96,-1587.5</points>
<connection>
<GID>6483</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-1612.5,112.5,-1448</points>
<connection>
<GID>6255</GID>
<name>N_in1</name></connection>
<connection>
<GID>6240</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 6</intersection>
<intersection>-1579 7</intersection>
<intersection>-1560 8</intersection>
<intersection>-1541.5 9</intersection>
<intersection>-1519.5 10</intersection>
<intersection>-1501 11</intersection>
<intersection>-1482 12</intersection>
<intersection>-1463.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109,-1597.5,112.5,-1597.5</points>
<connection>
<GID>6485</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>109,-1579,112.5,-1579</points>
<connection>
<GID>6158</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109,-1560,112.5,-1560</points>
<connection>
<GID>6198</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>109,-1541.5,112.5,-1541.5</points>
<connection>
<GID>6224</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>109,-1519.5,112.5,-1519.5</points>
<connection>
<GID>6341</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>109,-1501,112.5,-1501</points>
<connection>
<GID>6377</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109,-1482,112.5,-1482</points>
<connection>
<GID>6413</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>109,-1463.5,112.5,-1463.5</points>
<connection>
<GID>6449</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-1612.5,116.5,-1447.5</points>
<connection>
<GID>6256</GID>
<name>N_in1</name></connection>
<connection>
<GID>6241</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 13</intersection>
<intersection>-1569 12</intersection>
<intersection>-1550 11</intersection>
<intersection>-1531.5 10</intersection>
<intersection>-1509.5 9</intersection>
<intersection>-1491 8</intersection>
<intersection>-1472 7</intersection>
<intersection>-1453.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116.5,-1453.5,119,-1453.5</points>
<connection>
<GID>6451</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116.5,-1472,119,-1472</points>
<connection>
<GID>6415</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>116.5,-1491,119,-1491</points>
<connection>
<GID>6379</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116.5,-1509.5,119,-1509.5</points>
<connection>
<GID>6343</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116.5,-1531.5,119,-1531.5</points>
<connection>
<GID>6225</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>116.5,-1550,119,-1550</points>
<connection>
<GID>6201</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>116.5,-1569,119,-1569</points>
<connection>
<GID>6160</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>116.5,-1587.5,119,-1587.5</points>
<connection>
<GID>6124</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-1612.5,135,-1447.5</points>
<connection>
<GID>6257</GID>
<name>N_in1</name></connection>
<connection>
<GID>6242</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 6</intersection>
<intersection>-1579 7</intersection>
<intersection>-1560 8</intersection>
<intersection>-1541.5 9</intersection>
<intersection>-1519.5 10</intersection>
<intersection>-1501 11</intersection>
<intersection>-1482 12</intersection>
<intersection>-1463.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>132,-1597.5,135,-1597.5</points>
<connection>
<GID>6126</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>132,-1579,135,-1579</points>
<connection>
<GID>6162</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>132,-1560,135,-1560</points>
<connection>
<GID>6203</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>132,-1541.5,135,-1541.5</points>
<connection>
<GID>6226</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132,-1519.5,135,-1519.5</points>
<connection>
<GID>6345</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132,-1501,135,-1501</points>
<connection>
<GID>6381</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>132,-1482,135,-1482</points>
<connection>
<GID>6417</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132,-1463.5,135,-1463.5</points>
<connection>
<GID>6453</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>4454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-1612.5,139,-1447.5</points>
<connection>
<GID>6258</GID>
<name>N_in1</name></connection>
<connection>
<GID>6243</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 13</intersection>
<intersection>-1569 12</intersection>
<intersection>-1550 11</intersection>
<intersection>-1531.5 10</intersection>
<intersection>-1509.5 9</intersection>
<intersection>-1491 8</intersection>
<intersection>-1472 7</intersection>
<intersection>-1453.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-1453.5,142,-1453.5</points>
<connection>
<GID>6455</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,-1472,142,-1472</points>
<connection>
<GID>6419</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>139,-1491,142,-1491</points>
<connection>
<GID>6383</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>139,-1509.5,142,-1509.5</points>
<connection>
<GID>6347</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>139,-1531.5,142,-1531.5</points>
<connection>
<GID>6227</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139,-1550,142,-1550</points>
<connection>
<GID>6206</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>139,-1569,142,-1569</points>
<connection>
<GID>6164</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>139,-1587.5,142,-1587.5</points>
<connection>
<GID>6128</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>4455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-1612,158,-1447.5</points>
<connection>
<GID>6259</GID>
<name>N_in1</name></connection>
<connection>
<GID>6244</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 6</intersection>
<intersection>-1579 7</intersection>
<intersection>-1560 8</intersection>
<intersection>-1541.5 9</intersection>
<intersection>-1519.5 10</intersection>
<intersection>-1501 11</intersection>
<intersection>-1482 12</intersection>
<intersection>-1463.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>155,-1597.5,158,-1597.5</points>
<connection>
<GID>6130</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>155,-1579,158,-1579</points>
<connection>
<GID>6166</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>155,-1560,158,-1560</points>
<connection>
<GID>6208</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>155,-1541.5,158,-1541.5</points>
<connection>
<GID>6228</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>155,-1519.5,158,-1519.5</points>
<connection>
<GID>6349</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>155,-1501,158,-1501</points>
<connection>
<GID>6385</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>155,-1482,158,-1482</points>
<connection>
<GID>6421</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>155,-1463.5,158,-1463.5</points>
<connection>
<GID>6457</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>4456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-1612,163,-1447.5</points>
<connection>
<GID>6260</GID>
<name>N_in1</name></connection>
<connection>
<GID>6245</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 13</intersection>
<intersection>-1569 12</intersection>
<intersection>-1550 11</intersection>
<intersection>-1531.5 10</intersection>
<intersection>-1509.5 9</intersection>
<intersection>-1491 8</intersection>
<intersection>-1472 7</intersection>
<intersection>-1453.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>163,-1453.5,165,-1453.5</points>
<connection>
<GID>6459</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>163,-1472,165,-1472</points>
<connection>
<GID>6423</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>163,-1491,165,-1491</points>
<connection>
<GID>6387</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>163,-1509.5,165,-1509.5</points>
<connection>
<GID>6351</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>163,-1531.5,165,-1531.5</points>
<connection>
<GID>6229</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>163,-1550,165,-1550</points>
<connection>
<GID>6210</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>163,-1569,165,-1569</points>
<connection>
<GID>6168</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>163,-1587.5,165,-1587.5</points>
<connection>
<GID>6132</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>4457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-1611.5,181,-1447.5</points>
<connection>
<GID>6261</GID>
<name>N_in1</name></connection>
<connection>
<GID>6247</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 16</intersection>
<intersection>-1579 15</intersection>
<intersection>-1560 14</intersection>
<intersection>-1541.5 13</intersection>
<intersection>-1519.5 12</intersection>
<intersection>-1501 11</intersection>
<intersection>-1482 10</intersection>
<intersection>-1463.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>178,-1463.5,181,-1463.5</points>
<connection>
<GID>6461</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>178,-1482,181,-1482</points>
<connection>
<GID>6425</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>178,-1501,181,-1501</points>
<connection>
<GID>6389</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>178,-1519.5,181,-1519.5</points>
<connection>
<GID>6353</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>178,-1541.5,181,-1541.5</points>
<connection>
<GID>6230</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>178,-1560,181,-1560</points>
<connection>
<GID>6211</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>178,-1579,181,-1579</points>
<connection>
<GID>6170</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>178,-1597.5,181,-1597.5</points>
<connection>
<GID>6134</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>4458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-1611.5,185.5,-1447.5</points>
<connection>
<GID>6262</GID>
<name>N_in1</name></connection>
<connection>
<GID>6246</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 13</intersection>
<intersection>-1569 12</intersection>
<intersection>-1550 11</intersection>
<intersection>-1531.5 10</intersection>
<intersection>-1509.5 9</intersection>
<intersection>-1491 8</intersection>
<intersection>-1472 7</intersection>
<intersection>-1453.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>185.5,-1453.5,190,-1453.5</points>
<connection>
<GID>6463</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>185.5,-1472,190,-1472</points>
<connection>
<GID>6427</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>185.5,-1491,190,-1491</points>
<connection>
<GID>6391</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185.5,-1509.5,190,-1509.5</points>
<connection>
<GID>6355</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>185.5,-1531.5,190,-1531.5</points>
<connection>
<GID>6231</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>185.5,-1550,190,-1550</points>
<connection>
<GID>6213</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185.5,-1569,190,-1569</points>
<connection>
<GID>6172</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>185.5,-1587.5,190,-1587.5</points>
<connection>
<GID>6136</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-1611,206.5,-1448</points>
<connection>
<GID>6263</GID>
<name>N_in1</name></connection>
<connection>
<GID>6248</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 6</intersection>
<intersection>-1579 7</intersection>
<intersection>-1560 8</intersection>
<intersection>-1541.5 9</intersection>
<intersection>-1519.5 10</intersection>
<intersection>-1501 11</intersection>
<intersection>-1482 12</intersection>
<intersection>-1463.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>203,-1597.5,206.5,-1597.5</points>
<connection>
<GID>6138</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-1579,206.5,-1579</points>
<connection>
<GID>6174</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>203,-1560,206.5,-1560</points>
<connection>
<GID>6214</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>203,-1541.5,206.5,-1541.5</points>
<connection>
<GID>6232</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>203,-1519.5,206.5,-1519.5</points>
<connection>
<GID>6357</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-1501,206.5,-1501</points>
<connection>
<GID>6393</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>203,-1482,206.5,-1482</points>
<connection>
<GID>6429</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>203,-1463.5,206.5,-1463.5</points>
<connection>
<GID>6465</GID>
<name>OUT_0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-1611,210,-1448</points>
<connection>
<GID>6264</GID>
<name>N_in1</name></connection>
<connection>
<GID>6265</GID>
<name>N_in0</name></connection>
<intersection>-1587.5 11</intersection>
<intersection>-1569 10</intersection>
<intersection>-1550 9</intersection>
<intersection>-1531.5 7</intersection>
<intersection>-1509.5 6</intersection>
<intersection>-1491 5</intersection>
<intersection>-1472 4</intersection>
<intersection>-1453.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>210,-1453.5,213,-1453.5</points>
<connection>
<GID>6467</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>210,-1472,213,-1472</points>
<connection>
<GID>6431</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>210,-1491,213,-1491</points>
<connection>
<GID>6395</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>210,-1509.5,213,-1509.5</points>
<connection>
<GID>6359</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>210,-1531.5,213,-1531.5</points>
<connection>
<GID>6233</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>210,-1550,213,-1550</points>
<connection>
<GID>6215</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210,-1569,213,-1569</points>
<connection>
<GID>6176</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>210,-1587.5,213,-1587.5</points>
<connection>
<GID>6140</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>4461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,-1611,231,-1449</points>
<connection>
<GID>6266</GID>
<name>N_in1</name></connection>
<connection>
<GID>6249</GID>
<name>N_in0</name></connection>
<intersection>-1597.5 11</intersection>
<intersection>-1579 10</intersection>
<intersection>-1560 9</intersection>
<intersection>-1541.5 8</intersection>
<intersection>-1519.5 7</intersection>
<intersection>-1501 6</intersection>
<intersection>-1482 5</intersection>
<intersection>-1463.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>226,-1463.5,231,-1463.5</points>
<connection>
<GID>6469</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>226,-1482,231,-1482</points>
<connection>
<GID>6433</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>226,-1501,231,-1501</points>
<connection>
<GID>6397</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>226,-1519.5,231,-1519.5</points>
<connection>
<GID>6361</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>226,-1541.5,231,-1541.5</points>
<connection>
<GID>6234</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>226,-1560,231,-1560</points>
<connection>
<GID>6216</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>226,-1579,231,-1579</points>
<connection>
<GID>6178</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>226,-1597.5,231,-1597.5</points>
<connection>
<GID>6142</GID>
<name>OUT_0</name></connection>
<intersection>231 0</intersection></hsegment></shape></wire>
<wire>
<ID>4462</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-126,-1455.5,20.5,-1455.5</points>
<connection>
<GID>6435</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-1607,-126,-1455.5</points>
<connection>
<GID>6272</GID>
<name>OUT_15</name></connection>
<intersection>-1465 4</intersection>
<intersection>-1455.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-1465,32,-1465</points>
<connection>
<GID>6437</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>4463</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-125,-1474,20.5,-1474</points>
<connection>
<GID>6399</GID>
<name>IN_0</name></connection>
<intersection>-125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-125,-1608,-125,-1474</points>
<intersection>-1608 6</intersection>
<intersection>-1483.5 5</intersection>
<intersection>-1474 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-125,-1483.5,32,-1483.5</points>
<connection>
<GID>6401</GID>
<name>IN_0</name></connection>
<intersection>-125 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-126,-1608,-125,-1608</points>
<connection>
<GID>6272</GID>
<name>OUT_14</name></connection>
<intersection>-125 4</intersection></hsegment></shape></wire>
<wire>
<ID>4464</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-124,-1493,20.5,-1493</points>
<connection>
<GID>6363</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-1609,-124,-1493</points>
<intersection>-1609 6</intersection>
<intersection>-1502.5 4</intersection>
<intersection>-1493 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-1502.5,32,-1502.5</points>
<connection>
<GID>6365</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-126,-1609,-124,-1609</points>
<connection>
<GID>6272</GID>
<name>OUT_13</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>4465</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-123,-1511.5,20.5,-1511.5</points>
<connection>
<GID>6303</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-1610,-123,-1511.5</points>
<intersection>-1610 5</intersection>
<intersection>-1521 4</intersection>
<intersection>-1511.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-1521,32,-1521</points>
<connection>
<GID>6308</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1610,-123,-1610</points>
<connection>
<GID>6272</GID>
<name>OUT_12</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>4466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-1533.5,20.5,-1533.5</points>
<connection>
<GID>6217</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-1611,-122,-1533.5</points>
<intersection>-1611 6</intersection>
<intersection>-1543 4</intersection>
<intersection>-1533.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-1543,31.5,-1543</points>
<connection>
<GID>6218</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-126,-1611,-122,-1611</points>
<connection>
<GID>6272</GID>
<name>OUT_11</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>4467</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-1552,20.5,-1552</points>
<connection>
<GID>6181</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-1612,-121,-1552</points>
<intersection>-1612 5</intersection>
<intersection>-1561.5 4</intersection>
<intersection>-1552 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-1561.5,31.5,-1561.5</points>
<connection>
<GID>6183</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1612,-121,-1612</points>
<connection>
<GID>6272</GID>
<name>OUT_10</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4468</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-1571,20.5,-1571</points>
<connection>
<GID>6144</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-1613,-120,-1571</points>
<intersection>-1613 5</intersection>
<intersection>-1580.5 4</intersection>
<intersection>-1571 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-120,-1580.5,31.5,-1580.5</points>
<connection>
<GID>6146</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1613,-120,-1613</points>
<connection>
<GID>6272</GID>
<name>OUT_9</name></connection>
<intersection>-120 3</intersection></hsegment></shape></wire>
<wire>
<ID>4469</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,-1589.5,20.5,-1589.5</points>
<connection>
<GID>6471</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-1614,-119,-1589.5</points>
<intersection>-1614 5</intersection>
<intersection>-1599 4</intersection>
<intersection>-1589.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-1599,31.5,-1599</points>
<connection>
<GID>6473</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1614,-119,-1614</points>
<connection>
<GID>6272</GID>
<name>OUT_8</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>4470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-1613,19.5,-1448</points>
<connection>
<GID>6270</GID>
<name>N_in1</name></connection>
<connection>
<GID>6268</GID>
<name>N_in0</name></connection>
<intersection>-1591.5 10</intersection>
<intersection>-1573 9</intersection>
<intersection>-1554 8</intersection>
<intersection>-1535.5 7</intersection>
<intersection>-1513.5 6</intersection>
<intersection>-1495 5</intersection>
<intersection>-1476 4</intersection>
<intersection>-1457.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>19.5,-1457.5,20.5,-1457.5</points>
<connection>
<GID>6435</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>19.5,-1476,20.5,-1476</points>
<connection>
<GID>6399</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>19.5,-1495,20.5,-1495</points>
<connection>
<GID>6363</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>19.5,-1513.5,20.5,-1513.5</points>
<connection>
<GID>6303</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>19.5,-1535.5,20.5,-1535.5</points>
<connection>
<GID>6217</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>19.5,-1554,20.5,-1554</points>
<connection>
<GID>6181</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>19.5,-1573,20.5,-1573</points>
<connection>
<GID>6144</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>19.5,-1591.5,20.5,-1591.5</points>
<connection>
<GID>6471</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-1613,29.5,-1448</points>
<connection>
<GID>6269</GID>
<name>N_in1</name></connection>
<connection>
<GID>6267</GID>
<name>N_in0</name></connection>
<intersection>-1601 3</intersection>
<intersection>-1582.5 5</intersection>
<intersection>-1563.5 7</intersection>
<intersection>-1545 9</intersection>
<intersection>-1523 11</intersection>
<intersection>-1504.5 13</intersection>
<intersection>-1485.5 15</intersection>
<intersection>-1467 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-1601,31.5,-1601</points>
<connection>
<GID>6473</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>29.5,-1582.5,31.5,-1582.5</points>
<connection>
<GID>6146</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>29.5,-1563.5,31.5,-1563.5</points>
<connection>
<GID>6183</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>29.5,-1545,31.5,-1545</points>
<connection>
<GID>6218</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>29.5,-1523,32,-1523</points>
<connection>
<GID>6308</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>29.5,-1504.5,32,-1504.5</points>
<connection>
<GID>6365</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>29.5,-1485.5,32,-1485.5</points>
<connection>
<GID>6401</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>29.5,-1467,32,-1467</points>
<connection>
<GID>6437</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1700.5,61,-1700.5</points>
<connection>
<GID>6368</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1700.5,55,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1685,55,-1685</points>
<connection>
<GID>6356</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4473</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1700.5,84,-1700.5</points>
<connection>
<GID>6394</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1700.5,78,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1685,78,-1685</points>
<connection>
<GID>6392</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1700.5,109,-1700.5</points>
<connection>
<GID>6402</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1700.5,103,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1685,103,-1685</points>
<connection>
<GID>6398</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4475</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1700.5,132,-1700.5</points>
<connection>
<GID>6410</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1700.5,126,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1685,126,-1685</points>
<connection>
<GID>6406</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4476</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1700.5,155,-1700.5</points>
<connection>
<GID>6416</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1700.5,149,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1685,149,-1685</points>
<connection>
<GID>6412</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4477</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1700.5,178,-1700.5</points>
<connection>
<GID>6420</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1700.5,172,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1685,172,-1685</points>
<connection>
<GID>6418</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1700.5,203,-1700.5</points>
<connection>
<GID>6424</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1700.5,197,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1685,197,-1685</points>
<connection>
<GID>6422</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4479</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1700.5,226,-1700.5</points>
<connection>
<GID>6428</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1700.5,220,-1685</points>
<intersection>-1700.5 1</intersection>
<intersection>-1685 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1685,220,-1685</points>
<connection>
<GID>6426</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4480</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1688,213,-1688</points>
<connection>
<GID>6426</GID>
<name>clock</name></connection>
<connection>
<GID>6422</GID>
<name>clock</name></connection>
<connection>
<GID>6418</GID>
<name>clock</name></connection>
<connection>
<GID>6412</GID>
<name>clock</name></connection>
<connection>
<GID>6406</GID>
<name>clock</name></connection>
<connection>
<GID>6398</GID>
<name>clock</name></connection>
<connection>
<GID>6392</GID>
<name>clock</name></connection>
<connection>
<GID>6356</GID>
<name>clock</name></connection>
<connection>
<GID>6350</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4481</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1697.5,224,-1697.5</points>
<connection>
<GID>6428</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6424</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6420</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6416</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6410</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6402</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6394</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6368</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6352</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4482</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1682,61,-1682</points>
<connection>
<GID>6436</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1682,55,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1666.5,55,-1666.5</points>
<connection>
<GID>6434</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1682,84,-1682</points>
<connection>
<GID>6440</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1682,78,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1666.5,78,-1666.5</points>
<connection>
<GID>6438</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4484</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1682,109,-1682</points>
<connection>
<GID>6444</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1682,103,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1666.5,103,-1666.5</points>
<connection>
<GID>6442</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1682,132,-1682</points>
<connection>
<GID>6448</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1682,126,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1666.5,126,-1666.5</points>
<connection>
<GID>6446</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1682,155,-1682</points>
<connection>
<GID>6452</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1682,149,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1666.5,149,-1666.5</points>
<connection>
<GID>6450</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1682,178,-1682</points>
<connection>
<GID>6456</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1682,172,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1666.5,172,-1666.5</points>
<connection>
<GID>6454</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4488</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1682,203,-1682</points>
<connection>
<GID>6460</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1682,197,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1666.5,197,-1666.5</points>
<connection>
<GID>6458</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4489</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1682,226,-1682</points>
<connection>
<GID>6464</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1682,220,-1666.5</points>
<intersection>-1682 1</intersection>
<intersection>-1666.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1666.5,220,-1666.5</points>
<connection>
<GID>6462</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4490</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1669.5,213,-1669.5</points>
<connection>
<GID>6462</GID>
<name>clock</name></connection>
<connection>
<GID>6458</GID>
<name>clock</name></connection>
<connection>
<GID>6454</GID>
<name>clock</name></connection>
<connection>
<GID>6450</GID>
<name>clock</name></connection>
<connection>
<GID>6446</GID>
<name>clock</name></connection>
<connection>
<GID>6442</GID>
<name>clock</name></connection>
<connection>
<GID>6438</GID>
<name>clock</name></connection>
<connection>
<GID>6434</GID>
<name>clock</name></connection>
<connection>
<GID>6430</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1679,224,-1679</points>
<connection>
<GID>6464</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6460</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6456</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6452</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6448</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6444</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6440</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6436</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6432</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1663,61,-1663</points>
<connection>
<GID>6472</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1663,55,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1647.5,55,-1647.5</points>
<connection>
<GID>6470</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1663,84,-1663</points>
<connection>
<GID>6476</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1663,78,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1647.5,78,-1647.5</points>
<connection>
<GID>6474</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1663,109,-1663</points>
<connection>
<GID>6480</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1663,103,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1647.5,103,-1647.5</points>
<connection>
<GID>6478</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1663,132,-1663</points>
<connection>
<GID>6484</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1663,126,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1647.5,126,-1647.5</points>
<connection>
<GID>6482</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1663,155,-1663</points>
<connection>
<GID>6125</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1663,149,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1647.5,149,-1647.5</points>
<connection>
<GID>6486</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4497</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1663,178,-1663</points>
<connection>
<GID>6129</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1663,172,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1647.5,172,-1647.5</points>
<connection>
<GID>6127</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1663,203,-1663</points>
<connection>
<GID>6133</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1663,197,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1647.5,197,-1647.5</points>
<connection>
<GID>6131</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1663,226,-1663</points>
<connection>
<GID>6137</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1663,220,-1647.5</points>
<intersection>-1663 1</intersection>
<intersection>-1647.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1647.5,220,-1647.5</points>
<connection>
<GID>6135</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1650.5,213,-1650.5</points>
<connection>
<GID>6135</GID>
<name>clock</name></connection>
<connection>
<GID>6131</GID>
<name>clock</name></connection>
<connection>
<GID>6127</GID>
<name>clock</name></connection>
<connection>
<GID>6486</GID>
<name>clock</name></connection>
<connection>
<GID>6482</GID>
<name>clock</name></connection>
<connection>
<GID>6478</GID>
<name>clock</name></connection>
<connection>
<GID>6474</GID>
<name>clock</name></connection>
<connection>
<GID>6470</GID>
<name>clock</name></connection>
<connection>
<GID>6466</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1660,224,-1660</points>
<connection>
<GID>6137</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6133</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6129</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6125</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6484</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6480</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6476</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6472</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6468</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4502</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1644.5,61,-1644.5</points>
<connection>
<GID>6145</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1644.5,55,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1629,55,-1629</points>
<connection>
<GID>6143</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4503</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1644.5,84,-1644.5</points>
<connection>
<GID>6149</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1644.5,78,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1629,78,-1629</points>
<connection>
<GID>6147</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4504</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1644.5,109,-1644.5</points>
<connection>
<GID>6153</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1644.5,103,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1629,103,-1629</points>
<connection>
<GID>6151</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1644.5,132,-1644.5</points>
<connection>
<GID>6157</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1644.5,126,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1629,126,-1629</points>
<connection>
<GID>6155</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1644.5,155,-1644.5</points>
<connection>
<GID>6161</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1644.5,149,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1629,149,-1629</points>
<connection>
<GID>6159</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1644.5,178,-1644.5</points>
<connection>
<GID>6165</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1644.5,172,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1629,172,-1629</points>
<connection>
<GID>6163</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1644.5,203,-1644.5</points>
<connection>
<GID>6169</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1644.5,197,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1629,197,-1629</points>
<connection>
<GID>6167</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1644.5,226,-1644.5</points>
<connection>
<GID>6173</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1644.5,220,-1629</points>
<intersection>-1644.5 1</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1629,220,-1629</points>
<connection>
<GID>6171</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1632,213,-1632</points>
<connection>
<GID>6155</GID>
<name>clock</name></connection>
<connection>
<GID>6151</GID>
<name>clock</name></connection>
<connection>
<GID>6147</GID>
<name>clock</name></connection>
<connection>
<GID>6143</GID>
<name>clock</name></connection>
<connection>
<GID>6139</GID>
<name>OUT</name></connection>
<connection>
<GID>6171</GID>
<name>clock</name></connection>
<connection>
<GID>6167</GID>
<name>clock</name></connection>
<connection>
<GID>6163</GID>
<name>clock</name></connection>
<connection>
<GID>6159</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-1641.5,224,-1641.5</points>
<connection>
<GID>6157</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6153</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6149</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6145</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6141</GID>
<name>OUT</name></connection>
<connection>
<GID>6173</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6169</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6165</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6161</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1778.5,61,-1778.5</points>
<connection>
<GID>6182</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1778.5,55,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1763,55,-1763</points>
<connection>
<GID>6179</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1778.5,84,-1778.5</points>
<connection>
<GID>6187</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1778.5,78,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1763,78,-1763</points>
<connection>
<GID>6184</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1778.5,109,-1778.5</points>
<connection>
<GID>6192</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1778.5,103,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1763,103,-1763</points>
<connection>
<GID>6189</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4515</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1778.5,132,-1778.5</points>
<connection>
<GID>6197</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1778.5,126,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1763,126,-1763</points>
<connection>
<GID>6194</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1778.5,155,-1778.5</points>
<connection>
<GID>6202</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1778.5,149,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1763,149,-1763</points>
<connection>
<GID>6199</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1778.5,178,-1778.5</points>
<connection>
<GID>6207</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1778.5,172,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1763,172,-1763</points>
<connection>
<GID>6204</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1778.5,203,-1778.5</points>
<connection>
<GID>6274</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1778.5,197,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1763,197,-1763</points>
<connection>
<GID>6273</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4519</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1778.5,226,-1778.5</points>
<connection>
<GID>6276</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1778.5,220,-1763</points>
<intersection>-1778.5 1</intersection>
<intersection>-1763 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1763,220,-1763</points>
<connection>
<GID>6275</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1766,213,-1766</points>
<connection>
<GID>6275</GID>
<name>clock</name></connection>
<connection>
<GID>6273</GID>
<name>clock</name></connection>
<connection>
<GID>6204</GID>
<name>clock</name></connection>
<connection>
<GID>6199</GID>
<name>clock</name></connection>
<connection>
<GID>6194</GID>
<name>clock</name></connection>
<connection>
<GID>6189</GID>
<name>clock</name></connection>
<connection>
<GID>6184</GID>
<name>clock</name></connection>
<connection>
<GID>6179</GID>
<name>clock</name></connection>
<connection>
<GID>6175</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1775.5,224,-1775.5</points>
<connection>
<GID>6276</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6274</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6207</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6202</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6197</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6192</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6187</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6182</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6177</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1760,61,-1760</points>
<connection>
<GID>6280</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1760,55,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1744.5,55,-1744.5</points>
<connection>
<GID>6279</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1760,84,-1760</points>
<connection>
<GID>6282</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1760,78,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1744.5,78,-1744.5</points>
<connection>
<GID>6281</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1760,109,-1760</points>
<connection>
<GID>6284</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1760,103,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1744.5,103,-1744.5</points>
<connection>
<GID>6283</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1760,132,-1760</points>
<connection>
<GID>6286</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1760,126,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1744.5,126,-1744.5</points>
<connection>
<GID>6285</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1760,155,-1760</points>
<connection>
<GID>6288</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1760,149,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1744.5,149,-1744.5</points>
<connection>
<GID>6287</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1760,178,-1760</points>
<connection>
<GID>6290</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1760,172,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1744.5,172,-1744.5</points>
<connection>
<GID>6289</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1760,203,-1760</points>
<connection>
<GID>6292</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1760,197,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1744.5,197,-1744.5</points>
<connection>
<GID>6291</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1760,226,-1760</points>
<connection>
<GID>6294</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1760,220,-1744.5</points>
<intersection>-1760 1</intersection>
<intersection>-1744.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1744.5,220,-1744.5</points>
<connection>
<GID>6293</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1747.5,213,-1747.5</points>
<connection>
<GID>6293</GID>
<name>clock</name></connection>
<connection>
<GID>6291</GID>
<name>clock</name></connection>
<connection>
<GID>6289</GID>
<name>clock</name></connection>
<connection>
<GID>6287</GID>
<name>clock</name></connection>
<connection>
<GID>6285</GID>
<name>clock</name></connection>
<connection>
<GID>6283</GID>
<name>clock</name></connection>
<connection>
<GID>6281</GID>
<name>clock</name></connection>
<connection>
<GID>6279</GID>
<name>clock</name></connection>
<connection>
<GID>6277</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1757,224,-1757</points>
<connection>
<GID>6294</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6292</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6290</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6288</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6286</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6284</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6282</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6280</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6278</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1741,61,-1741</points>
<connection>
<GID>6190</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1741,55,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1725.5,55,-1725.5</points>
<connection>
<GID>6185</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1741,84,-1741</points>
<connection>
<GID>6200</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1741,78,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1725.5,78,-1725.5</points>
<connection>
<GID>6195</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1741,109,-1741</points>
<connection>
<GID>6209</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1741,103,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1725.5,103,-1725.5</points>
<connection>
<GID>6205</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1741,132,-1741</points>
<connection>
<GID>6296</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1741,126,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1725.5,126,-1725.5</points>
<connection>
<GID>6212</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1741,155,-1741</points>
<connection>
<GID>6298</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1741,149,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1725.5,149,-1725.5</points>
<connection>
<GID>6297</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1741,178,-1741</points>
<connection>
<GID>6300</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1741,172,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1725.5,172,-1725.5</points>
<connection>
<GID>6299</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4538</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1741,203,-1741</points>
<connection>
<GID>6302</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1741,197,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1725.5,197,-1725.5</points>
<connection>
<GID>6301</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1741,226,-1741</points>
<connection>
<GID>6305</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1741,220,-1725.5</points>
<intersection>-1741 1</intersection>
<intersection>-1725.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1725.5,220,-1725.5</points>
<connection>
<GID>6304</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4540</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1728.5,213,-1728.5</points>
<connection>
<GID>6304</GID>
<name>clock</name></connection>
<connection>
<GID>6301</GID>
<name>clock</name></connection>
<connection>
<GID>6299</GID>
<name>clock</name></connection>
<connection>
<GID>6297</GID>
<name>clock</name></connection>
<connection>
<GID>6295</GID>
<name>OUT</name></connection>
<connection>
<GID>6212</GID>
<name>clock</name></connection>
<connection>
<GID>6205</GID>
<name>clock</name></connection>
<connection>
<GID>6195</GID>
<name>clock</name></connection>
<connection>
<GID>6185</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4541</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1738,224,-1738</points>
<connection>
<GID>6305</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6302</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6300</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6298</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6296</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6209</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6200</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6190</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6180</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4542</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-1722.5,61,-1722.5</points>
<connection>
<GID>6310</GID>
<name>IN_0</name></connection>
<intersection>55 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55,-1722.5,55,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>54,-1707,55,-1707</points>
<connection>
<GID>6309</GID>
<name>OUT_0</name></connection>
<intersection>55 2</intersection></hsegment></shape></wire>
<wire>
<ID>4543</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-1722.5,84,-1722.5</points>
<connection>
<GID>6312</GID>
<name>IN_0</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-1722.5,78,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-1707,78,-1707</points>
<connection>
<GID>6311</GID>
<name>OUT_0</name></connection>
<intersection>78 2</intersection></hsegment></shape></wire>
<wire>
<ID>4544</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-1722.5,109,-1722.5</points>
<connection>
<GID>6315</GID>
<name>IN_0</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-1722.5,103,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>102,-1707,103,-1707</points>
<connection>
<GID>6314</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>4545</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-1722.5,132,-1722.5</points>
<connection>
<GID>6317</GID>
<name>IN_0</name></connection>
<intersection>126 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-1722.5,126,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>125,-1707,126,-1707</points>
<connection>
<GID>6316</GID>
<name>OUT_0</name></connection>
<intersection>126 2</intersection></hsegment></shape></wire>
<wire>
<ID>4546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149,-1722.5,155,-1722.5</points>
<connection>
<GID>6320</GID>
<name>IN_0</name></connection>
<intersection>149 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>149,-1722.5,149,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>148,-1707,149,-1707</points>
<connection>
<GID>6318</GID>
<name>OUT_0</name></connection>
<intersection>149 2</intersection></hsegment></shape></wire>
<wire>
<ID>4547</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-1722.5,178,-1722.5</points>
<connection>
<GID>6322</GID>
<name>IN_0</name></connection>
<intersection>172 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172,-1722.5,172,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171,-1707,172,-1707</points>
<connection>
<GID>6321</GID>
<name>OUT_0</name></connection>
<intersection>172 2</intersection></hsegment></shape></wire>
<wire>
<ID>4548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-1722.5,203,-1722.5</points>
<connection>
<GID>6324</GID>
<name>IN_0</name></connection>
<intersection>197 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>197,-1722.5,197,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>196,-1707,197,-1707</points>
<connection>
<GID>6323</GID>
<name>OUT_0</name></connection>
<intersection>197 2</intersection></hsegment></shape></wire>
<wire>
<ID>4549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-1722.5,226,-1722.5</points>
<connection>
<GID>6326</GID>
<name>IN_0</name></connection>
<intersection>220 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>220,-1722.5,220,-1707</points>
<intersection>-1722.5 1</intersection>
<intersection>-1707 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>219,-1707,220,-1707</points>
<connection>
<GID>6325</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection></hsegment></shape></wire>
<wire>
<ID>4550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1710,213,-1710</points>
<connection>
<GID>6325</GID>
<name>clock</name></connection>
<connection>
<GID>6323</GID>
<name>clock</name></connection>
<connection>
<GID>6321</GID>
<name>clock</name></connection>
<connection>
<GID>6318</GID>
<name>clock</name></connection>
<connection>
<GID>6316</GID>
<name>clock</name></connection>
<connection>
<GID>6314</GID>
<name>clock</name></connection>
<connection>
<GID>6311</GID>
<name>clock</name></connection>
<connection>
<GID>6309</GID>
<name>clock</name></connection>
<connection>
<GID>6306</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4551</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1719.5,224,-1719.5</points>
<connection>
<GID>6326</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6324</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6322</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6320</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6317</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6315</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6312</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6310</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6307</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-1788.5,42.5,-1623.5</points>
<connection>
<GID>6354</GID>
<name>N_in1</name></connection>
<connection>
<GID>6327</GID>
<name>N_in0</name></connection>
<intersection>-1763 12</intersection>
<intersection>-1744.5 11</intersection>
<intersection>-1725.5 10</intersection>
<intersection>-1707 9</intersection>
<intersection>-1685 8</intersection>
<intersection>-1666.5 7</intersection>
<intersection>-1647.5 6</intersection>
<intersection>-1629 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-1629,48,-1629</points>
<connection>
<GID>6143</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>42.5,-1647.5,48,-1647.5</points>
<connection>
<GID>6470</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>42.5,-1666.5,48,-1666.5</points>
<connection>
<GID>6434</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>42.5,-1685,48,-1685</points>
<connection>
<GID>6356</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42.5,-1707,48,-1707</points>
<connection>
<GID>6309</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>42.5,-1725.5,48,-1725.5</points>
<connection>
<GID>6185</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>42.5,-1744.5,48,-1744.5</points>
<connection>
<GID>6279</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>42.5,-1763,48,-1763</points>
<connection>
<GID>6179</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-1788,65.5,-1623</points>
<connection>
<GID>6358</GID>
<name>N_in1</name></connection>
<connection>
<GID>6328</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 4</intersection>
<intersection>-1754 5</intersection>
<intersection>-1735 6</intersection>
<intersection>-1716.5 7</intersection>
<intersection>-1694.5 8</intersection>
<intersection>-1676 9</intersection>
<intersection>-1657 10</intersection>
<intersection>-1638.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>61,-1772.5,65.5,-1772.5</points>
<intersection>61 12</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61,-1754,65.5,-1754</points>
<intersection>61 14</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61,-1735,65.5,-1735</points>
<intersection>61 13</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61,-1716.5,65.5,-1716.5</points>
<intersection>61 15</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61,-1694.5,65.5,-1694.5</points>
<intersection>61 18</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61,-1676,65.5,-1676</points>
<intersection>61 19</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61,-1657,65.5,-1657</points>
<intersection>61 20</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>61,-1638.5,65.5,-1638.5</points>
<intersection>61 21</intersection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>61,-1773,61,-1772.5</points>
<connection>
<GID>6182</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>61,-1735.5,61,-1735</points>
<connection>
<GID>6190</GID>
<name>OUT_0</name></connection>
<intersection>-1735 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>61,-1754.5,61,-1754</points>
<connection>
<GID>6280</GID>
<name>OUT_0</name></connection>
<intersection>-1754 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>61,-1717,61,-1716.5</points>
<connection>
<GID>6310</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>61,-1695,61,-1694.5</points>
<connection>
<GID>6368</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>61,-1676.5,61,-1676</points>
<connection>
<GID>6436</GID>
<name>OUT_0</name></connection>
<intersection>-1676 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>61,-1657.5,61,-1657</points>
<connection>
<GID>6472</GID>
<name>OUT_0</name></connection>
<intersection>-1657 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>61,-1639,61,-1638.5</points>
<connection>
<GID>6145</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>4554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-1788,68.5,-1623.5</points>
<connection>
<GID>6360</GID>
<name>N_in1</name></connection>
<connection>
<GID>6329</GID>
<name>N_in0</name></connection>
<intersection>-1763 10</intersection>
<intersection>-1744.5 9</intersection>
<intersection>-1725.5 8</intersection>
<intersection>-1707 7</intersection>
<intersection>-1685 6</intersection>
<intersection>-1666.5 5</intersection>
<intersection>-1647.5 4</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>68.5,-1629,71,-1629</points>
<connection>
<GID>6147</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-1647.5,71,-1647.5</points>
<connection>
<GID>6474</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68.5,-1666.5,71,-1666.5</points>
<connection>
<GID>6438</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68.5,-1685,71,-1685</points>
<connection>
<GID>6392</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68.5,-1707,71,-1707</points>
<connection>
<GID>6311</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-1725.5,71,-1725.5</points>
<connection>
<GID>6195</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68.5,-1744.5,71,-1744.5</points>
<connection>
<GID>6281</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68.5,-1763,71,-1763</points>
<connection>
<GID>6184</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-1788,88,-1623</points>
<connection>
<GID>6362</GID>
<name>N_in1</name></connection>
<connection>
<GID>6330</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 6</intersection>
<intersection>-1754 7</intersection>
<intersection>-1735 8</intersection>
<intersection>-1716.5 9</intersection>
<intersection>-1694.5 10</intersection>
<intersection>-1676 11</intersection>
<intersection>-1657 12</intersection>
<intersection>-1638.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84,-1772.5,88,-1772.5</points>
<intersection>84 14</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84,-1754,88,-1754</points>
<intersection>84 16</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>84,-1735,88,-1735</points>
<intersection>84 15</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84,-1716.5,88,-1716.5</points>
<intersection>84 17</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84,-1694.5,88,-1694.5</points>
<intersection>84 20</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84,-1676,88,-1676</points>
<intersection>84 21</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>84,-1657,88,-1657</points>
<intersection>84 22</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>84,-1638.5,88,-1638.5</points>
<intersection>84 23</intersection>
<intersection>88 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>84,-1773,84,-1772.5</points>
<connection>
<GID>6187</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>84,-1735.5,84,-1735</points>
<connection>
<GID>6200</GID>
<name>OUT_0</name></connection>
<intersection>-1735 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>84,-1754.5,84,-1754</points>
<connection>
<GID>6282</GID>
<name>OUT_0</name></connection>
<intersection>-1754 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>84,-1717,84,-1716.5</points>
<connection>
<GID>6312</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>84,-1695,84,-1694.5</points>
<connection>
<GID>6394</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>84,-1676.5,84,-1676</points>
<connection>
<GID>6440</GID>
<name>OUT_0</name></connection>
<intersection>-1676 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>84,-1657.5,84,-1657</points>
<connection>
<GID>6476</GID>
<name>OUT_0</name></connection>
<intersection>-1657 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>84,-1639,84,-1638.5</points>
<connection>
<GID>6149</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-1788,91.5,-1623</points>
<connection>
<GID>6364</GID>
<name>N_in1</name></connection>
<connection>
<GID>6331</GID>
<name>N_in0</name></connection>
<intersection>-1763 13</intersection>
<intersection>-1744.5 12</intersection>
<intersection>-1725.5 11</intersection>
<intersection>-1707 10</intersection>
<intersection>-1685 9</intersection>
<intersection>-1666.5 8</intersection>
<intersection>-1647.5 7</intersection>
<intersection>-1629 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>91.5,-1629,96,-1629</points>
<connection>
<GID>6151</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>91.5,-1647.5,96,-1647.5</points>
<connection>
<GID>6478</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>91.5,-1666.5,96,-1666.5</points>
<connection>
<GID>6442</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>91.5,-1685,96,-1685</points>
<connection>
<GID>6398</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>91.5,-1707,96,-1707</points>
<connection>
<GID>6314</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>91.5,-1725.5,96,-1725.5</points>
<connection>
<GID>6205</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>91.5,-1744.5,96,-1744.5</points>
<connection>
<GID>6283</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>91.5,-1763,96,-1763</points>
<connection>
<GID>6189</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-1788,112.5,-1623.5</points>
<connection>
<GID>6366</GID>
<name>N_in1</name></connection>
<connection>
<GID>6332</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 6</intersection>
<intersection>-1754 7</intersection>
<intersection>-1735 8</intersection>
<intersection>-1716.5 9</intersection>
<intersection>-1694.5 10</intersection>
<intersection>-1676 11</intersection>
<intersection>-1657 12</intersection>
<intersection>-1638.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109,-1772.5,112.5,-1772.5</points>
<intersection>109 14</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>109,-1754,112.5,-1754</points>
<intersection>109 16</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109,-1735,112.5,-1735</points>
<intersection>109 15</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>109,-1716.5,112.5,-1716.5</points>
<intersection>109 17</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>109,-1694.5,112.5,-1694.5</points>
<intersection>109 20</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>109,-1676,112.5,-1676</points>
<intersection>109 21</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109,-1657,112.5,-1657</points>
<intersection>109 22</intersection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>109,-1638.5,112.5,-1638.5</points>
<intersection>109 23</intersection>
<intersection>112.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>109,-1773,109,-1772.5</points>
<connection>
<GID>6192</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>109,-1735.5,109,-1735</points>
<connection>
<GID>6209</GID>
<name>OUT_0</name></connection>
<intersection>-1735 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>109,-1754.5,109,-1754</points>
<connection>
<GID>6284</GID>
<name>OUT_0</name></connection>
<intersection>-1754 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>109,-1717,109,-1716.5</points>
<connection>
<GID>6315</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>109,-1695,109,-1694.5</points>
<connection>
<GID>6402</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>109,-1676.5,109,-1676</points>
<connection>
<GID>6444</GID>
<name>OUT_0</name></connection>
<intersection>-1676 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>109,-1657.5,109,-1657</points>
<connection>
<GID>6480</GID>
<name>OUT_0</name></connection>
<intersection>-1657 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>109,-1639,109,-1638.5</points>
<connection>
<GID>6153</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-1788,116.5,-1623</points>
<connection>
<GID>6370</GID>
<name>N_in1</name></connection>
<connection>
<GID>6333</GID>
<name>N_in0</name></connection>
<intersection>-1763 13</intersection>
<intersection>-1744.5 12</intersection>
<intersection>-1725.5 11</intersection>
<intersection>-1707 10</intersection>
<intersection>-1685 9</intersection>
<intersection>-1666.5 8</intersection>
<intersection>-1647.5 7</intersection>
<intersection>-1629 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116.5,-1629,119,-1629</points>
<connection>
<GID>6155</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116.5,-1647.5,119,-1647.5</points>
<connection>
<GID>6482</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>116.5,-1666.5,119,-1666.5</points>
<connection>
<GID>6446</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116.5,-1685,119,-1685</points>
<connection>
<GID>6406</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116.5,-1707,119,-1707</points>
<connection>
<GID>6316</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>116.5,-1725.5,119,-1725.5</points>
<connection>
<GID>6212</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>116.5,-1744.5,119,-1744.5</points>
<connection>
<GID>6285</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>116.5,-1763,119,-1763</points>
<connection>
<GID>6194</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-1788,135,-1623</points>
<connection>
<GID>6372</GID>
<name>N_in1</name></connection>
<connection>
<GID>6334</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 6</intersection>
<intersection>-1754 7</intersection>
<intersection>-1735 8</intersection>
<intersection>-1716.5 9</intersection>
<intersection>-1694.5 10</intersection>
<intersection>-1676 11</intersection>
<intersection>-1657 12</intersection>
<intersection>-1638.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>132,-1772.5,135,-1772.5</points>
<intersection>132 14</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>132,-1754,135,-1754</points>
<intersection>132 15</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>132,-1735,135,-1735</points>
<intersection>132 16</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>132,-1716.5,135,-1716.5</points>
<intersection>132 17</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132,-1694.5,135,-1694.5</points>
<intersection>132 20</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132,-1676,135,-1676</points>
<intersection>132 21</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>132,-1657,135,-1657</points>
<intersection>132 22</intersection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132,-1638.5,135,-1638.5</points>
<intersection>132 23</intersection>
<intersection>135 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>132,-1773,132,-1772.5</points>
<connection>
<GID>6197</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>132,-1754.5,132,-1754</points>
<connection>
<GID>6286</GID>
<name>OUT_0</name></connection>
<intersection>-1754 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>132,-1735.5,132,-1735</points>
<connection>
<GID>6296</GID>
<name>OUT_0</name></connection>
<intersection>-1735 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>132,-1717,132,-1716.5</points>
<connection>
<GID>6317</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>132,-1695,132,-1694.5</points>
<connection>
<GID>6410</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>132,-1676.5,132,-1676</points>
<connection>
<GID>6448</GID>
<name>OUT_0</name></connection>
<intersection>-1676 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>132,-1657.5,132,-1657</points>
<connection>
<GID>6484</GID>
<name>OUT_0</name></connection>
<intersection>-1657 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>132,-1639,132,-1638.5</points>
<connection>
<GID>6157</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-1788,139,-1623</points>
<connection>
<GID>6374</GID>
<name>N_in1</name></connection>
<connection>
<GID>6336</GID>
<name>N_in0</name></connection>
<intersection>-1763 13</intersection>
<intersection>-1744.5 12</intersection>
<intersection>-1725.5 11</intersection>
<intersection>-1707 10</intersection>
<intersection>-1685 9</intersection>
<intersection>-1666.5 8</intersection>
<intersection>-1647.5 7</intersection>
<intersection>-1629 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-1629,142,-1629</points>
<connection>
<GID>6159</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,-1647.5,142,-1647.5</points>
<connection>
<GID>6486</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>139,-1666.5,142,-1666.5</points>
<connection>
<GID>6450</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>139,-1685,142,-1685</points>
<connection>
<GID>6412</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>139,-1707,142,-1707</points>
<connection>
<GID>6318</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139,-1725.5,142,-1725.5</points>
<connection>
<GID>6297</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>139,-1744.5,142,-1744.5</points>
<connection>
<GID>6287</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>139,-1763,142,-1763</points>
<connection>
<GID>6199</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>4561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-1787.5,158,-1623</points>
<connection>
<GID>6376</GID>
<name>N_in1</name></connection>
<connection>
<GID>6338</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 6</intersection>
<intersection>-1754 7</intersection>
<intersection>-1735 8</intersection>
<intersection>-1716.5 9</intersection>
<intersection>-1694.5 10</intersection>
<intersection>-1676 11</intersection>
<intersection>-1657 12</intersection>
<intersection>-1638.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>155,-1772.5,158,-1772.5</points>
<intersection>155 15</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>155,-1754,158,-1754</points>
<intersection>155 16</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>155,-1735,158,-1735</points>
<intersection>155 17</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>155,-1716.5,158,-1716.5</points>
<intersection>155 18</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>155,-1694.5,158,-1694.5</points>
<intersection>155 21</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>155,-1676,158,-1676</points>
<intersection>155 22</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>155,-1657,158,-1657</points>
<intersection>155 23</intersection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>155,-1638.5,158,-1638.5</points>
<intersection>155 14</intersection>
<intersection>158 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>155,-1639,155,-1638.5</points>
<connection>
<GID>6161</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>155,-1773,155,-1772.5</points>
<connection>
<GID>6202</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>155,-1754.5,155,-1754</points>
<connection>
<GID>6288</GID>
<name>OUT_0</name></connection>
<intersection>-1754 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>155,-1735.5,155,-1735</points>
<connection>
<GID>6298</GID>
<name>OUT_0</name></connection>
<intersection>-1735 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>155,-1717,155,-1716.5</points>
<connection>
<GID>6320</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>155,-1695,155,-1694.5</points>
<connection>
<GID>6416</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>155,-1676.5,155,-1676</points>
<connection>
<GID>6452</GID>
<name>OUT_0</name></connection>
<intersection>-1676 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>155,-1657.5,155,-1657</points>
<connection>
<GID>6125</GID>
<name>OUT_0</name></connection>
<intersection>-1657 12</intersection></vsegment></shape></wire>
<wire>
<ID>4562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-1787.5,163,-1623</points>
<connection>
<GID>6378</GID>
<name>N_in1</name></connection>
<connection>
<GID>6340</GID>
<name>N_in0</name></connection>
<intersection>-1763 13</intersection>
<intersection>-1744.5 12</intersection>
<intersection>-1725.5 11</intersection>
<intersection>-1707 10</intersection>
<intersection>-1685 9</intersection>
<intersection>-1666.5 8</intersection>
<intersection>-1647.5 7</intersection>
<intersection>-1629 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>163,-1629,165,-1629</points>
<connection>
<GID>6163</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>163,-1647.5,165,-1647.5</points>
<connection>
<GID>6127</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>163,-1666.5,165,-1666.5</points>
<connection>
<GID>6454</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>163,-1685,165,-1685</points>
<connection>
<GID>6418</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>163,-1707,165,-1707</points>
<connection>
<GID>6321</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>163,-1725.5,165,-1725.5</points>
<connection>
<GID>6299</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>163,-1744.5,165,-1744.5</points>
<connection>
<GID>6289</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>163,-1763,165,-1763</points>
<connection>
<GID>6204</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>4563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-1787,181,-1623</points>
<connection>
<GID>6380</GID>
<name>N_in1</name></connection>
<connection>
<GID>6344</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 16</intersection>
<intersection>-1754 15</intersection>
<intersection>-1735 14</intersection>
<intersection>-1716.5 13</intersection>
<intersection>-1694.5 12</intersection>
<intersection>-1676 11</intersection>
<intersection>-1657 10</intersection>
<intersection>-1638.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>178,-1638.5,181,-1638.5</points>
<intersection>178 17</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>178,-1657,181,-1657</points>
<intersection>178 26</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>178,-1676,181,-1676</points>
<intersection>178 25</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>178,-1694.5,181,-1694.5</points>
<intersection>178 24</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>178,-1716.5,181,-1716.5</points>
<intersection>178 21</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>178,-1735,181,-1735</points>
<intersection>178 20</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>178,-1754,181,-1754</points>
<intersection>178 19</intersection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>178,-1772.5,181,-1772.5</points>
<intersection>178 18</intersection>
<intersection>181 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>178,-1639,178,-1638.5</points>
<connection>
<GID>6165</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>178,-1773,178,-1772.5</points>
<connection>
<GID>6207</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>178,-1754.5,178,-1754</points>
<connection>
<GID>6290</GID>
<name>OUT_0</name></connection>
<intersection>-1754 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>178,-1735.5,178,-1735</points>
<connection>
<GID>6300</GID>
<name>OUT_0</name></connection>
<intersection>-1735 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>178,-1717,178,-1716.5</points>
<connection>
<GID>6322</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>178,-1695,178,-1694.5</points>
<connection>
<GID>6420</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>178,-1676.5,178,-1676</points>
<connection>
<GID>6456</GID>
<name>OUT_0</name></connection>
<intersection>-1676 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>178,-1657.5,178,-1657</points>
<connection>
<GID>6129</GID>
<name>OUT_0</name></connection>
<intersection>-1657 10</intersection></vsegment></shape></wire>
<wire>
<ID>4564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-1787,185.5,-1623</points>
<connection>
<GID>6382</GID>
<name>N_in1</name></connection>
<connection>
<GID>6342</GID>
<name>N_in0</name></connection>
<intersection>-1763 13</intersection>
<intersection>-1744.5 12</intersection>
<intersection>-1725.5 11</intersection>
<intersection>-1707 10</intersection>
<intersection>-1685 9</intersection>
<intersection>-1666.5 8</intersection>
<intersection>-1647.5 7</intersection>
<intersection>-1629 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>185.5,-1629,190,-1629</points>
<connection>
<GID>6167</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>185.5,-1647.5,190,-1647.5</points>
<connection>
<GID>6131</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>185.5,-1666.5,190,-1666.5</points>
<connection>
<GID>6458</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185.5,-1685,190,-1685</points>
<connection>
<GID>6422</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>185.5,-1707,190,-1707</points>
<connection>
<GID>6323</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>185.5,-1725.5,190,-1725.5</points>
<connection>
<GID>6301</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>185.5,-1744.5,190,-1744.5</points>
<connection>
<GID>6291</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>185.5,-1763,190,-1763</points>
<connection>
<GID>6273</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-1786.5,206.5,-1623.5</points>
<connection>
<GID>6384</GID>
<name>N_in1</name></connection>
<connection>
<GID>6346</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 6</intersection>
<intersection>-1754 7</intersection>
<intersection>-1735 8</intersection>
<intersection>-1716.5 9</intersection>
<intersection>-1694.5 10</intersection>
<intersection>-1676 11</intersection>
<intersection>-1657 12</intersection>
<intersection>-1638.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>203,-1772.5,206.5,-1772.5</points>
<intersection>203 15</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-1754,206.5,-1754</points>
<intersection>203 16</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>203,-1735,206.5,-1735</points>
<intersection>203 17</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>203,-1716.5,206.5,-1716.5</points>
<intersection>203 18</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>203,-1694.5,206.5,-1694.5</points>
<intersection>203 21</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-1676,206.5,-1676</points>
<intersection>203 22</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>203,-1657,206.5,-1657</points>
<intersection>203 23</intersection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>203,-1638.5,206.5,-1638.5</points>
<intersection>203 14</intersection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>203,-1639,203,-1638.5</points>
<connection>
<GID>6169</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>203,-1773,203,-1772.5</points>
<connection>
<GID>6274</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>203,-1754.5,203,-1754</points>
<connection>
<GID>6292</GID>
<name>OUT_0</name></connection>
<intersection>-1754 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>203,-1735.5,203,-1735</points>
<connection>
<GID>6302</GID>
<name>OUT_0</name></connection>
<intersection>-1735 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>203,-1717,203,-1716.5</points>
<connection>
<GID>6324</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>203,-1695,203,-1694.5</points>
<connection>
<GID>6424</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>203,-1676.5,203,-1676</points>
<connection>
<GID>6460</GID>
<name>OUT_0</name></connection>
<intersection>-1676 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>203,-1657.5,203,-1657</points>
<connection>
<GID>6133</GID>
<name>OUT_0</name></connection>
<intersection>-1657 12</intersection></vsegment></shape></wire>
<wire>
<ID>4566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-1786.5,210,-1623.5</points>
<connection>
<GID>6386</GID>
<name>N_in1</name></connection>
<connection>
<GID>6388</GID>
<name>N_in0</name></connection>
<intersection>-1763 11</intersection>
<intersection>-1744.5 10</intersection>
<intersection>-1725.5 9</intersection>
<intersection>-1707 7</intersection>
<intersection>-1685 6</intersection>
<intersection>-1666.5 5</intersection>
<intersection>-1647.5 4</intersection>
<intersection>-1629 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>210,-1629,213,-1629</points>
<connection>
<GID>6171</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>210,-1647.5,213,-1647.5</points>
<connection>
<GID>6135</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>210,-1666.5,213,-1666.5</points>
<connection>
<GID>6462</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>210,-1685,213,-1685</points>
<connection>
<GID>6426</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>210,-1707,213,-1707</points>
<connection>
<GID>6325</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>210,-1725.5,213,-1725.5</points>
<connection>
<GID>6304</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210,-1744.5,213,-1744.5</points>
<connection>
<GID>6293</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>210,-1763,213,-1763</points>
<connection>
<GID>6275</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>4567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,-1786.5,231,-1624.5</points>
<connection>
<GID>6390</GID>
<name>N_in1</name></connection>
<connection>
<GID>6348</GID>
<name>N_in0</name></connection>
<intersection>-1772.5 11</intersection>
<intersection>-1754 10</intersection>
<intersection>-1735 9</intersection>
<intersection>-1716.5 8</intersection>
<intersection>-1694.5 7</intersection>
<intersection>-1676 6</intersection>
<intersection>-1657 5</intersection>
<intersection>-1638.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>226,-1638.5,231,-1638.5</points>
<intersection>226 12</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>226,-1657,231,-1657</points>
<intersection>226 21</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>226,-1676,231,-1676</points>
<intersection>226 20</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>226,-1694.5,231,-1694.5</points>
<intersection>226 19</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>226,-1716.5,231,-1716.5</points>
<intersection>226 16</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>226,-1735,231,-1735</points>
<intersection>226 15</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>226,-1754,231,-1754</points>
<intersection>226 14</intersection>
<intersection>231 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>226,-1772.5,231,-1772.5</points>
<intersection>226 13</intersection>
<intersection>231 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>226,-1639,226,-1638.5</points>
<connection>
<GID>6173</GID>
<name>OUT_0</name></connection>
<intersection>-1638.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>226,-1773,226,-1772.5</points>
<connection>
<GID>6276</GID>
<name>OUT_0</name></connection>
<intersection>-1772.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>226,-1754.5,226,-1754</points>
<connection>
<GID>6294</GID>
<name>OUT_0</name></connection>
<intersection>-1754 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>226,-1735.5,226,-1735</points>
<connection>
<GID>6305</GID>
<name>OUT_0</name></connection>
<intersection>-1735 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>226,-1717,226,-1716.5</points>
<connection>
<GID>6326</GID>
<name>OUT_0</name></connection>
<intersection>-1716.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>226,-1695,226,-1694.5</points>
<connection>
<GID>6428</GID>
<name>OUT_0</name></connection>
<intersection>-1694.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>226,-1676.5,226,-1676</points>
<connection>
<GID>6464</GID>
<name>OUT_0</name></connection>
<intersection>-1676 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>226,-1657.5,226,-1657</points>
<connection>
<GID>6137</GID>
<name>OUT_0</name></connection>
<intersection>-1657 5</intersection></vsegment></shape></wire>
<wire>
<ID>4568</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-119,-1631,20.5,-1631</points>
<connection>
<GID>6139</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-1640.5,-119,-1615</points>
<intersection>-1640.5 4</intersection>
<intersection>-1631 2</intersection>
<intersection>-1615 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-1640.5,32,-1640.5</points>
<connection>
<GID>6141</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-126,-1615,-119,-1615</points>
<connection>
<GID>6272</GID>
<name>OUT_7</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>4569</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-120,-1649.5,20.5,-1649.5</points>
<connection>
<GID>6466</GID>
<name>IN_0</name></connection>
<intersection>-120 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-120,-1659,-120,-1616</points>
<intersection>-1659 5</intersection>
<intersection>-1649.5 2</intersection>
<intersection>-1616 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-120,-1659,32,-1659</points>
<connection>
<GID>6468</GID>
<name>IN_0</name></connection>
<intersection>-120 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-126,-1616,-120,-1616</points>
<connection>
<GID>6272</GID>
<name>OUT_6</name></connection>
<intersection>-120 4</intersection></hsegment></shape></wire>
<wire>
<ID>4570</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-121,-1668.5,20.5,-1668.5</points>
<connection>
<GID>6430</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-1678,-121,-1617</points>
<intersection>-1678 4</intersection>
<intersection>-1668.5 2</intersection>
<intersection>-1617 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-1678,32,-1678</points>
<connection>
<GID>6432</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-126,-1617,-121,-1617</points>
<connection>
<GID>6272</GID>
<name>OUT_5</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4571</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-122,-1687,20.5,-1687</points>
<connection>
<GID>6350</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-1696.5,-122,-1618</points>
<intersection>-1696.5 4</intersection>
<intersection>-1687 2</intersection>
<intersection>-1618 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-1696.5,32,-1696.5</points>
<connection>
<GID>6352</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1618,-122,-1618</points>
<connection>
<GID>6272</GID>
<name>OUT_4</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>4572</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123,-1709,20.5,-1709</points>
<connection>
<GID>6306</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-1718.5,-123,-1619</points>
<intersection>-1718.5 4</intersection>
<intersection>-1709 1</intersection>
<intersection>-1619 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-1718.5,31.5,-1718.5</points>
<connection>
<GID>6307</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1619,-123,-1619</points>
<connection>
<GID>6272</GID>
<name>OUT_3</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>4573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,-1727.5,20.5,-1727.5</points>
<connection>
<GID>6295</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-1737,-124,-1620</points>
<intersection>-1737 4</intersection>
<intersection>-1727.5 1</intersection>
<intersection>-1620 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-1737,31.5,-1737</points>
<connection>
<GID>6180</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1620,-124,-1620</points>
<connection>
<GID>6272</GID>
<name>OUT_2</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>4574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125,-1746.5,20.5,-1746.5</points>
<connection>
<GID>6277</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-125,-1756,-125,-1621</points>
<intersection>-1756 4</intersection>
<intersection>-1746.5 1</intersection>
<intersection>-1621 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-125,-1756,31.5,-1756</points>
<connection>
<GID>6278</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-126,-1621,-125,-1621</points>
<connection>
<GID>6272</GID>
<name>OUT_1</name></connection>
<intersection>-125 3</intersection></hsegment></shape></wire>
<wire>
<ID>4575</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,-1765,20.5,-1765</points>
<connection>
<GID>6175</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-1774.5,-126,-1622</points>
<connection>
<GID>6272</GID>
<name>OUT_0</name></connection>
<intersection>-1774.5 4</intersection>
<intersection>-1765 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-1774.5,31.5,-1774.5</points>
<connection>
<GID>6177</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>4576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-1788.5,19.5,-1623.5</points>
<connection>
<GID>6408</GID>
<name>N_in1</name></connection>
<connection>
<GID>6400</GID>
<name>N_in0</name></connection>
<intersection>-1767 10</intersection>
<intersection>-1748.5 9</intersection>
<intersection>-1729.5 8</intersection>
<intersection>-1711 7</intersection>
<intersection>-1689 6</intersection>
<intersection>-1670.5 5</intersection>
<intersection>-1651.5 4</intersection>
<intersection>-1633 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>19.5,-1633,20.5,-1633</points>
<connection>
<GID>6139</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>19.5,-1651.5,20.5,-1651.5</points>
<connection>
<GID>6466</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>19.5,-1670.5,20.5,-1670.5</points>
<connection>
<GID>6430</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>19.5,-1689,20.5,-1689</points>
<connection>
<GID>6350</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>19.5,-1711,20.5,-1711</points>
<connection>
<GID>6306</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>19.5,-1729.5,20.5,-1729.5</points>
<connection>
<GID>6295</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>19.5,-1748.5,20.5,-1748.5</points>
<connection>
<GID>6277</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>19.5,-1767,20.5,-1767</points>
<connection>
<GID>6175</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-1788.5,29.5,-1623.5</points>
<connection>
<GID>6404</GID>
<name>N_in1</name></connection>
<connection>
<GID>6396</GID>
<name>N_in0</name></connection>
<intersection>-1776.5 3</intersection>
<intersection>-1758 5</intersection>
<intersection>-1739 7</intersection>
<intersection>-1720.5 9</intersection>
<intersection>-1698.5 11</intersection>
<intersection>-1680 13</intersection>
<intersection>-1661 15</intersection>
<intersection>-1642.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-1776.5,31.5,-1776.5</points>
<connection>
<GID>6177</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>29.5,-1758,31.5,-1758</points>
<connection>
<GID>6278</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>29.5,-1739,31.5,-1739</points>
<connection>
<GID>6180</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>29.5,-1720.5,31.5,-1720.5</points>
<connection>
<GID>6307</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>29.5,-1698.5,32,-1698.5</points>
<connection>
<GID>6352</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>29.5,-1680,32,-1680</points>
<connection>
<GID>6432</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>29.5,-1661,32,-1661</points>
<connection>
<GID>6468</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>29.5,-1642.5,32,-1642.5</points>
<connection>
<GID>6141</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-1621.5,19.5,-1615</points>
<connection>
<GID>6400</GID>
<name>N_in1</name></connection>
<connection>
<GID>6270</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-1621.5,29.5,-1615</points>
<connection>
<GID>6396</GID>
<name>N_in1</name></connection>
<connection>
<GID>6269</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-1621.5,42.5,-1615</points>
<connection>
<GID>6327</GID>
<name>N_in1</name></connection>
<connection>
<GID>6250</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-1621,65.5,-1614.5</points>
<connection>
<GID>6328</GID>
<name>N_in1</name></connection>
<connection>
<GID>6251</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4582</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-1621.5,68.5,-1614.5</points>
<connection>
<GID>6329</GID>
<name>N_in1</name></connection>
<connection>
<GID>6252</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-1621,88,-1614.5</points>
<connection>
<GID>6330</GID>
<name>N_in1</name></connection>
<connection>
<GID>6253</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-1621,91.5,-1614.5</points>
<connection>
<GID>6331</GID>
<name>N_in1</name></connection>
<connection>
<GID>6254</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-1621.5,112.5,-1614.5</points>
<connection>
<GID>6332</GID>
<name>N_in1</name></connection>
<connection>
<GID>6255</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-1621,116.5,-1614.5</points>
<connection>
<GID>6333</GID>
<name>N_in1</name></connection>
<connection>
<GID>6256</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-1621,135,-1614.5</points>
<connection>
<GID>6334</GID>
<name>N_in1</name></connection>
<connection>
<GID>6257</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-1621,139,-1614.5</points>
<connection>
<GID>6336</GID>
<name>N_in1</name></connection>
<connection>
<GID>6258</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-1621,158,-1614</points>
<connection>
<GID>6338</GID>
<name>N_in1</name></connection>
<connection>
<GID>6259</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-1621,163,-1614</points>
<connection>
<GID>6340</GID>
<name>N_in1</name></connection>
<connection>
<GID>6260</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-1621,181,-1613.5</points>
<connection>
<GID>6344</GID>
<name>N_in1</name></connection>
<connection>
<GID>6261</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-1621,185.5,-1613.5</points>
<connection>
<GID>6342</GID>
<name>N_in1</name></connection>
<connection>
<GID>6262</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-1621.5,206.5,-1613</points>
<connection>
<GID>6346</GID>
<name>N_in1</name></connection>
<connection>
<GID>6263</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-1621.5,210,-1613</points>
<connection>
<GID>6388</GID>
<name>N_in1</name></connection>
<connection>
<GID>6264</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,-1622.5,231,-1613</points>
<connection>
<GID>6348</GID>
<name>N_in1</name></connection>
<connection>
<GID>6266</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4596</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1898,59,-1898</points>
<connection>
<GID>6684</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1898,53,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1882.5,53,-1882.5</points>
<connection>
<GID>6678</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1898,82,-1898</points>
<connection>
<GID>6702</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1898,76,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1882.5,76,-1882.5</points>
<connection>
<GID>6700</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4598</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1898,107,-1898</points>
<connection>
<GID>6706</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1898,101,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1882.5,101,-1882.5</points>
<connection>
<GID>6704</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1898,130,-1898</points>
<connection>
<GID>6710</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1898,124,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1882.5,124,-1882.5</points>
<connection>
<GID>6708</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4600</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1898,153,-1898</points>
<connection>
<GID>6714</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1898,147,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1882.5,147,-1882.5</points>
<connection>
<GID>6712</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4601</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1898,176,-1898</points>
<connection>
<GID>6718</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1898,170,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1882.5,170,-1882.5</points>
<connection>
<GID>6716</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4602</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1898,201,-1898</points>
<connection>
<GID>6722</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1898,195,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1882.5,195,-1882.5</points>
<connection>
<GID>6720</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4603</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1898,224,-1898</points>
<connection>
<GID>6726</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1898,218,-1882.5</points>
<intersection>-1898 1</intersection>
<intersection>-1882.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1882.5,218,-1882.5</points>
<connection>
<GID>6724</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4604</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1885.5,211,-1885.5</points>
<connection>
<GID>6668</GID>
<name>OUT</name></connection>
<connection>
<GID>6678</GID>
<name>clock</name></connection>
<connection>
<GID>6700</GID>
<name>clock</name></connection>
<connection>
<GID>6704</GID>
<name>clock</name></connection>
<connection>
<GID>6708</GID>
<name>clock</name></connection>
<connection>
<GID>6712</GID>
<name>clock</name></connection>
<connection>
<GID>6716</GID>
<name>clock</name></connection>
<connection>
<GID>6720</GID>
<name>clock</name></connection>
<connection>
<GID>6724</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4605</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-1895,222,-1895</points>
<connection>
<GID>6673</GID>
<name>OUT</name></connection>
<connection>
<GID>6684</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6702</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6706</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6710</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6714</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6718</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6722</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6726</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4606</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1879.5,59,-1879.5</points>
<connection>
<GID>6734</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1879.5,53,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1864,53,-1864</points>
<connection>
<GID>6732</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4607</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1879.5,82,-1879.5</points>
<connection>
<GID>6738</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1879.5,76,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1864,76,-1864</points>
<connection>
<GID>6736</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4608</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1879.5,107,-1879.5</points>
<connection>
<GID>6742</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1879.5,101,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1864,101,-1864</points>
<connection>
<GID>6740</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4609</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1879.5,130,-1879.5</points>
<connection>
<GID>6746</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1879.5,124,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1864,124,-1864</points>
<connection>
<GID>6744</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4610</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1879.5,153,-1879.5</points>
<connection>
<GID>6750</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1879.5,147,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1864,147,-1864</points>
<connection>
<GID>6748</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4611</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1879.5,176,-1879.5</points>
<connection>
<GID>6754</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1879.5,170,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1864,170,-1864</points>
<connection>
<GID>6752</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4612</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1879.5,201,-1879.5</points>
<connection>
<GID>6758</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1879.5,195,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1864,195,-1864</points>
<connection>
<GID>6756</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4613</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1879.5,224,-1879.5</points>
<connection>
<GID>6762</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1879.5,218,-1864</points>
<intersection>-1879.5 1</intersection>
<intersection>-1864 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1864,218,-1864</points>
<connection>
<GID>6760</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4614</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1867,211,-1867</points>
<connection>
<GID>6728</GID>
<name>OUT</name></connection>
<connection>
<GID>6732</GID>
<name>clock</name></connection>
<connection>
<GID>6736</GID>
<name>clock</name></connection>
<connection>
<GID>6740</GID>
<name>clock</name></connection>
<connection>
<GID>6744</GID>
<name>clock</name></connection>
<connection>
<GID>6748</GID>
<name>clock</name></connection>
<connection>
<GID>6752</GID>
<name>clock</name></connection>
<connection>
<GID>6756</GID>
<name>clock</name></connection>
<connection>
<GID>6760</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4615</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-1876.5,222,-1876.5</points>
<connection>
<GID>6730</GID>
<name>OUT</name></connection>
<connection>
<GID>6734</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6738</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6742</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6746</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6754</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6758</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6762</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4616</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1860.5,59,-1860.5</points>
<connection>
<GID>6770</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1860.5,53,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1845,53,-1845</points>
<connection>
<GID>6768</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4617</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1860.5,82,-1860.5</points>
<connection>
<GID>6774</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1860.5,76,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1845,76,-1845</points>
<connection>
<GID>6772</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1860.5,107,-1860.5</points>
<connection>
<GID>6778</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1860.5,101,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1845,101,-1845</points>
<connection>
<GID>6776</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4619</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1860.5,130,-1860.5</points>
<connection>
<GID>6782</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1860.5,124,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1845,124,-1845</points>
<connection>
<GID>6780</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4620</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1860.5,153,-1860.5</points>
<connection>
<GID>6786</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1860.5,147,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1845,147,-1845</points>
<connection>
<GID>6784</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4621</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1860.5,176,-1860.5</points>
<connection>
<GID>6790</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1860.5,170,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1845,170,-1845</points>
<connection>
<GID>6788</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1860.5,201,-1860.5</points>
<connection>
<GID>6794</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1860.5,195,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1845,195,-1845</points>
<connection>
<GID>6792</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4623</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1860.5,224,-1860.5</points>
<connection>
<GID>6798</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1860.5,218,-1845</points>
<intersection>-1860.5 1</intersection>
<intersection>-1845 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1845,218,-1845</points>
<connection>
<GID>6796</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4624</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1848,211,-1848</points>
<connection>
<GID>6764</GID>
<name>OUT</name></connection>
<connection>
<GID>6768</GID>
<name>clock</name></connection>
<connection>
<GID>6772</GID>
<name>clock</name></connection>
<connection>
<GID>6776</GID>
<name>clock</name></connection>
<connection>
<GID>6780</GID>
<name>clock</name></connection>
<connection>
<GID>6784</GID>
<name>clock</name></connection>
<connection>
<GID>6788</GID>
<name>clock</name></connection>
<connection>
<GID>6792</GID>
<name>clock</name></connection>
<connection>
<GID>6796</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-1857.5,222,-1857.5</points>
<connection>
<GID>6766</GID>
<name>OUT</name></connection>
<connection>
<GID>6770</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6774</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6778</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6782</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6786</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6790</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6794</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6798</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1842,59,-1842</points>
<connection>
<GID>6806</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1842,53,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1826.5,53,-1826.5</points>
<connection>
<GID>6804</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1842,82,-1842</points>
<connection>
<GID>6810</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1842,76,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1826.5,76,-1826.5</points>
<connection>
<GID>6808</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4628</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1842,107,-1842</points>
<connection>
<GID>6814</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1842,101,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1826.5,101,-1826.5</points>
<connection>
<GID>6812</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1842,130,-1842</points>
<connection>
<GID>6818</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1842,124,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1826.5,124,-1826.5</points>
<connection>
<GID>6816</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4630</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1842,153,-1842</points>
<connection>
<GID>6822</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1842,147,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1826.5,147,-1826.5</points>
<connection>
<GID>6820</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1842,176,-1842</points>
<connection>
<GID>6826</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1842,170,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1826.5,170,-1826.5</points>
<connection>
<GID>6824</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4632</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1842,201,-1842</points>
<connection>
<GID>6830</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1842,195,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1826.5,195,-1826.5</points>
<connection>
<GID>6828</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4633</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1842,224,-1842</points>
<connection>
<GID>6834</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1842,218,-1826.5</points>
<intersection>-1842 1</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1826.5,218,-1826.5</points>
<connection>
<GID>6832</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4634</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1829.5,211,-1829.5</points>
<connection>
<GID>6800</GID>
<name>OUT</name></connection>
<connection>
<GID>6804</GID>
<name>clock</name></connection>
<connection>
<GID>6808</GID>
<name>clock</name></connection>
<connection>
<GID>6812</GID>
<name>clock</name></connection>
<connection>
<GID>6816</GID>
<name>clock</name></connection>
<connection>
<GID>6820</GID>
<name>clock</name></connection>
<connection>
<GID>6824</GID>
<name>clock</name></connection>
<connection>
<GID>6828</GID>
<name>clock</name></connection>
<connection>
<GID>6832</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-1839,222,-1839</points>
<connection>
<GID>6802</GID>
<name>OUT</name></connection>
<connection>
<GID>6806</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6810</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6814</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6818</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6822</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6826</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6830</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6834</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4636</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1976,59,-1976</points>
<connection>
<GID>6842</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1976,53,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1960.5,53,-1960.5</points>
<connection>
<GID>6840</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1976,82,-1976</points>
<connection>
<GID>6846</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1976,76,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1960.5,76,-1960.5</points>
<connection>
<GID>6844</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1976,107,-1976</points>
<connection>
<GID>6850</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1976,101,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1960.5,101,-1960.5</points>
<connection>
<GID>6848</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1976,130,-1976</points>
<connection>
<GID>6491</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1976,124,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1960.5,124,-1960.5</points>
<connection>
<GID>6489</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4640</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1976,153,-1976</points>
<connection>
<GID>6495</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1976,147,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1960.5,147,-1960.5</points>
<connection>
<GID>6493</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4641</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1976,176,-1976</points>
<connection>
<GID>6499</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1976,170,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1960.5,170,-1960.5</points>
<connection>
<GID>6497</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4642</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1976,201,-1976</points>
<connection>
<GID>6503</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1976,195,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1960.5,195,-1960.5</points>
<connection>
<GID>6501</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4643</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1976,224,-1976</points>
<connection>
<GID>6507</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1976,218,-1960.5</points>
<intersection>-1976 1</intersection>
<intersection>-1960.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1960.5,218,-1960.5</points>
<connection>
<GID>6505</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4644</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1963.5,211,-1963.5</points>
<connection>
<GID>6848</GID>
<name>clock</name></connection>
<connection>
<GID>6844</GID>
<name>clock</name></connection>
<connection>
<GID>6840</GID>
<name>clock</name></connection>
<connection>
<GID>6836</GID>
<name>OUT</name></connection>
<connection>
<GID>6505</GID>
<name>clock</name></connection>
<connection>
<GID>6501</GID>
<name>clock</name></connection>
<connection>
<GID>6497</GID>
<name>clock</name></connection>
<connection>
<GID>6493</GID>
<name>clock</name></connection>
<connection>
<GID>6489</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-1973,222,-1973</points>
<connection>
<GID>6850</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6846</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6842</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6838</GID>
<name>OUT</name></connection>
<connection>
<GID>6507</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6503</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6499</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6495</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6491</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1957.5,59,-1957.5</points>
<connection>
<GID>6515</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1957.5,53,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1942,53,-1942</points>
<connection>
<GID>6513</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1957.5,82,-1957.5</points>
<connection>
<GID>6519</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1957.5,76,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1942,76,-1942</points>
<connection>
<GID>6517</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1957.5,107,-1957.5</points>
<connection>
<GID>6523</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1957.5,101,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1942,101,-1942</points>
<connection>
<GID>6521</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4649</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1957.5,130,-1957.5</points>
<connection>
<GID>6527</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1957.5,124,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1942,124,-1942</points>
<connection>
<GID>6525</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1957.5,153,-1957.5</points>
<connection>
<GID>6531</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1957.5,147,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1942,147,-1942</points>
<connection>
<GID>6529</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1957.5,176,-1957.5</points>
<connection>
<GID>6535</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1957.5,170,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1942,170,-1942</points>
<connection>
<GID>6533</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4652</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1957.5,201,-1957.5</points>
<connection>
<GID>6539</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1957.5,195,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1942,195,-1942</points>
<connection>
<GID>6537</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1957.5,224,-1957.5</points>
<connection>
<GID>6543</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1957.5,218,-1942</points>
<intersection>-1957.5 1</intersection>
<intersection>-1942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1942,218,-1942</points>
<connection>
<GID>6541</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4654</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1945,211,-1945</points>
<connection>
<GID>6509</GID>
<name>OUT</name></connection>
<connection>
<GID>6513</GID>
<name>clock</name></connection>
<connection>
<GID>6517</GID>
<name>clock</name></connection>
<connection>
<GID>6521</GID>
<name>clock</name></connection>
<connection>
<GID>6525</GID>
<name>clock</name></connection>
<connection>
<GID>6529</GID>
<name>clock</name></connection>
<connection>
<GID>6533</GID>
<name>clock</name></connection>
<connection>
<GID>6537</GID>
<name>clock</name></connection>
<connection>
<GID>6541</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4655</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-1954.5,222,-1954.5</points>
<connection>
<GID>6511</GID>
<name>OUT</name></connection>
<connection>
<GID>6515</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6519</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6523</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6527</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6531</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6535</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6539</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6543</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4656</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1938.5,59,-1938.5</points>
<connection>
<GID>6553</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1938.5,53,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1923,53,-1923</points>
<connection>
<GID>6551</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4657</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1938.5,82,-1938.5</points>
<connection>
<GID>6558</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1938.5,76,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1923,76,-1923</points>
<connection>
<GID>6556</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1938.5,107,-1938.5</points>
<connection>
<GID>6563</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1938.5,101,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1923,101,-1923</points>
<connection>
<GID>6561</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4659</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1938.5,130,-1938.5</points>
<connection>
<GID>6568</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1938.5,124,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1923,124,-1923</points>
<connection>
<GID>6566</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4660</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1938.5,153,-1938.5</points>
<connection>
<GID>6573</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1938.5,147,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1923,147,-1923</points>
<connection>
<GID>6571</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4661</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1938.5,176,-1938.5</points>
<connection>
<GID>6576</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1938.5,170,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1923,170,-1923</points>
<connection>
<GID>6575</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4662</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1938.5,201,-1938.5</points>
<connection>
<GID>6579</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1938.5,195,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1923,195,-1923</points>
<connection>
<GID>6578</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4663</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1938.5,224,-1938.5</points>
<connection>
<GID>6581</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1938.5,218,-1923</points>
<intersection>-1938.5 1</intersection>
<intersection>-1923 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1923,218,-1923</points>
<connection>
<GID>6580</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4664</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1926,211,-1926</points>
<connection>
<GID>6546</GID>
<name>OUT</name></connection>
<connection>
<GID>6551</GID>
<name>clock</name></connection>
<connection>
<GID>6556</GID>
<name>clock</name></connection>
<connection>
<GID>6561</GID>
<name>clock</name></connection>
<connection>
<GID>6566</GID>
<name>clock</name></connection>
<connection>
<GID>6571</GID>
<name>clock</name></connection>
<connection>
<GID>6575</GID>
<name>clock</name></connection>
<connection>
<GID>6578</GID>
<name>clock</name></connection>
<connection>
<GID>6580</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4665</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-1935.5,222,-1935.5</points>
<connection>
<GID>6548</GID>
<name>OUT</name></connection>
<connection>
<GID>6553</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6558</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6563</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6568</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6573</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6576</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6579</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6581</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4666</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-1920,59,-1920</points>
<connection>
<GID>6585</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-1920,53,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-1904.5,53,-1904.5</points>
<connection>
<GID>6584</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4667</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-1920,82,-1920</points>
<connection>
<GID>6587</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-1920,76,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-1904.5,76,-1904.5</points>
<connection>
<GID>6586</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-1920,107,-1920</points>
<connection>
<GID>6589</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-1920,101,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-1904.5,101,-1904.5</points>
<connection>
<GID>6588</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-1920,130,-1920</points>
<connection>
<GID>6591</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-1920,124,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-1904.5,124,-1904.5</points>
<connection>
<GID>6590</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4670</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-1920,153,-1920</points>
<connection>
<GID>6593</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-1920,147,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-1904.5,147,-1904.5</points>
<connection>
<GID>6592</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4671</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-1920,176,-1920</points>
<connection>
<GID>6595</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-1920,170,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-1904.5,170,-1904.5</points>
<connection>
<GID>6594</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4672</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-1920,201,-1920</points>
<connection>
<GID>6597</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-1920,195,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-1904.5,195,-1904.5</points>
<connection>
<GID>6596</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4673</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-1920,224,-1920</points>
<connection>
<GID>6599</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-1920,218,-1904.5</points>
<intersection>-1920 1</intersection>
<intersection>-1904.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-1904.5,218,-1904.5</points>
<connection>
<GID>6598</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4674</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-1907.5,211,-1907.5</points>
<connection>
<GID>6582</GID>
<name>OUT</name></connection>
<connection>
<GID>6584</GID>
<name>clock</name></connection>
<connection>
<GID>6586</GID>
<name>clock</name></connection>
<connection>
<GID>6588</GID>
<name>clock</name></connection>
<connection>
<GID>6590</GID>
<name>clock</name></connection>
<connection>
<GID>6592</GID>
<name>clock</name></connection>
<connection>
<GID>6594</GID>
<name>clock</name></connection>
<connection>
<GID>6596</GID>
<name>clock</name></connection>
<connection>
<GID>6598</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4675</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-1917,222,-1917</points>
<connection>
<GID>6583</GID>
<name>OUT</name></connection>
<connection>
<GID>6585</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6587</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6589</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6591</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6593</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6595</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6597</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6599</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-1986,40.5,-1821</points>
<connection>
<GID>6615</GID>
<name>N_in1</name></connection>
<connection>
<GID>6600</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 12</intersection>
<intersection>-1942 11</intersection>
<intersection>-1923 10</intersection>
<intersection>-1904.5 9</intersection>
<intersection>-1882.5 8</intersection>
<intersection>-1864 7</intersection>
<intersection>-1845 6</intersection>
<intersection>-1826.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-1826.5,46,-1826.5</points>
<connection>
<GID>6804</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40.5,-1845,46,-1845</points>
<connection>
<GID>6768</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>40.5,-1864,46,-1864</points>
<connection>
<GID>6732</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>40.5,-1882.5,46,-1882.5</points>
<connection>
<GID>6678</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>40.5,-1904.5,46,-1904.5</points>
<connection>
<GID>6584</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>40.5,-1923,46,-1923</points>
<connection>
<GID>6551</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>40.5,-1942,46,-1942</points>
<connection>
<GID>6513</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>40.5,-1960.5,46,-1960.5</points>
<connection>
<GID>6840</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-1985.5,63.5,-1820.5</points>
<connection>
<GID>6616</GID>
<name>N_in1</name></connection>
<connection>
<GID>6601</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 4</intersection>
<intersection>-1951 5</intersection>
<intersection>-1932 6</intersection>
<intersection>-1913.5 7</intersection>
<intersection>-1891.5 8</intersection>
<intersection>-1873 9</intersection>
<intersection>-1854 10</intersection>
<intersection>-1835.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>59,-1969.5,63.5,-1969.5</points>
<intersection>59 12</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>59,-1951,63.5,-1951</points>
<intersection>59 13</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59,-1932,63.5,-1932</points>
<intersection>59 14</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59,-1913.5,63.5,-1913.5</points>
<intersection>59 15</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>59,-1891.5,63.5,-1891.5</points>
<intersection>59 18</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>59,-1873,63.5,-1873</points>
<intersection>59 19</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>59,-1854,63.5,-1854</points>
<intersection>59 20</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>59,-1835.5,63.5,-1835.5</points>
<intersection>59 21</intersection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>59,-1970.5,59,-1969.5</points>
<connection>
<GID>6842</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>59,-1952,59,-1951</points>
<connection>
<GID>6515</GID>
<name>OUT_0</name></connection>
<intersection>-1951 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>59,-1933,59,-1932</points>
<connection>
<GID>6553</GID>
<name>OUT_0</name></connection>
<intersection>-1932 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>59,-1914.5,59,-1913.5</points>
<connection>
<GID>6585</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>59,-1892.5,59,-1891.5</points>
<connection>
<GID>6684</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>59,-1874,59,-1873</points>
<connection>
<GID>6734</GID>
<name>OUT_0</name></connection>
<intersection>-1873 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>59,-1855,59,-1854</points>
<connection>
<GID>6770</GID>
<name>OUT_0</name></connection>
<intersection>-1854 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>59,-1836.5,59,-1835.5</points>
<connection>
<GID>6806</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>4678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-1985.5,66.5,-1821</points>
<connection>
<GID>6617</GID>
<name>N_in1</name></connection>
<connection>
<GID>6602</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 10</intersection>
<intersection>-1942 9</intersection>
<intersection>-1923 8</intersection>
<intersection>-1904.5 7</intersection>
<intersection>-1882.5 6</intersection>
<intersection>-1864 5</intersection>
<intersection>-1845 4</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>66.5,-1826.5,69,-1826.5</points>
<connection>
<GID>6808</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-1845,69,-1845</points>
<connection>
<GID>6772</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66.5,-1864,69,-1864</points>
<connection>
<GID>6736</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66.5,-1882.5,69,-1882.5</points>
<connection>
<GID>6700</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66.5,-1904.5,69,-1904.5</points>
<connection>
<GID>6586</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-1923,69,-1923</points>
<connection>
<GID>6556</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66.5,-1942,69,-1942</points>
<connection>
<GID>6517</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>66.5,-1960.5,69,-1960.5</points>
<connection>
<GID>6844</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-1985.5,86,-1820.5</points>
<connection>
<GID>6618</GID>
<name>N_in1</name></connection>
<connection>
<GID>6603</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 6</intersection>
<intersection>-1951 7</intersection>
<intersection>-1932 8</intersection>
<intersection>-1913.5 9</intersection>
<intersection>-1891.5 10</intersection>
<intersection>-1873 11</intersection>
<intersection>-1854 12</intersection>
<intersection>-1835.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>82,-1969.5,86,-1969.5</points>
<intersection>82 14</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82,-1951,86,-1951</points>
<intersection>82 15</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>82,-1932,86,-1932</points>
<intersection>82 16</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82,-1913.5,86,-1913.5</points>
<intersection>82 17</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>82,-1891.5,86,-1891.5</points>
<intersection>82 20</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>82,-1873,86,-1873</points>
<intersection>82 21</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>82,-1854,86,-1854</points>
<intersection>82 22</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>82,-1835.5,86,-1835.5</points>
<intersection>82 23</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>82,-1970.5,82,-1969.5</points>
<connection>
<GID>6846</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>82,-1952,82,-1951</points>
<connection>
<GID>6519</GID>
<name>OUT_0</name></connection>
<intersection>-1951 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>82,-1933,82,-1932</points>
<connection>
<GID>6558</GID>
<name>OUT_0</name></connection>
<intersection>-1932 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>82,-1914.5,82,-1913.5</points>
<connection>
<GID>6587</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>82,-1892.5,82,-1891.5</points>
<connection>
<GID>6702</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>82,-1874,82,-1873</points>
<connection>
<GID>6738</GID>
<name>OUT_0</name></connection>
<intersection>-1873 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>82,-1855,82,-1854</points>
<connection>
<GID>6774</GID>
<name>OUT_0</name></connection>
<intersection>-1854 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>82,-1836.5,82,-1835.5</points>
<connection>
<GID>6810</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-1985.5,89.5,-1820.5</points>
<connection>
<GID>6619</GID>
<name>N_in1</name></connection>
<connection>
<GID>6604</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 13</intersection>
<intersection>-1942 12</intersection>
<intersection>-1923 11</intersection>
<intersection>-1904.5 10</intersection>
<intersection>-1882.5 9</intersection>
<intersection>-1864 8</intersection>
<intersection>-1845 7</intersection>
<intersection>-1826.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-1826.5,94,-1826.5</points>
<connection>
<GID>6812</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-1845,94,-1845</points>
<connection>
<GID>6776</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89.5,-1864,94,-1864</points>
<connection>
<GID>6740</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-1882.5,94,-1882.5</points>
<connection>
<GID>6704</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>89.5,-1904.5,94,-1904.5</points>
<connection>
<GID>6588</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89.5,-1923,94,-1923</points>
<connection>
<GID>6561</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>89.5,-1942,94,-1942</points>
<connection>
<GID>6521</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>89.5,-1960.5,94,-1960.5</points>
<connection>
<GID>6848</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-1985.5,110.5,-1821</points>
<connection>
<GID>6620</GID>
<name>N_in1</name></connection>
<connection>
<GID>6605</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 6</intersection>
<intersection>-1951 7</intersection>
<intersection>-1932 8</intersection>
<intersection>-1913.5 9</intersection>
<intersection>-1891.5 10</intersection>
<intersection>-1873 11</intersection>
<intersection>-1854 12</intersection>
<intersection>-1835.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>107,-1969.5,110.5,-1969.5</points>
<intersection>107 14</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>107,-1951,110.5,-1951</points>
<intersection>107 15</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>107,-1932,110.5,-1932</points>
<intersection>107 16</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>107,-1913.5,110.5,-1913.5</points>
<intersection>107 17</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>107,-1891.5,110.5,-1891.5</points>
<intersection>107 20</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>107,-1873,110.5,-1873</points>
<intersection>107 21</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>107,-1854,110.5,-1854</points>
<intersection>107 22</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>107,-1835.5,110.5,-1835.5</points>
<intersection>107 23</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>107,-1970.5,107,-1969.5</points>
<connection>
<GID>6850</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>107,-1952,107,-1951</points>
<connection>
<GID>6523</GID>
<name>OUT_0</name></connection>
<intersection>-1951 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>107,-1933,107,-1932</points>
<connection>
<GID>6563</GID>
<name>OUT_0</name></connection>
<intersection>-1932 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>107,-1914.5,107,-1913.5</points>
<connection>
<GID>6589</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>107,-1892.5,107,-1891.5</points>
<connection>
<GID>6706</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>107,-1874,107,-1873</points>
<connection>
<GID>6742</GID>
<name>OUT_0</name></connection>
<intersection>-1873 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>107,-1855,107,-1854</points>
<connection>
<GID>6778</GID>
<name>OUT_0</name></connection>
<intersection>-1854 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>107,-1836.5,107,-1835.5</points>
<connection>
<GID>6814</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-1985.5,114.5,-1820.5</points>
<connection>
<GID>6621</GID>
<name>N_in1</name></connection>
<connection>
<GID>6606</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 13</intersection>
<intersection>-1942 12</intersection>
<intersection>-1923 11</intersection>
<intersection>-1904.5 10</intersection>
<intersection>-1882.5 9</intersection>
<intersection>-1864 8</intersection>
<intersection>-1845 7</intersection>
<intersection>-1826.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>114.5,-1826.5,117,-1826.5</points>
<connection>
<GID>6816</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-1845,117,-1845</points>
<connection>
<GID>6780</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-1864,117,-1864</points>
<connection>
<GID>6744</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114.5,-1882.5,117,-1882.5</points>
<connection>
<GID>6708</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114.5,-1904.5,117,-1904.5</points>
<connection>
<GID>6590</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>114.5,-1923,117,-1923</points>
<connection>
<GID>6566</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114.5,-1942,117,-1942</points>
<connection>
<GID>6525</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>114.5,-1960.5,117,-1960.5</points>
<connection>
<GID>6489</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1985.5,133,-1820.5</points>
<connection>
<GID>6622</GID>
<name>N_in1</name></connection>
<connection>
<GID>6607</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 6</intersection>
<intersection>-1951 7</intersection>
<intersection>-1932 8</intersection>
<intersection>-1913.5 9</intersection>
<intersection>-1891.5 10</intersection>
<intersection>-1873 11</intersection>
<intersection>-1854 12</intersection>
<intersection>-1835.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>130,-1969.5,133,-1969.5</points>
<intersection>130 14</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-1951,133,-1951</points>
<intersection>130 15</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>130,-1932,133,-1932</points>
<intersection>130 16</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>130,-1913.5,133,-1913.5</points>
<intersection>130 17</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>130,-1891.5,133,-1891.5</points>
<intersection>130 20</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>130,-1873,133,-1873</points>
<intersection>130 21</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>130,-1854,133,-1854</points>
<intersection>130 22</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>130,-1835.5,133,-1835.5</points>
<intersection>130 23</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>130,-1970.5,130,-1969.5</points>
<connection>
<GID>6491</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>130,-1952,130,-1951</points>
<connection>
<GID>6527</GID>
<name>OUT_0</name></connection>
<intersection>-1951 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>130,-1933,130,-1932</points>
<connection>
<GID>6568</GID>
<name>OUT_0</name></connection>
<intersection>-1932 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>130,-1914.5,130,-1913.5</points>
<connection>
<GID>6591</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>130,-1892.5,130,-1891.5</points>
<connection>
<GID>6710</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>130,-1874,130,-1873</points>
<connection>
<GID>6746</GID>
<name>OUT_0</name></connection>
<intersection>-1873 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>130,-1855,130,-1854</points>
<connection>
<GID>6782</GID>
<name>OUT_0</name></connection>
<intersection>-1854 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>130,-1836.5,130,-1835.5</points>
<connection>
<GID>6818</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-1985.5,137,-1820.5</points>
<connection>
<GID>6623</GID>
<name>N_in1</name></connection>
<connection>
<GID>6608</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 13</intersection>
<intersection>-1942 12</intersection>
<intersection>-1923 11</intersection>
<intersection>-1904.5 10</intersection>
<intersection>-1882.5 9</intersection>
<intersection>-1864 8</intersection>
<intersection>-1845 7</intersection>
<intersection>-1826.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>137,-1826.5,140,-1826.5</points>
<connection>
<GID>6820</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137,-1845,140,-1845</points>
<connection>
<GID>6784</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-1864,140,-1864</points>
<connection>
<GID>6748</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137,-1882.5,140,-1882.5</points>
<connection>
<GID>6712</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-1904.5,140,-1904.5</points>
<connection>
<GID>6592</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>137,-1923,140,-1923</points>
<connection>
<GID>6571</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137,-1942,140,-1942</points>
<connection>
<GID>6529</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-1960.5,140,-1960.5</points>
<connection>
<GID>6493</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>4685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-1985,156,-1820.5</points>
<connection>
<GID>6624</GID>
<name>N_in1</name></connection>
<connection>
<GID>6609</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 6</intersection>
<intersection>-1951 7</intersection>
<intersection>-1932 8</intersection>
<intersection>-1913.5 9</intersection>
<intersection>-1891.5 10</intersection>
<intersection>-1873 11</intersection>
<intersection>-1854 12</intersection>
<intersection>-1835.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>153,-1969.5,156,-1969.5</points>
<intersection>153 14</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>153,-1951,156,-1951</points>
<intersection>153 15</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>153,-1932,156,-1932</points>
<intersection>153 16</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>153,-1913.5,156,-1913.5</points>
<intersection>153 17</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>153,-1891.5,156,-1891.5</points>
<intersection>153 20</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>153,-1873,156,-1873</points>
<intersection>153 21</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>153,-1854,156,-1854</points>
<intersection>153 22</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>153,-1835.5,156,-1835.5</points>
<intersection>153 23</intersection>
<intersection>156 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>153,-1970.5,153,-1969.5</points>
<connection>
<GID>6495</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>153,-1952,153,-1951</points>
<connection>
<GID>6531</GID>
<name>OUT_0</name></connection>
<intersection>-1951 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>153,-1933,153,-1932</points>
<connection>
<GID>6573</GID>
<name>OUT_0</name></connection>
<intersection>-1932 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>153,-1914.5,153,-1913.5</points>
<connection>
<GID>6593</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>153,-1892.5,153,-1891.5</points>
<connection>
<GID>6714</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>153,-1874,153,-1873</points>
<connection>
<GID>6750</GID>
<name>OUT_0</name></connection>
<intersection>-1873 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>153,-1855,153,-1854</points>
<connection>
<GID>6786</GID>
<name>OUT_0</name></connection>
<intersection>-1854 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>153,-1836.5,153,-1835.5</points>
<connection>
<GID>6822</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-1985,161,-1820.5</points>
<connection>
<GID>6625</GID>
<name>N_in1</name></connection>
<connection>
<GID>6610</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 13</intersection>
<intersection>-1942 12</intersection>
<intersection>-1923 11</intersection>
<intersection>-1904.5 10</intersection>
<intersection>-1882.5 9</intersection>
<intersection>-1864 8</intersection>
<intersection>-1845 7</intersection>
<intersection>-1826.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>161,-1826.5,163,-1826.5</points>
<connection>
<GID>6824</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>161,-1845,163,-1845</points>
<connection>
<GID>6788</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>161,-1864,163,-1864</points>
<connection>
<GID>6752</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>161,-1882.5,163,-1882.5</points>
<connection>
<GID>6716</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>161,-1904.5,163,-1904.5</points>
<connection>
<GID>6594</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>161,-1923,163,-1923</points>
<connection>
<GID>6575</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>161,-1942,163,-1942</points>
<connection>
<GID>6533</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>161,-1960.5,163,-1960.5</points>
<connection>
<GID>6497</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>4687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-1984.5,179,-1820.5</points>
<connection>
<GID>6626</GID>
<name>N_in1</name></connection>
<connection>
<GID>6612</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 16</intersection>
<intersection>-1951 15</intersection>
<intersection>-1932 14</intersection>
<intersection>-1913.5 13</intersection>
<intersection>-1891.5 12</intersection>
<intersection>-1873 11</intersection>
<intersection>-1854 10</intersection>
<intersection>-1835.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>176,-1835.5,179,-1835.5</points>
<intersection>176 26</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>176,-1854,179,-1854</points>
<intersection>176 25</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>176,-1873,179,-1873</points>
<intersection>176 24</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>176,-1891.5,179,-1891.5</points>
<intersection>176 23</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>176,-1913.5,179,-1913.5</points>
<intersection>176 20</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>176,-1932,179,-1932</points>
<intersection>176 19</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>176,-1951,179,-1951</points>
<intersection>176 18</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>176,-1969.5,179,-1969.5</points>
<intersection>176 17</intersection>
<intersection>179 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>176,-1970.5,176,-1969.5</points>
<connection>
<GID>6499</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>176,-1952,176,-1951</points>
<connection>
<GID>6535</GID>
<name>OUT_0</name></connection>
<intersection>-1951 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>176,-1933,176,-1932</points>
<connection>
<GID>6576</GID>
<name>OUT_0</name></connection>
<intersection>-1932 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>176,-1914.5,176,-1913.5</points>
<connection>
<GID>6595</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>176,-1892.5,176,-1891.5</points>
<connection>
<GID>6718</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>176,-1874,176,-1873</points>
<connection>
<GID>6754</GID>
<name>OUT_0</name></connection>
<intersection>-1873 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>176,-1855,176,-1854</points>
<connection>
<GID>6790</GID>
<name>OUT_0</name></connection>
<intersection>-1854 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>176,-1836.5,176,-1835.5</points>
<connection>
<GID>6826</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>4688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-1984.5,183.5,-1820.5</points>
<connection>
<GID>6627</GID>
<name>N_in1</name></connection>
<connection>
<GID>6611</GID>
<name>N_in0</name></connection>
<intersection>-1960.5 13</intersection>
<intersection>-1942 12</intersection>
<intersection>-1923 11</intersection>
<intersection>-1904.5 10</intersection>
<intersection>-1882.5 9</intersection>
<intersection>-1864 8</intersection>
<intersection>-1845 7</intersection>
<intersection>-1826.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>183.5,-1826.5,188,-1826.5</points>
<connection>
<GID>6828</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>183.5,-1845,188,-1845</points>
<connection>
<GID>6792</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>183.5,-1864,188,-1864</points>
<connection>
<GID>6756</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>183.5,-1882.5,188,-1882.5</points>
<connection>
<GID>6720</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183.5,-1904.5,188,-1904.5</points>
<connection>
<GID>6596</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183.5,-1923,188,-1923</points>
<connection>
<GID>6578</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183.5,-1942,188,-1942</points>
<connection>
<GID>6537</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183.5,-1960.5,188,-1960.5</points>
<connection>
<GID>6501</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-1984,204.5,-1821</points>
<connection>
<GID>6628</GID>
<name>N_in1</name></connection>
<connection>
<GID>6613</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 6</intersection>
<intersection>-1951 7</intersection>
<intersection>-1932 8</intersection>
<intersection>-1913.5 9</intersection>
<intersection>-1891.5 10</intersection>
<intersection>-1873 11</intersection>
<intersection>-1854 12</intersection>
<intersection>-1835.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>201,-1969.5,204.5,-1969.5</points>
<intersection>201 14</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>201,-1951,204.5,-1951</points>
<intersection>201 15</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>201,-1932,204.5,-1932</points>
<intersection>201 16</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>201,-1913.5,204.5,-1913.5</points>
<intersection>201 17</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>201,-1891.5,204.5,-1891.5</points>
<intersection>201 20</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>201,-1873,204.5,-1873</points>
<intersection>201 21</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>201,-1854,204.5,-1854</points>
<intersection>201 22</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>201,-1835.5,204.5,-1835.5</points>
<intersection>201 23</intersection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>201,-1970.5,201,-1969.5</points>
<connection>
<GID>6503</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201,-1952,201,-1951</points>
<connection>
<GID>6539</GID>
<name>OUT_0</name></connection>
<intersection>-1951 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>201,-1933,201,-1932</points>
<connection>
<GID>6579</GID>
<name>OUT_0</name></connection>
<intersection>-1932 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>201,-1914.5,201,-1913.5</points>
<connection>
<GID>6597</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>201,-1892.5,201,-1891.5</points>
<connection>
<GID>6722</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>201,-1874,201,-1873</points>
<connection>
<GID>6758</GID>
<name>OUT_0</name></connection>
<intersection>-1873 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>201,-1855,201,-1854</points>
<connection>
<GID>6794</GID>
<name>OUT_0</name></connection>
<intersection>-1854 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>201,-1836.5,201,-1835.5</points>
<connection>
<GID>6830</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-1984,208,-1821</points>
<connection>
<GID>6630</GID>
<name>N_in0</name></connection>
<connection>
<GID>6629</GID>
<name>N_in1</name></connection>
<intersection>-1960.5 11</intersection>
<intersection>-1942 10</intersection>
<intersection>-1923 9</intersection>
<intersection>-1904.5 7</intersection>
<intersection>-1882.5 6</intersection>
<intersection>-1864 5</intersection>
<intersection>-1845 4</intersection>
<intersection>-1826.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208,-1826.5,211,-1826.5</points>
<connection>
<GID>6832</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208,-1845,211,-1845</points>
<connection>
<GID>6796</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>208,-1864,211,-1864</points>
<connection>
<GID>6760</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>208,-1882.5,211,-1882.5</points>
<connection>
<GID>6724</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>208,-1904.5,211,-1904.5</points>
<connection>
<GID>6598</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>208,-1923,211,-1923</points>
<connection>
<GID>6580</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>208,-1942,211,-1942</points>
<connection>
<GID>6541</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>208,-1960.5,211,-1960.5</points>
<connection>
<GID>6505</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>4691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-1984,229,-1822</points>
<connection>
<GID>6631</GID>
<name>N_in1</name></connection>
<connection>
<GID>6614</GID>
<name>N_in0</name></connection>
<intersection>-1969.5 11</intersection>
<intersection>-1951 10</intersection>
<intersection>-1932 9</intersection>
<intersection>-1913.5 8</intersection>
<intersection>-1891.5 7</intersection>
<intersection>-1873 6</intersection>
<intersection>-1854 5</intersection>
<intersection>-1835.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>224,-1835.5,229,-1835.5</points>
<intersection>224 21</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>224,-1854,229,-1854</points>
<intersection>224 20</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>224,-1873,229,-1873</points>
<intersection>224 19</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>224,-1891.5,229,-1891.5</points>
<intersection>224 18</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>224,-1913.5,229,-1913.5</points>
<intersection>224 15</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>224,-1932,229,-1932</points>
<intersection>224 14</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>224,-1951,229,-1951</points>
<intersection>224 13</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>224,-1969.5,229,-1969.5</points>
<intersection>224 12</intersection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>224,-1970.5,224,-1969.5</points>
<connection>
<GID>6507</GID>
<name>OUT_0</name></connection>
<intersection>-1969.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>224,-1952,224,-1951</points>
<connection>
<GID>6543</GID>
<name>OUT_0</name></connection>
<intersection>-1951 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>224,-1933,224,-1932</points>
<connection>
<GID>6581</GID>
<name>OUT_0</name></connection>
<intersection>-1932 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>224,-1914.5,224,-1913.5</points>
<connection>
<GID>6599</GID>
<name>OUT_0</name></connection>
<intersection>-1913.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>224,-1892.5,224,-1891.5</points>
<connection>
<GID>6726</GID>
<name>OUT_0</name></connection>
<intersection>-1891.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>224,-1874,224,-1873</points>
<connection>
<GID>6762</GID>
<name>OUT_0</name></connection>
<intersection>-1873 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>224,-1855,224,-1854</points>
<connection>
<GID>6798</GID>
<name>OUT_0</name></connection>
<intersection>-1854 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>224,-1836.5,224,-1835.5</points>
<connection>
<GID>6834</GID>
<name>OUT_0</name></connection>
<intersection>-1835.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>4692</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-128,-1828.5,18.5,-1828.5</points>
<connection>
<GID>6800</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-1980,-128,-1828.5</points>
<connection>
<GID>6637</GID>
<name>OUT_15</name></connection>
<intersection>-1838 4</intersection>
<intersection>-1828.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-1838,30,-1838</points>
<connection>
<GID>6802</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>4693</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-127,-1847,18.5,-1847</points>
<connection>
<GID>6764</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-127,-1981,-127,-1847</points>
<intersection>-1981 6</intersection>
<intersection>-1856.5 5</intersection>
<intersection>-1847 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-127,-1856.5,30,-1856.5</points>
<connection>
<GID>6766</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-1981,-127,-1981</points>
<connection>
<GID>6637</GID>
<name>OUT_14</name></connection>
<intersection>-127 4</intersection></hsegment></shape></wire>
<wire>
<ID>4694</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-126,-1866,18.5,-1866</points>
<connection>
<GID>6728</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-1982,-126,-1866</points>
<intersection>-1982 6</intersection>
<intersection>-1875.5 4</intersection>
<intersection>-1866 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-1875.5,30,-1875.5</points>
<connection>
<GID>6730</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-1982,-126,-1982</points>
<connection>
<GID>6637</GID>
<name>OUT_13</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>4695</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-125,-1884.5,18.5,-1884.5</points>
<connection>
<GID>6668</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-125,-1983,-125,-1884.5</points>
<intersection>-1983 5</intersection>
<intersection>-1894 4</intersection>
<intersection>-1884.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-125,-1894,30,-1894</points>
<connection>
<GID>6673</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1983,-125,-1983</points>
<connection>
<GID>6637</GID>
<name>OUT_12</name></connection>
<intersection>-125 3</intersection></hsegment></shape></wire>
<wire>
<ID>4696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,-1906.5,18.5,-1906.5</points>
<connection>
<GID>6582</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-1984,-124,-1906.5</points>
<intersection>-1984 6</intersection>
<intersection>-1916 4</intersection>
<intersection>-1906.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-1916,29.5,-1916</points>
<connection>
<GID>6583</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-1984,-124,-1984</points>
<connection>
<GID>6637</GID>
<name>OUT_11</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>4697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123,-1925,18.5,-1925</points>
<connection>
<GID>6546</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-1985,-123,-1925</points>
<intersection>-1985 5</intersection>
<intersection>-1934.5 4</intersection>
<intersection>-1925 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-1934.5,29.5,-1934.5</points>
<connection>
<GID>6548</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1985,-123,-1985</points>
<connection>
<GID>6637</GID>
<name>OUT_10</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>4698</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-1944,18.5,-1944</points>
<connection>
<GID>6509</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-1986,-122,-1944</points>
<intersection>-1986 5</intersection>
<intersection>-1953.5 4</intersection>
<intersection>-1944 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-1953.5,29.5,-1953.5</points>
<connection>
<GID>6511</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1986,-122,-1986</points>
<connection>
<GID>6637</GID>
<name>OUT_9</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>4699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-1962.5,18.5,-1962.5</points>
<connection>
<GID>6836</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-1987,-121,-1962.5</points>
<intersection>-1987 5</intersection>
<intersection>-1972 4</intersection>
<intersection>-1962.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-1972,29.5,-1972</points>
<connection>
<GID>6838</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1987,-121,-1987</points>
<connection>
<GID>6637</GID>
<name>OUT_8</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-1986,17.5,-1821</points>
<connection>
<GID>6635</GID>
<name>N_in1</name></connection>
<connection>
<GID>6633</GID>
<name>N_in0</name></connection>
<intersection>-1964.5 10</intersection>
<intersection>-1946 9</intersection>
<intersection>-1927 8</intersection>
<intersection>-1908.5 7</intersection>
<intersection>-1886.5 6</intersection>
<intersection>-1868 5</intersection>
<intersection>-1849 4</intersection>
<intersection>-1830.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-1830.5,18.5,-1830.5</points>
<connection>
<GID>6800</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-1849,18.5,-1849</points>
<connection>
<GID>6764</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>17.5,-1868,18.5,-1868</points>
<connection>
<GID>6728</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>17.5,-1886.5,18.5,-1886.5</points>
<connection>
<GID>6668</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>17.5,-1908.5,18.5,-1908.5</points>
<connection>
<GID>6582</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>17.5,-1927,18.5,-1927</points>
<connection>
<GID>6546</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>17.5,-1946,18.5,-1946</points>
<connection>
<GID>6509</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>17.5,-1964.5,18.5,-1964.5</points>
<connection>
<GID>6836</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-1986,27.5,-1821</points>
<connection>
<GID>6634</GID>
<name>N_in1</name></connection>
<connection>
<GID>6632</GID>
<name>N_in0</name></connection>
<intersection>-1974 3</intersection>
<intersection>-1955.5 5</intersection>
<intersection>-1936.5 7</intersection>
<intersection>-1918 9</intersection>
<intersection>-1896 11</intersection>
<intersection>-1877.5 13</intersection>
<intersection>-1858.5 15</intersection>
<intersection>-1840 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-1974,29.5,-1974</points>
<connection>
<GID>6838</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-1955.5,29.5,-1955.5</points>
<connection>
<GID>6511</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-1936.5,29.5,-1936.5</points>
<connection>
<GID>6548</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>27.5,-1918,29.5,-1918</points>
<connection>
<GID>6583</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>27.5,-1896,30,-1896</points>
<connection>
<GID>6673</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>27.5,-1877.5,30,-1877.5</points>
<connection>
<GID>6730</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>27.5,-1858.5,30,-1858.5</points>
<connection>
<GID>6766</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>27.5,-1840,30,-1840</points>
<connection>
<GID>6802</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4702</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2073.5,59,-2073.5</points>
<connection>
<GID>6733</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2073.5,53,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2058,53,-2058</points>
<connection>
<GID>6721</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2073.5,82,-2073.5</points>
<connection>
<GID>6759</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2073.5,76,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2058,76,-2058</points>
<connection>
<GID>6757</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4704</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2073.5,107,-2073.5</points>
<connection>
<GID>6767</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2073.5,101,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2058,101,-2058</points>
<connection>
<GID>6763</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2073.5,130,-2073.5</points>
<connection>
<GID>6775</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2073.5,124,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2058,124,-2058</points>
<connection>
<GID>6771</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4706</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2073.5,153,-2073.5</points>
<connection>
<GID>6781</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2073.5,147,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2058,147,-2058</points>
<connection>
<GID>6777</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4707</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2073.5,176,-2073.5</points>
<connection>
<GID>6785</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2073.5,170,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2058,170,-2058</points>
<connection>
<GID>6783</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4708</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2073.5,201,-2073.5</points>
<connection>
<GID>6789</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2073.5,195,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2058,195,-2058</points>
<connection>
<GID>6787</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4709</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2073.5,224,-2073.5</points>
<connection>
<GID>6793</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2073.5,218,-2058</points>
<intersection>-2073.5 1</intersection>
<intersection>-2058 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2058,218,-2058</points>
<connection>
<GID>6791</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4710</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2061,211,-2061</points>
<connection>
<GID>6715</GID>
<name>OUT</name></connection>
<connection>
<GID>6721</GID>
<name>clock</name></connection>
<connection>
<GID>6757</GID>
<name>clock</name></connection>
<connection>
<GID>6763</GID>
<name>clock</name></connection>
<connection>
<GID>6771</GID>
<name>clock</name></connection>
<connection>
<GID>6777</GID>
<name>clock</name></connection>
<connection>
<GID>6783</GID>
<name>clock</name></connection>
<connection>
<GID>6787</GID>
<name>clock</name></connection>
<connection>
<GID>6791</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4711</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2070.5,222,-2070.5</points>
<connection>
<GID>6717</GID>
<name>OUT</name></connection>
<connection>
<GID>6733</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6759</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6767</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6775</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6781</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6785</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6789</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6793</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4712</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2055,59,-2055</points>
<connection>
<GID>6801</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2055,53,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2039.5,53,-2039.5</points>
<connection>
<GID>6799</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2055,82,-2055</points>
<connection>
<GID>6805</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2055,76,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2039.5,76,-2039.5</points>
<connection>
<GID>6803</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4714</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2055,107,-2055</points>
<connection>
<GID>6809</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2055,101,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2039.5,101,-2039.5</points>
<connection>
<GID>6807</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4715</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2055,130,-2055</points>
<connection>
<GID>6813</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2055,124,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2039.5,124,-2039.5</points>
<connection>
<GID>6811</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4716</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2055,153,-2055</points>
<connection>
<GID>6817</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2055,147,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2039.5,147,-2039.5</points>
<connection>
<GID>6815</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4717</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2055,176,-2055</points>
<connection>
<GID>6821</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2055,170,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2039.5,170,-2039.5</points>
<connection>
<GID>6819</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2055,201,-2055</points>
<connection>
<GID>6825</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2055,195,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2039.5,195,-2039.5</points>
<connection>
<GID>6823</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4719</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2055,224,-2055</points>
<connection>
<GID>6829</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2055,218,-2039.5</points>
<intersection>-2055 1</intersection>
<intersection>-2039.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2039.5,218,-2039.5</points>
<connection>
<GID>6827</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4720</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2042.5,211,-2042.5</points>
<connection>
<GID>6795</GID>
<name>OUT</name></connection>
<connection>
<GID>6799</GID>
<name>clock</name></connection>
<connection>
<GID>6803</GID>
<name>clock</name></connection>
<connection>
<GID>6807</GID>
<name>clock</name></connection>
<connection>
<GID>6811</GID>
<name>clock</name></connection>
<connection>
<GID>6815</GID>
<name>clock</name></connection>
<connection>
<GID>6819</GID>
<name>clock</name></connection>
<connection>
<GID>6823</GID>
<name>clock</name></connection>
<connection>
<GID>6827</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1642</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-247.5,220,-247.5</points>
<connection>
<GID>1685</GID>
<name>clock</name></connection>
<connection>
<GID>1683</GID>
<name>clock</name></connection>
<connection>
<GID>1681</GID>
<name>clock</name></connection>
<connection>
<GID>1679</GID>
<name>clock</name></connection>
<connection>
<GID>1677</GID>
<name>clock</name></connection>
<connection>
<GID>1675</GID>
<name>clock</name></connection>
<connection>
<GID>1673</GID>
<name>clock</name></connection>
<connection>
<GID>1671</GID>
<name>clock</name></connection>
<connection>
<GID>1669</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2052,222,-2052</points>
<connection>
<GID>6797</GID>
<name>OUT</name></connection>
<connection>
<GID>6801</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6805</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6809</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6813</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6817</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6821</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6825</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6829</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1643</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-257,231,-257</points>
<connection>
<GID>1686</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1684</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1682</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1678</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1676</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1674</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1672</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1670</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4722</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2036,59,-2036</points>
<connection>
<GID>6837</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2036,53,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2020.5,53,-2020.5</points>
<connection>
<GID>6835</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>1644</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-241,68,-241</points>
<connection>
<GID>1959</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-241,62,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61,-225.5,62,-225.5</points>
<connection>
<GID>1957</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>4723</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2036,82,-2036</points>
<connection>
<GID>6841</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2036,76,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2020.5,76,-2020.5</points>
<connection>
<GID>6839</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>1645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-241,91,-241</points>
<connection>
<GID>1963</GID>
<name>IN_0</name></connection>
<intersection>85 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85,-241,85,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-225.5,85,-225.5</points>
<connection>
<GID>1961</GID>
<name>OUT_0</name></connection>
<intersection>85 2</intersection></hsegment></shape></wire>
<wire>
<ID>4724</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2036,107,-2036</points>
<connection>
<GID>6845</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2036,101,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2020.5,101,-2020.5</points>
<connection>
<GID>6843</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>1646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-241,116,-241</points>
<connection>
<GID>1967</GID>
<name>IN_0</name></connection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,-241,110,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109,-225.5,110,-225.5</points>
<connection>
<GID>1965</GID>
<name>OUT_0</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>4725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2036,130,-2036</points>
<connection>
<GID>6849</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2036,124,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2020.5,124,-2020.5</points>
<connection>
<GID>6847</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>1647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-241,139,-241</points>
<connection>
<GID>2204</GID>
<name>IN_0</name></connection>
<intersection>133 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133,-241,133,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132,-225.5,133,-225.5</points>
<connection>
<GID>1969</GID>
<name>OUT_0</name></connection>
<intersection>133 2</intersection></hsegment></shape></wire>
<wire>
<ID>4726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2036,153,-2036</points>
<connection>
<GID>6490</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2036,147,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2020.5,147,-2020.5</points>
<connection>
<GID>6851</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>1648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-241,162,-241</points>
<connection>
<GID>2206</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-241,156,-225.5</points>
<intersection>-241 1</intersection>
<intersection>-225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>155,-225.5,156,-225.5</points>
<connection>
<GID>2205</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>4727</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2036,176,-2036</points>
<connection>
<GID>6494</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2036,170,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2020.5,170,-2020.5</points>
<connection>
<GID>6492</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4728</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2036,201,-2036</points>
<connection>
<GID>6498</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2036,195,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2020.5,195,-2020.5</points>
<connection>
<GID>6496</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4729</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2036,224,-2036</points>
<connection>
<GID>6502</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2036,218,-2020.5</points>
<intersection>-2036 1</intersection>
<intersection>-2020.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2020.5,218,-2020.5</points>
<connection>
<GID>6500</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2023.5,211,-2023.5</points>
<connection>
<GID>6851</GID>
<name>clock</name></connection>
<connection>
<GID>6847</GID>
<name>clock</name></connection>
<connection>
<GID>6843</GID>
<name>clock</name></connection>
<connection>
<GID>6839</GID>
<name>clock</name></connection>
<connection>
<GID>6835</GID>
<name>clock</name></connection>
<connection>
<GID>6831</GID>
<name>OUT</name></connection>
<connection>
<GID>6500</GID>
<name>clock</name></connection>
<connection>
<GID>6496</GID>
<name>clock</name></connection>
<connection>
<GID>6492</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4731</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2033,222,-2033</points>
<connection>
<GID>6849</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6845</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6841</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6837</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6833</GID>
<name>OUT</name></connection>
<connection>
<GID>6502</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6498</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6494</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6490</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4732</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2017.5,59,-2017.5</points>
<connection>
<GID>6510</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2017.5,53,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2002,53,-2002</points>
<connection>
<GID>6508</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4733</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2017.5,82,-2017.5</points>
<connection>
<GID>6514</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2017.5,76,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2002,76,-2002</points>
<connection>
<GID>6512</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2017.5,107,-2017.5</points>
<connection>
<GID>6518</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2017.5,101,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2002,101,-2002</points>
<connection>
<GID>6516</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4735</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2017.5,130,-2017.5</points>
<connection>
<GID>6522</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2017.5,124,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2002,124,-2002</points>
<connection>
<GID>6520</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4736</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2017.5,153,-2017.5</points>
<connection>
<GID>6526</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2017.5,147,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2002,147,-2002</points>
<connection>
<GID>6524</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4737</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2017.5,176,-2017.5</points>
<connection>
<GID>6530</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2017.5,170,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2002,170,-2002</points>
<connection>
<GID>6528</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2017.5,201,-2017.5</points>
<connection>
<GID>6534</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2017.5,195,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2002,195,-2002</points>
<connection>
<GID>6532</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2017.5,224,-2017.5</points>
<connection>
<GID>6538</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2017.5,218,-2002</points>
<intersection>-2017.5 1</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2002,218,-2002</points>
<connection>
<GID>6536</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4740</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2005,211,-2005</points>
<connection>
<GID>6504</GID>
<name>OUT</name></connection>
<connection>
<GID>6508</GID>
<name>clock</name></connection>
<connection>
<GID>6512</GID>
<name>clock</name></connection>
<connection>
<GID>6516</GID>
<name>clock</name></connection>
<connection>
<GID>6520</GID>
<name>clock</name></connection>
<connection>
<GID>6524</GID>
<name>clock</name></connection>
<connection>
<GID>6528</GID>
<name>clock</name></connection>
<connection>
<GID>6532</GID>
<name>clock</name></connection>
<connection>
<GID>6536</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2014.5,222,-2014.5</points>
<connection>
<GID>6506</GID>
<name>OUT</name></connection>
<connection>
<GID>6510</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6514</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6518</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6522</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6526</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6530</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6534</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6538</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2151.5,59,-2151.5</points>
<connection>
<GID>6547</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2151.5,53,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2136,53,-2136</points>
<connection>
<GID>6544</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4743</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2151.5,82,-2151.5</points>
<connection>
<GID>6552</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2151.5,76,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2136,76,-2136</points>
<connection>
<GID>6549</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2151.5,107,-2151.5</points>
<connection>
<GID>6557</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2151.5,101,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2136,101,-2136</points>
<connection>
<GID>6554</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4745</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2151.5,130,-2151.5</points>
<connection>
<GID>6562</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2151.5,124,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2136,124,-2136</points>
<connection>
<GID>6559</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4746</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2151.5,153,-2151.5</points>
<connection>
<GID>6567</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2151.5,147,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2136,147,-2136</points>
<connection>
<GID>6564</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4747</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2151.5,176,-2151.5</points>
<connection>
<GID>6572</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2151.5,170,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2136,170,-2136</points>
<connection>
<GID>6569</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4748</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2151.5,201,-2151.5</points>
<connection>
<GID>6639</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2151.5,195,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2136,195,-2136</points>
<connection>
<GID>6638</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4749</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2151.5,224,-2151.5</points>
<connection>
<GID>6641</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2151.5,218,-2136</points>
<intersection>-2151.5 1</intersection>
<intersection>-2136 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2136,218,-2136</points>
<connection>
<GID>6640</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4750</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2139,211,-2139</points>
<connection>
<GID>6540</GID>
<name>OUT</name></connection>
<connection>
<GID>6544</GID>
<name>clock</name></connection>
<connection>
<GID>6549</GID>
<name>clock</name></connection>
<connection>
<GID>6554</GID>
<name>clock</name></connection>
<connection>
<GID>6559</GID>
<name>clock</name></connection>
<connection>
<GID>6564</GID>
<name>clock</name></connection>
<connection>
<GID>6569</GID>
<name>clock</name></connection>
<connection>
<GID>6638</GID>
<name>clock</name></connection>
<connection>
<GID>6640</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4751</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2148.5,222,-2148.5</points>
<connection>
<GID>6542</GID>
<name>OUT</name></connection>
<connection>
<GID>6547</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6552</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6557</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6562</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6567</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6572</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6639</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6641</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4752</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2133,59,-2133</points>
<connection>
<GID>6645</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2133,53,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2117.5,53,-2117.5</points>
<connection>
<GID>6644</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4753</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2133,82,-2133</points>
<connection>
<GID>6647</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2133,76,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2117.5,76,-2117.5</points>
<connection>
<GID>6646</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4754</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2133,107,-2133</points>
<connection>
<GID>6649</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2133,101,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2117.5,101,-2117.5</points>
<connection>
<GID>6648</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4755</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2133,130,-2133</points>
<connection>
<GID>6651</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2133,124,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2117.5,124,-2117.5</points>
<connection>
<GID>6650</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4756</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2133,153,-2133</points>
<connection>
<GID>6653</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2133,147,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2117.5,147,-2117.5</points>
<connection>
<GID>6652</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4757</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2133,176,-2133</points>
<connection>
<GID>6655</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2133,170,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2117.5,170,-2117.5</points>
<connection>
<GID>6654</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4758</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2133,201,-2133</points>
<connection>
<GID>6657</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2133,195,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2117.5,195,-2117.5</points>
<connection>
<GID>6656</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4759</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2133,224,-2133</points>
<connection>
<GID>6659</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2133,218,-2117.5</points>
<intersection>-2133 1</intersection>
<intersection>-2117.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2117.5,218,-2117.5</points>
<connection>
<GID>6658</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4760</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2120.5,211,-2120.5</points>
<connection>
<GID>6642</GID>
<name>OUT</name></connection>
<connection>
<GID>6644</GID>
<name>clock</name></connection>
<connection>
<GID>6646</GID>
<name>clock</name></connection>
<connection>
<GID>6648</GID>
<name>clock</name></connection>
<connection>
<GID>6650</GID>
<name>clock</name></connection>
<connection>
<GID>6652</GID>
<name>clock</name></connection>
<connection>
<GID>6654</GID>
<name>clock</name></connection>
<connection>
<GID>6656</GID>
<name>clock</name></connection>
<connection>
<GID>6658</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4761</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2130,222,-2130</points>
<connection>
<GID>6643</GID>
<name>OUT</name></connection>
<connection>
<GID>6645</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6647</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6649</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6651</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6653</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6655</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6657</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6659</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4762</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2114,59,-2114</points>
<connection>
<GID>6555</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2114,53,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2098.5,53,-2098.5</points>
<connection>
<GID>6550</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4763</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2114,82,-2114</points>
<connection>
<GID>6565</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2114,76,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2098.5,76,-2098.5</points>
<connection>
<GID>6560</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4764</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2114,107,-2114</points>
<connection>
<GID>6574</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2114,101,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2098.5,101,-2098.5</points>
<connection>
<GID>6570</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4765</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2114,130,-2114</points>
<connection>
<GID>6661</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2114,124,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2098.5,124,-2098.5</points>
<connection>
<GID>6577</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2114,153,-2114</points>
<connection>
<GID>6663</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2114,147,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2098.5,147,-2098.5</points>
<connection>
<GID>6662</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4767</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2114,176,-2114</points>
<connection>
<GID>6665</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2114,170,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2098.5,170,-2098.5</points>
<connection>
<GID>6664</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4768</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2114,201,-2114</points>
<connection>
<GID>6667</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2114,195,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2098.5,195,-2098.5</points>
<connection>
<GID>6666</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2114,224,-2114</points>
<connection>
<GID>6670</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2114,218,-2098.5</points>
<intersection>-2114 1</intersection>
<intersection>-2098.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2098.5,218,-2098.5</points>
<connection>
<GID>6669</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2101.5,211,-2101.5</points>
<connection>
<GID>6669</GID>
<name>clock</name></connection>
<connection>
<GID>6666</GID>
<name>clock</name></connection>
<connection>
<GID>6664</GID>
<name>clock</name></connection>
<connection>
<GID>6662</GID>
<name>clock</name></connection>
<connection>
<GID>6660</GID>
<name>OUT</name></connection>
<connection>
<GID>6577</GID>
<name>clock</name></connection>
<connection>
<GID>6570</GID>
<name>clock</name></connection>
<connection>
<GID>6560</GID>
<name>clock</name></connection>
<connection>
<GID>6550</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4771</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2111,222,-2111</points>
<connection>
<GID>6545</GID>
<name>OUT</name></connection>
<connection>
<GID>6555</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6565</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6574</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6661</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6663</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6665</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6667</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6670</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4772</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2095.5,59,-2095.5</points>
<connection>
<GID>6675</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2095.5,53,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2080,53,-2080</points>
<connection>
<GID>6674</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4773</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2095.5,82,-2095.5</points>
<connection>
<GID>6677</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2095.5,76,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2080,76,-2080</points>
<connection>
<GID>6676</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4774</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2095.5,107,-2095.5</points>
<connection>
<GID>6680</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2095.5,101,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2080,101,-2080</points>
<connection>
<GID>6679</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4775</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2095.5,130,-2095.5</points>
<connection>
<GID>6682</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2095.5,124,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2080,124,-2080</points>
<connection>
<GID>6681</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4776</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2095.5,153,-2095.5</points>
<connection>
<GID>6685</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2095.5,147,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2080,147,-2080</points>
<connection>
<GID>6683</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4777</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2095.5,176,-2095.5</points>
<connection>
<GID>6687</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2095.5,170,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2080,170,-2080</points>
<connection>
<GID>6686</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4778</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2095.5,201,-2095.5</points>
<connection>
<GID>6689</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2095.5,195,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2080,195,-2080</points>
<connection>
<GID>6688</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4779</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2095.5,224,-2095.5</points>
<connection>
<GID>6691</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2095.5,218,-2080</points>
<intersection>-2095.5 1</intersection>
<intersection>-2080 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2080,218,-2080</points>
<connection>
<GID>6690</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4780</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2083,211,-2083</points>
<connection>
<GID>6671</GID>
<name>OUT</name></connection>
<connection>
<GID>6674</GID>
<name>clock</name></connection>
<connection>
<GID>6676</GID>
<name>clock</name></connection>
<connection>
<GID>6679</GID>
<name>clock</name></connection>
<connection>
<GID>6681</GID>
<name>clock</name></connection>
<connection>
<GID>6683</GID>
<name>clock</name></connection>
<connection>
<GID>6686</GID>
<name>clock</name></connection>
<connection>
<GID>6688</GID>
<name>clock</name></connection>
<connection>
<GID>6690</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4781</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2092.5,222,-2092.5</points>
<connection>
<GID>6672</GID>
<name>OUT</name></connection>
<connection>
<GID>6675</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6677</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6682</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6685</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6687</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6689</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6691</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-2161.5,40.5,-1996.5</points>
<connection>
<GID>6719</GID>
<name>N_in1</name></connection>
<connection>
<GID>6692</GID>
<name>N_in0</name></connection>
<intersection>-2136 12</intersection>
<intersection>-2117.5 11</intersection>
<intersection>-2098.5 10</intersection>
<intersection>-2080 9</intersection>
<intersection>-2058 8</intersection>
<intersection>-2039.5 7</intersection>
<intersection>-2020.5 6</intersection>
<intersection>-2002 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-2002,46,-2002</points>
<connection>
<GID>6508</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40.5,-2020.5,46,-2020.5</points>
<connection>
<GID>6835</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>40.5,-2039.5,46,-2039.5</points>
<connection>
<GID>6799</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>40.5,-2058,46,-2058</points>
<connection>
<GID>6721</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>40.5,-2080,46,-2080</points>
<connection>
<GID>6674</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>40.5,-2098.5,46,-2098.5</points>
<connection>
<GID>6550</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>40.5,-2117.5,46,-2117.5</points>
<connection>
<GID>6644</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>40.5,-2136,46,-2136</points>
<connection>
<GID>6544</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-2161,63.5,-1996</points>
<connection>
<GID>6723</GID>
<name>N_in1</name></connection>
<connection>
<GID>6693</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 4</intersection>
<intersection>-2126 5</intersection>
<intersection>-2107 6</intersection>
<intersection>-2088.5 7</intersection>
<intersection>-2066.5 8</intersection>
<intersection>-2048 9</intersection>
<intersection>-2029 10</intersection>
<intersection>-2010.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>59,-2144.5,63.5,-2144.5</points>
<intersection>59 12</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>59,-2126,63.5,-2126</points>
<intersection>59 14</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59,-2107,63.5,-2107</points>
<intersection>59 13</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59,-2088.5,63.5,-2088.5</points>
<intersection>59 15</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>59,-2066.5,63.5,-2066.5</points>
<intersection>59 18</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>59,-2048,63.5,-2048</points>
<intersection>59 19</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>59,-2029,63.5,-2029</points>
<intersection>59 20</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>59,-2010.5,63.5,-2010.5</points>
<intersection>59 21</intersection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>59,-2146,59,-2144.5</points>
<connection>
<GID>6547</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>59,-2108.5,59,-2107</points>
<connection>
<GID>6555</GID>
<name>OUT_0</name></connection>
<intersection>-2107 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>59,-2127.5,59,-2126</points>
<connection>
<GID>6645</GID>
<name>OUT_0</name></connection>
<intersection>-2126 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>59,-2090,59,-2088.5</points>
<connection>
<GID>6675</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>59,-2068,59,-2066.5</points>
<connection>
<GID>6733</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>59,-2049.5,59,-2048</points>
<connection>
<GID>6801</GID>
<name>OUT_0</name></connection>
<intersection>-2048 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>59,-2030.5,59,-2029</points>
<connection>
<GID>6837</GID>
<name>OUT_0</name></connection>
<intersection>-2029 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>59,-2012,59,-2010.5</points>
<connection>
<GID>6510</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>4784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-2161,66.5,-1996.5</points>
<connection>
<GID>6725</GID>
<name>N_in1</name></connection>
<connection>
<GID>6694</GID>
<name>N_in0</name></connection>
<intersection>-2136 10</intersection>
<intersection>-2117.5 9</intersection>
<intersection>-2098.5 8</intersection>
<intersection>-2080 7</intersection>
<intersection>-2058 6</intersection>
<intersection>-2039.5 5</intersection>
<intersection>-2020.5 4</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>66.5,-2002,69,-2002</points>
<connection>
<GID>6512</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-2020.5,69,-2020.5</points>
<connection>
<GID>6839</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66.5,-2039.5,69,-2039.5</points>
<connection>
<GID>6803</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66.5,-2058,69,-2058</points>
<connection>
<GID>6757</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66.5,-2080,69,-2080</points>
<connection>
<GID>6676</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-2098.5,69,-2098.5</points>
<connection>
<GID>6560</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66.5,-2117.5,69,-2117.5</points>
<connection>
<GID>6646</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>66.5,-2136,69,-2136</points>
<connection>
<GID>6549</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-2161,86,-1996</points>
<connection>
<GID>6727</GID>
<name>N_in1</name></connection>
<connection>
<GID>6695</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 6</intersection>
<intersection>-2126 7</intersection>
<intersection>-2107 8</intersection>
<intersection>-2088.5 9</intersection>
<intersection>-2066.5 10</intersection>
<intersection>-2048 11</intersection>
<intersection>-2029 12</intersection>
<intersection>-2010.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>82,-2144.5,86,-2144.5</points>
<intersection>82 14</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82,-2126,86,-2126</points>
<intersection>82 16</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>82,-2107,86,-2107</points>
<intersection>82 15</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82,-2088.5,86,-2088.5</points>
<intersection>82 17</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>82,-2066.5,86,-2066.5</points>
<intersection>82 20</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>82,-2048,86,-2048</points>
<intersection>82 21</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>82,-2029,86,-2029</points>
<intersection>82 22</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>82,-2010.5,86,-2010.5</points>
<intersection>82 23</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>82,-2146,82,-2144.5</points>
<connection>
<GID>6552</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>82,-2108.5,82,-2107</points>
<connection>
<GID>6565</GID>
<name>OUT_0</name></connection>
<intersection>-2107 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>82,-2127.5,82,-2126</points>
<connection>
<GID>6647</GID>
<name>OUT_0</name></connection>
<intersection>-2126 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>82,-2090,82,-2088.5</points>
<connection>
<GID>6677</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>82,-2068,82,-2066.5</points>
<connection>
<GID>6759</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>82,-2049.5,82,-2048</points>
<connection>
<GID>6805</GID>
<name>OUT_0</name></connection>
<intersection>-2048 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>82,-2030.5,82,-2029</points>
<connection>
<GID>6841</GID>
<name>OUT_0</name></connection>
<intersection>-2029 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>82,-2012,82,-2010.5</points>
<connection>
<GID>6514</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-2161,89.5,-1996</points>
<connection>
<GID>6729</GID>
<name>N_in1</name></connection>
<connection>
<GID>6696</GID>
<name>N_in0</name></connection>
<intersection>-2136 13</intersection>
<intersection>-2117.5 12</intersection>
<intersection>-2098.5 11</intersection>
<intersection>-2080 10</intersection>
<intersection>-2058 9</intersection>
<intersection>-2039.5 8</intersection>
<intersection>-2020.5 7</intersection>
<intersection>-2002 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-2002,94,-2002</points>
<connection>
<GID>6516</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-2020.5,94,-2020.5</points>
<connection>
<GID>6843</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89.5,-2039.5,94,-2039.5</points>
<connection>
<GID>6807</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-2058,94,-2058</points>
<connection>
<GID>6763</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>89.5,-2080,94,-2080</points>
<connection>
<GID>6679</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89.5,-2098.5,94,-2098.5</points>
<connection>
<GID>6570</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>89.5,-2117.5,94,-2117.5</points>
<connection>
<GID>6648</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>89.5,-2136,94,-2136</points>
<connection>
<GID>6554</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-2161,110.5,-1996.5</points>
<connection>
<GID>6731</GID>
<name>N_in1</name></connection>
<connection>
<GID>6697</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 6</intersection>
<intersection>-2126 7</intersection>
<intersection>-2107 8</intersection>
<intersection>-2088.5 9</intersection>
<intersection>-2066.5 10</intersection>
<intersection>-2048 11</intersection>
<intersection>-2029 12</intersection>
<intersection>-2010.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>107,-2144.5,110.5,-2144.5</points>
<intersection>107 14</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>107,-2126,110.5,-2126</points>
<intersection>107 16</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>107,-2107,110.5,-2107</points>
<intersection>107 15</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>107,-2088.5,110.5,-2088.5</points>
<intersection>107 17</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>107,-2066.5,110.5,-2066.5</points>
<intersection>107 20</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>107,-2048,110.5,-2048</points>
<intersection>107 21</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>107,-2029,110.5,-2029</points>
<intersection>107 22</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>107,-2010.5,110.5,-2010.5</points>
<intersection>107 23</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>107,-2146,107,-2144.5</points>
<connection>
<GID>6557</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>107,-2108.5,107,-2107</points>
<connection>
<GID>6574</GID>
<name>OUT_0</name></connection>
<intersection>-2107 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>107,-2127.5,107,-2126</points>
<connection>
<GID>6649</GID>
<name>OUT_0</name></connection>
<intersection>-2126 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>107,-2090,107,-2088.5</points>
<connection>
<GID>6680</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>107,-2068,107,-2066.5</points>
<connection>
<GID>6767</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>107,-2049.5,107,-2048</points>
<connection>
<GID>6809</GID>
<name>OUT_0</name></connection>
<intersection>-2048 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>107,-2030.5,107,-2029</points>
<connection>
<GID>6845</GID>
<name>OUT_0</name></connection>
<intersection>-2029 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>107,-2012,107,-2010.5</points>
<connection>
<GID>6518</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2161,114.5,-1996</points>
<connection>
<GID>6735</GID>
<name>N_in1</name></connection>
<connection>
<GID>6698</GID>
<name>N_in0</name></connection>
<intersection>-2136 13</intersection>
<intersection>-2117.5 12</intersection>
<intersection>-2098.5 11</intersection>
<intersection>-2080 10</intersection>
<intersection>-2058 9</intersection>
<intersection>-2039.5 8</intersection>
<intersection>-2020.5 7</intersection>
<intersection>-2002 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>114.5,-2002,117,-2002</points>
<connection>
<GID>6520</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-2020.5,117,-2020.5</points>
<connection>
<GID>6847</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-2039.5,117,-2039.5</points>
<connection>
<GID>6811</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114.5,-2058,117,-2058</points>
<connection>
<GID>6771</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114.5,-2080,117,-2080</points>
<connection>
<GID>6681</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>114.5,-2098.5,117,-2098.5</points>
<connection>
<GID>6577</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114.5,-2117.5,117,-2117.5</points>
<connection>
<GID>6650</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>114.5,-2136,117,-2136</points>
<connection>
<GID>6559</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4789</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-2161,133,-1996</points>
<connection>
<GID>6737</GID>
<name>N_in1</name></connection>
<connection>
<GID>6699</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 6</intersection>
<intersection>-2126 7</intersection>
<intersection>-2107 8</intersection>
<intersection>-2088.5 9</intersection>
<intersection>-2066.5 10</intersection>
<intersection>-2048 11</intersection>
<intersection>-2029 12</intersection>
<intersection>-2010.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>130,-2144.5,133,-2144.5</points>
<intersection>130 14</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-2126,133,-2126</points>
<intersection>130 15</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>130,-2107,133,-2107</points>
<intersection>130 16</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>130,-2088.5,133,-2088.5</points>
<intersection>130 17</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>130,-2066.5,133,-2066.5</points>
<intersection>130 20</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>130,-2048,133,-2048</points>
<intersection>130 21</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>130,-2029,133,-2029</points>
<intersection>130 22</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>130,-2010.5,133,-2010.5</points>
<intersection>130 23</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>130,-2146,130,-2144.5</points>
<connection>
<GID>6562</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>130,-2127.5,130,-2126</points>
<connection>
<GID>6651</GID>
<name>OUT_0</name></connection>
<intersection>-2126 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>130,-2108.5,130,-2107</points>
<connection>
<GID>6661</GID>
<name>OUT_0</name></connection>
<intersection>-2107 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>130,-2090,130,-2088.5</points>
<connection>
<GID>6682</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>130,-2068,130,-2066.5</points>
<connection>
<GID>6775</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>130,-2049.5,130,-2048</points>
<connection>
<GID>6813</GID>
<name>OUT_0</name></connection>
<intersection>-2048 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>130,-2030.5,130,-2029</points>
<connection>
<GID>6849</GID>
<name>OUT_0</name></connection>
<intersection>-2029 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>130,-2012,130,-2010.5</points>
<connection>
<GID>6522</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2161,137,-1996</points>
<connection>
<GID>6739</GID>
<name>N_in1</name></connection>
<connection>
<GID>6701</GID>
<name>N_in0</name></connection>
<intersection>-2136 13</intersection>
<intersection>-2117.5 12</intersection>
<intersection>-2098.5 11</intersection>
<intersection>-2080 10</intersection>
<intersection>-2058 9</intersection>
<intersection>-2039.5 8</intersection>
<intersection>-2020.5 7</intersection>
<intersection>-2002 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>137,-2002,140,-2002</points>
<connection>
<GID>6524</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137,-2020.5,140,-2020.5</points>
<connection>
<GID>6851</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-2039.5,140,-2039.5</points>
<connection>
<GID>6815</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137,-2058,140,-2058</points>
<connection>
<GID>6777</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-2080,140,-2080</points>
<connection>
<GID>6683</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>137,-2098.5,140,-2098.5</points>
<connection>
<GID>6662</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137,-2117.5,140,-2117.5</points>
<connection>
<GID>6652</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-2136,140,-2136</points>
<connection>
<GID>6564</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>4791</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-2160.5,156,-1996</points>
<connection>
<GID>6741</GID>
<name>N_in1</name></connection>
<connection>
<GID>6703</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 6</intersection>
<intersection>-2126 7</intersection>
<intersection>-2107 8</intersection>
<intersection>-2088.5 9</intersection>
<intersection>-2066.5 10</intersection>
<intersection>-2048 11</intersection>
<intersection>-2029 12</intersection>
<intersection>-2010.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>153,-2144.5,156,-2144.5</points>
<intersection>153 15</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>153,-2126,156,-2126</points>
<intersection>153 16</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>153,-2107,156,-2107</points>
<intersection>153 17</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>153,-2088.5,156,-2088.5</points>
<intersection>153 18</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>153,-2066.5,156,-2066.5</points>
<intersection>153 21</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>153,-2048,156,-2048</points>
<intersection>153 22</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>153,-2029,156,-2029</points>
<intersection>153 23</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>153,-2010.5,156,-2010.5</points>
<intersection>153 14</intersection>
<intersection>156 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>153,-2012,153,-2010.5</points>
<connection>
<GID>6526</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>153,-2146,153,-2144.5</points>
<connection>
<GID>6567</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>153,-2127.5,153,-2126</points>
<connection>
<GID>6653</GID>
<name>OUT_0</name></connection>
<intersection>-2126 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>153,-2108.5,153,-2107</points>
<connection>
<GID>6663</GID>
<name>OUT_0</name></connection>
<intersection>-2107 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>153,-2090,153,-2088.5</points>
<connection>
<GID>6685</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>153,-2068,153,-2066.5</points>
<connection>
<GID>6781</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>153,-2049.5,153,-2048</points>
<connection>
<GID>6817</GID>
<name>OUT_0</name></connection>
<intersection>-2048 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>153,-2030.5,153,-2029</points>
<connection>
<GID>6490</GID>
<name>OUT_0</name></connection>
<intersection>-2029 12</intersection></vsegment></shape></wire>
<wire>
<ID>4792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-2160.5,161,-1996</points>
<connection>
<GID>6743</GID>
<name>N_in1</name></connection>
<connection>
<GID>6705</GID>
<name>N_in0</name></connection>
<intersection>-2136 13</intersection>
<intersection>-2117.5 12</intersection>
<intersection>-2098.5 11</intersection>
<intersection>-2080 10</intersection>
<intersection>-2058 9</intersection>
<intersection>-2039.5 8</intersection>
<intersection>-2020.5 7</intersection>
<intersection>-2002 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>161,-2002,163,-2002</points>
<connection>
<GID>6528</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>161,-2020.5,163,-2020.5</points>
<connection>
<GID>6492</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>161,-2039.5,163,-2039.5</points>
<connection>
<GID>6819</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>161,-2058,163,-2058</points>
<connection>
<GID>6783</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>161,-2080,163,-2080</points>
<connection>
<GID>6686</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>161,-2098.5,163,-2098.5</points>
<connection>
<GID>6664</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>161,-2117.5,163,-2117.5</points>
<connection>
<GID>6654</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>161,-2136,163,-2136</points>
<connection>
<GID>6569</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>4793</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-2160,179,-1996</points>
<connection>
<GID>6745</GID>
<name>N_in1</name></connection>
<connection>
<GID>6709</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 16</intersection>
<intersection>-2126 15</intersection>
<intersection>-2107 14</intersection>
<intersection>-2088.5 13</intersection>
<intersection>-2066.5 12</intersection>
<intersection>-2048 11</intersection>
<intersection>-2029 10</intersection>
<intersection>-2010.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>176,-2010.5,179,-2010.5</points>
<intersection>176 17</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>176,-2029,179,-2029</points>
<intersection>176 26</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>176,-2048,179,-2048</points>
<intersection>176 25</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>176,-2066.5,179,-2066.5</points>
<intersection>176 24</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>176,-2088.5,179,-2088.5</points>
<intersection>176 21</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>176,-2107,179,-2107</points>
<intersection>176 20</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>176,-2126,179,-2126</points>
<intersection>176 19</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>176,-2144.5,179,-2144.5</points>
<intersection>176 18</intersection>
<intersection>179 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>176,-2012,176,-2010.5</points>
<connection>
<GID>6530</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>176,-2146,176,-2144.5</points>
<connection>
<GID>6572</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>176,-2127.5,176,-2126</points>
<connection>
<GID>6655</GID>
<name>OUT_0</name></connection>
<intersection>-2126 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>176,-2108.5,176,-2107</points>
<connection>
<GID>6665</GID>
<name>OUT_0</name></connection>
<intersection>-2107 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>176,-2090,176,-2088.5</points>
<connection>
<GID>6687</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>176,-2068,176,-2066.5</points>
<connection>
<GID>6785</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>176,-2049.5,176,-2048</points>
<connection>
<GID>6821</GID>
<name>OUT_0</name></connection>
<intersection>-2048 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>176,-2030.5,176,-2029</points>
<connection>
<GID>6494</GID>
<name>OUT_0</name></connection>
<intersection>-2029 10</intersection></vsegment></shape></wire>
<wire>
<ID>4794</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2160,183.5,-1996</points>
<connection>
<GID>6747</GID>
<name>N_in1</name></connection>
<connection>
<GID>6707</GID>
<name>N_in0</name></connection>
<intersection>-2136 13</intersection>
<intersection>-2117.5 12</intersection>
<intersection>-2098.5 11</intersection>
<intersection>-2080 10</intersection>
<intersection>-2058 9</intersection>
<intersection>-2039.5 8</intersection>
<intersection>-2020.5 7</intersection>
<intersection>-2002 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>183.5,-2002,188,-2002</points>
<connection>
<GID>6532</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>183.5,-2020.5,188,-2020.5</points>
<connection>
<GID>6496</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>183.5,-2039.5,188,-2039.5</points>
<connection>
<GID>6823</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>183.5,-2058,188,-2058</points>
<connection>
<GID>6787</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183.5,-2080,188,-2080</points>
<connection>
<GID>6688</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183.5,-2098.5,188,-2098.5</points>
<connection>
<GID>6666</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183.5,-2117.5,188,-2117.5</points>
<connection>
<GID>6656</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183.5,-2136,188,-2136</points>
<connection>
<GID>6638</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-2159.5,204.5,-1996.5</points>
<connection>
<GID>6749</GID>
<name>N_in1</name></connection>
<connection>
<GID>6711</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 6</intersection>
<intersection>-2126 7</intersection>
<intersection>-2107 8</intersection>
<intersection>-2088.5 9</intersection>
<intersection>-2066.5 10</intersection>
<intersection>-2048 11</intersection>
<intersection>-2029 12</intersection>
<intersection>-2010.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>201,-2144.5,204.5,-2144.5</points>
<intersection>201 15</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>201,-2126,204.5,-2126</points>
<intersection>201 16</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>201,-2107,204.5,-2107</points>
<intersection>201 17</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>201,-2088.5,204.5,-2088.5</points>
<intersection>201 18</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>201,-2066.5,204.5,-2066.5</points>
<intersection>201 21</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>201,-2048,204.5,-2048</points>
<intersection>201 22</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>201,-2029,204.5,-2029</points>
<intersection>201 23</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>201,-2010.5,204.5,-2010.5</points>
<intersection>201 14</intersection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>201,-2012,201,-2010.5</points>
<connection>
<GID>6534</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201,-2146,201,-2144.5</points>
<connection>
<GID>6639</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>201,-2127.5,201,-2126</points>
<connection>
<GID>6657</GID>
<name>OUT_0</name></connection>
<intersection>-2126 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>201,-2108.5,201,-2107</points>
<connection>
<GID>6667</GID>
<name>OUT_0</name></connection>
<intersection>-2107 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>201,-2090,201,-2088.5</points>
<connection>
<GID>6689</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>201,-2068,201,-2066.5</points>
<connection>
<GID>6789</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>201,-2049.5,201,-2048</points>
<connection>
<GID>6825</GID>
<name>OUT_0</name></connection>
<intersection>-2048 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>201,-2030.5,201,-2029</points>
<connection>
<GID>6498</GID>
<name>OUT_0</name></connection>
<intersection>-2029 12</intersection></vsegment></shape></wire>
<wire>
<ID>4796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-2159.5,208,-1996.5</points>
<connection>
<GID>6753</GID>
<name>N_in0</name></connection>
<connection>
<GID>6751</GID>
<name>N_in1</name></connection>
<intersection>-2136 11</intersection>
<intersection>-2117.5 10</intersection>
<intersection>-2098.5 9</intersection>
<intersection>-2080 7</intersection>
<intersection>-2058 6</intersection>
<intersection>-2039.5 5</intersection>
<intersection>-2020.5 4</intersection>
<intersection>-2002 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208,-2002,211,-2002</points>
<connection>
<GID>6536</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208,-2020.5,211,-2020.5</points>
<connection>
<GID>6500</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>208,-2039.5,211,-2039.5</points>
<connection>
<GID>6827</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>208,-2058,211,-2058</points>
<connection>
<GID>6791</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>208,-2080,211,-2080</points>
<connection>
<GID>6690</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>208,-2098.5,211,-2098.5</points>
<connection>
<GID>6669</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>208,-2117.5,211,-2117.5</points>
<connection>
<GID>6658</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>208,-2136,211,-2136</points>
<connection>
<GID>6640</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>4797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-2159.5,229,-1997.5</points>
<connection>
<GID>6755</GID>
<name>N_in1</name></connection>
<connection>
<GID>6713</GID>
<name>N_in0</name></connection>
<intersection>-2144.5 11</intersection>
<intersection>-2126 10</intersection>
<intersection>-2107 9</intersection>
<intersection>-2088.5 8</intersection>
<intersection>-2066.5 7</intersection>
<intersection>-2048 6</intersection>
<intersection>-2029 5</intersection>
<intersection>-2010.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>224,-2010.5,229,-2010.5</points>
<intersection>224 12</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>224,-2029,229,-2029</points>
<intersection>224 21</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>224,-2048,229,-2048</points>
<intersection>224 20</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>224,-2066.5,229,-2066.5</points>
<intersection>224 19</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>224,-2088.5,229,-2088.5</points>
<intersection>224 16</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>224,-2107,229,-2107</points>
<intersection>224 15</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>224,-2126,229,-2126</points>
<intersection>224 14</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>224,-2144.5,229,-2144.5</points>
<intersection>224 13</intersection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>224,-2012,224,-2010.5</points>
<connection>
<GID>6538</GID>
<name>OUT_0</name></connection>
<intersection>-2010.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>224,-2146,224,-2144.5</points>
<connection>
<GID>6641</GID>
<name>OUT_0</name></connection>
<intersection>-2144.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>224,-2127.5,224,-2126</points>
<connection>
<GID>6659</GID>
<name>OUT_0</name></connection>
<intersection>-2126 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>224,-2108.5,224,-2107</points>
<connection>
<GID>6670</GID>
<name>OUT_0</name></connection>
<intersection>-2107 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>224,-2090,224,-2088.5</points>
<connection>
<GID>6691</GID>
<name>OUT_0</name></connection>
<intersection>-2088.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>224,-2068,224,-2066.5</points>
<connection>
<GID>6793</GID>
<name>OUT_0</name></connection>
<intersection>-2066.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>224,-2049.5,224,-2048</points>
<connection>
<GID>6829</GID>
<name>OUT_0</name></connection>
<intersection>-2048 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>224,-2030.5,224,-2029</points>
<connection>
<GID>6502</GID>
<name>OUT_0</name></connection>
<intersection>-2029 5</intersection></vsegment></shape></wire>
<wire>
<ID>4798</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-121,-2004,18.5,-2004</points>
<connection>
<GID>6504</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-2013.5,-121,-1988</points>
<intersection>-2013.5 4</intersection>
<intersection>-2004 2</intersection>
<intersection>-1988 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-2013.5,30,-2013.5</points>
<connection>
<GID>6506</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-1988,-121,-1988</points>
<connection>
<GID>6637</GID>
<name>OUT_7</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4799</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-122,-2022.5,18.5,-2022.5</points>
<connection>
<GID>6831</GID>
<name>IN_0</name></connection>
<intersection>-122 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-122,-2032,-122,-1989</points>
<intersection>-2032 5</intersection>
<intersection>-2022.5 2</intersection>
<intersection>-1989 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-122,-2032,30,-2032</points>
<connection>
<GID>6833</GID>
<name>IN_0</name></connection>
<intersection>-122 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-1989,-122,-1989</points>
<connection>
<GID>6637</GID>
<name>OUT_6</name></connection>
<intersection>-122 4</intersection></hsegment></shape></wire>
<wire>
<ID>4800</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-123,-2041.5,18.5,-2041.5</points>
<connection>
<GID>6795</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-2051,-123,-1990</points>
<intersection>-2051 4</intersection>
<intersection>-2041.5 2</intersection>
<intersection>-1990 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-2051,30,-2051</points>
<connection>
<GID>6797</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-1990,-123,-1990</points>
<connection>
<GID>6637</GID>
<name>OUT_5</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>4801</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-124,-2060,18.5,-2060</points>
<connection>
<GID>6715</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-2069.5,-124,-1991</points>
<intersection>-2069.5 4</intersection>
<intersection>-2060 2</intersection>
<intersection>-1991 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-2069.5,30,-2069.5</points>
<connection>
<GID>6717</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1991,-124,-1991</points>
<connection>
<GID>6637</GID>
<name>OUT_4</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>4802</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125,-2082,18.5,-2082</points>
<connection>
<GID>6671</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-125,-2091.5,-125,-1992</points>
<intersection>-2091.5 4</intersection>
<intersection>-2082 1</intersection>
<intersection>-1992 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-125,-2091.5,29.5,-2091.5</points>
<connection>
<GID>6672</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1992,-125,-1992</points>
<connection>
<GID>6637</GID>
<name>OUT_3</name></connection>
<intersection>-125 3</intersection></hsegment></shape></wire>
<wire>
<ID>4803</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,-2100.5,18.5,-2100.5</points>
<connection>
<GID>6660</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-2110,-126,-1993</points>
<intersection>-2110 4</intersection>
<intersection>-2100.5 1</intersection>
<intersection>-1993 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-2110,29.5,-2110</points>
<connection>
<GID>6545</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1993,-126,-1993</points>
<connection>
<GID>6637</GID>
<name>OUT_2</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>4804</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127,-2119.5,18.5,-2119.5</points>
<connection>
<GID>6642</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-127,-2129,-127,-1994</points>
<intersection>-2129 4</intersection>
<intersection>-2119.5 1</intersection>
<intersection>-1994 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-127,-2129,29.5,-2129</points>
<connection>
<GID>6643</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1994,-127,-1994</points>
<connection>
<GID>6637</GID>
<name>OUT_1</name></connection>
<intersection>-127 3</intersection></hsegment></shape></wire>
<wire>
<ID>4805</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-128,-2138,18.5,-2138</points>
<connection>
<GID>6540</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-2147.5,-128,-1995</points>
<connection>
<GID>6637</GID>
<name>OUT_0</name></connection>
<intersection>-2147.5 4</intersection>
<intersection>-2138 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-2147.5,29.5,-2147.5</points>
<connection>
<GID>6542</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>4806</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-2161.5,17.5,-1996.5</points>
<connection>
<GID>6773</GID>
<name>N_in1</name></connection>
<connection>
<GID>6765</GID>
<name>N_in0</name></connection>
<intersection>-2140 10</intersection>
<intersection>-2121.5 9</intersection>
<intersection>-2102.5 8</intersection>
<intersection>-2084 7</intersection>
<intersection>-2062 6</intersection>
<intersection>-2043.5 5</intersection>
<intersection>-2024.5 4</intersection>
<intersection>-2006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-2006,18.5,-2006</points>
<connection>
<GID>6504</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-2024.5,18.5,-2024.5</points>
<connection>
<GID>6831</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>17.5,-2043.5,18.5,-2043.5</points>
<connection>
<GID>6795</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>17.5,-2062,18.5,-2062</points>
<connection>
<GID>6715</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>17.5,-2084,18.5,-2084</points>
<connection>
<GID>6671</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>17.5,-2102.5,18.5,-2102.5</points>
<connection>
<GID>6660</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>17.5,-2121.5,18.5,-2121.5</points>
<connection>
<GID>6642</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>17.5,-2140,18.5,-2140</points>
<connection>
<GID>6540</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-2161.5,27.5,-1996.5</points>
<connection>
<GID>6769</GID>
<name>N_in1</name></connection>
<connection>
<GID>6761</GID>
<name>N_in0</name></connection>
<intersection>-2149.5 3</intersection>
<intersection>-2131 5</intersection>
<intersection>-2112 7</intersection>
<intersection>-2093.5 9</intersection>
<intersection>-2071.5 11</intersection>
<intersection>-2053 13</intersection>
<intersection>-2034 15</intersection>
<intersection>-2015.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-2149.5,29.5,-2149.5</points>
<connection>
<GID>6542</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-2131,29.5,-2131</points>
<connection>
<GID>6643</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-2112,29.5,-2112</points>
<connection>
<GID>6545</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>27.5,-2093.5,29.5,-2093.5</points>
<connection>
<GID>6672</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>27.5,-2071.5,30,-2071.5</points>
<connection>
<GID>6717</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>27.5,-2053,30,-2053</points>
<connection>
<GID>6797</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>27.5,-2034,30,-2034</points>
<connection>
<GID>6833</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>27.5,-2015.5,30,-2015.5</points>
<connection>
<GID>6506</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-1994.5,17.5,-1988</points>
<connection>
<GID>6765</GID>
<name>N_in1</name></connection>
<connection>
<GID>6635</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-1994.5,27.5,-1988</points>
<connection>
<GID>6761</GID>
<name>N_in1</name></connection>
<connection>
<GID>6634</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4810</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-1994.5,40.5,-1988</points>
<connection>
<GID>6692</GID>
<name>N_in1</name></connection>
<connection>
<GID>6615</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-1994,63.5,-1987.5</points>
<connection>
<GID>6693</GID>
<name>N_in1</name></connection>
<connection>
<GID>6616</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-1994.5,66.5,-1987.5</points>
<connection>
<GID>6694</GID>
<name>N_in1</name></connection>
<connection>
<GID>6617</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4813</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-1994,86,-1987.5</points>
<connection>
<GID>6695</GID>
<name>N_in1</name></connection>
<connection>
<GID>6618</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-1994,89.5,-1987.5</points>
<connection>
<GID>6696</GID>
<name>N_in1</name></connection>
<connection>
<GID>6619</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-1994.5,110.5,-1987.5</points>
<connection>
<GID>6697</GID>
<name>N_in1</name></connection>
<connection>
<GID>6620</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4816</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-1994,114.5,-1987.5</points>
<connection>
<GID>6698</GID>
<name>N_in1</name></connection>
<connection>
<GID>6621</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4817</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1994,133,-1987.5</points>
<connection>
<GID>6699</GID>
<name>N_in1</name></connection>
<connection>
<GID>6622</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-1994,137,-1987.5</points>
<connection>
<GID>6701</GID>
<name>N_in1</name></connection>
<connection>
<GID>6623</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4819</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-1994,156,-1987</points>
<connection>
<GID>6703</GID>
<name>N_in1</name></connection>
<connection>
<GID>6624</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-1994,161,-1987</points>
<connection>
<GID>6705</GID>
<name>N_in1</name></connection>
<connection>
<GID>6625</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4821</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-1994,179,-1986.5</points>
<connection>
<GID>6709</GID>
<name>N_in1</name></connection>
<connection>
<GID>6626</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-1994,183.5,-1986.5</points>
<connection>
<GID>6707</GID>
<name>N_in1</name></connection>
<connection>
<GID>6627</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4823</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-1994.5,204.5,-1986</points>
<connection>
<GID>6711</GID>
<name>N_in1</name></connection>
<connection>
<GID>6628</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-1994.5,208,-1986</points>
<connection>
<GID>6753</GID>
<name>N_in1</name></connection>
<connection>
<GID>6629</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4825</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-1995.5,229,-1986</points>
<connection>
<GID>6713</GID>
<name>N_in1</name></connection>
<connection>
<GID>6631</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2258,59,-2258</points>
<connection>
<GID>7049</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2258,53,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2242.5,53,-2242.5</points>
<connection>
<GID>7043</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4827</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2258,82,-2258</points>
<connection>
<GID>7067</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2258,76,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2242.5,76,-2242.5</points>
<connection>
<GID>7065</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4828</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2258,107,-2258</points>
<connection>
<GID>7071</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2258,101,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2242.5,101,-2242.5</points>
<connection>
<GID>7069</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4829</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2258,130,-2258</points>
<connection>
<GID>7075</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2258,124,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2242.5,124,-2242.5</points>
<connection>
<GID>7073</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4830</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2258,153,-2258</points>
<connection>
<GID>7079</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2258,147,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2242.5,147,-2242.5</points>
<connection>
<GID>7077</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4831</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2258,176,-2258</points>
<connection>
<GID>7083</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2258,170,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2242.5,170,-2242.5</points>
<connection>
<GID>7081</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4832</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2258,201,-2258</points>
<connection>
<GID>7087</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2258,195,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2242.5,195,-2242.5</points>
<connection>
<GID>7085</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4833</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2258,224,-2258</points>
<connection>
<GID>7091</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2258,218,-2242.5</points>
<intersection>-2258 1</intersection>
<intersection>-2242.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2242.5,218,-2242.5</points>
<connection>
<GID>7089</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4834</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2245.5,211,-2245.5</points>
<connection>
<GID>7033</GID>
<name>OUT</name></connection>
<connection>
<GID>7043</GID>
<name>clock</name></connection>
<connection>
<GID>7065</GID>
<name>clock</name></connection>
<connection>
<GID>7069</GID>
<name>clock</name></connection>
<connection>
<GID>7073</GID>
<name>clock</name></connection>
<connection>
<GID>7077</GID>
<name>clock</name></connection>
<connection>
<GID>7081</GID>
<name>clock</name></connection>
<connection>
<GID>7085</GID>
<name>clock</name></connection>
<connection>
<GID>7089</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4835</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2255,222,-2255</points>
<connection>
<GID>7038</GID>
<name>OUT</name></connection>
<connection>
<GID>7049</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7067</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7071</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7075</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7079</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7083</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7087</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7091</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4836</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2239.5,59,-2239.5</points>
<connection>
<GID>7099</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2239.5,53,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2224,53,-2224</points>
<connection>
<GID>7097</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4837</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2239.5,82,-2239.5</points>
<connection>
<GID>7103</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2239.5,76,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2224,76,-2224</points>
<connection>
<GID>7101</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4838</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2239.5,107,-2239.5</points>
<connection>
<GID>7107</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2239.5,101,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2224,101,-2224</points>
<connection>
<GID>7105</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4839</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2239.5,130,-2239.5</points>
<connection>
<GID>7111</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2239.5,124,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2224,124,-2224</points>
<connection>
<GID>7109</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4840</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2239.5,153,-2239.5</points>
<connection>
<GID>7115</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2239.5,147,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2224,147,-2224</points>
<connection>
<GID>7113</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4841</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2239.5,176,-2239.5</points>
<connection>
<GID>7119</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2239.5,170,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2224,170,-2224</points>
<connection>
<GID>7117</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4842</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2239.5,201,-2239.5</points>
<connection>
<GID>7123</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2239.5,195,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2224,195,-2224</points>
<connection>
<GID>7121</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4843</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2239.5,224,-2239.5</points>
<connection>
<GID>7127</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2239.5,218,-2224</points>
<intersection>-2239.5 1</intersection>
<intersection>-2224 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2224,218,-2224</points>
<connection>
<GID>7125</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4844</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2227,211,-2227</points>
<connection>
<GID>7093</GID>
<name>OUT</name></connection>
<connection>
<GID>7097</GID>
<name>clock</name></connection>
<connection>
<GID>7101</GID>
<name>clock</name></connection>
<connection>
<GID>7105</GID>
<name>clock</name></connection>
<connection>
<GID>7109</GID>
<name>clock</name></connection>
<connection>
<GID>7113</GID>
<name>clock</name></connection>
<connection>
<GID>7117</GID>
<name>clock</name></connection>
<connection>
<GID>7121</GID>
<name>clock</name></connection>
<connection>
<GID>7125</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4845</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2236.5,222,-2236.5</points>
<connection>
<GID>7095</GID>
<name>OUT</name></connection>
<connection>
<GID>7099</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7103</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7107</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7111</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7115</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7119</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7123</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7127</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4846</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2220.5,59,-2220.5</points>
<connection>
<GID>7135</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2220.5,53,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2205,53,-2205</points>
<connection>
<GID>7133</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4847</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2220.5,82,-2220.5</points>
<connection>
<GID>7139</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2220.5,76,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2205,76,-2205</points>
<connection>
<GID>7137</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4848</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2220.5,107,-2220.5</points>
<connection>
<GID>7143</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2220.5,101,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2205,101,-2205</points>
<connection>
<GID>7141</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4849</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2220.5,130,-2220.5</points>
<connection>
<GID>7147</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2220.5,124,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2205,124,-2205</points>
<connection>
<GID>7145</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4850</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2220.5,153,-2220.5</points>
<connection>
<GID>7151</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2220.5,147,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2205,147,-2205</points>
<connection>
<GID>7149</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4851</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2220.5,176,-2220.5</points>
<connection>
<GID>7155</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2220.5,170,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2205,170,-2205</points>
<connection>
<GID>7153</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4852</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2220.5,201,-2220.5</points>
<connection>
<GID>7159</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2220.5,195,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2205,195,-2205</points>
<connection>
<GID>7157</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4853</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2220.5,224,-2220.5</points>
<connection>
<GID>7163</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2220.5,218,-2205</points>
<intersection>-2220.5 1</intersection>
<intersection>-2205 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2205,218,-2205</points>
<connection>
<GID>7161</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4854</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2208,211,-2208</points>
<connection>
<GID>7129</GID>
<name>OUT</name></connection>
<connection>
<GID>7133</GID>
<name>clock</name></connection>
<connection>
<GID>7137</GID>
<name>clock</name></connection>
<connection>
<GID>7141</GID>
<name>clock</name></connection>
<connection>
<GID>7145</GID>
<name>clock</name></connection>
<connection>
<GID>7149</GID>
<name>clock</name></connection>
<connection>
<GID>7153</GID>
<name>clock</name></connection>
<connection>
<GID>7157</GID>
<name>clock</name></connection>
<connection>
<GID>7161</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4855</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2217.5,222,-2217.5</points>
<connection>
<GID>7131</GID>
<name>OUT</name></connection>
<connection>
<GID>7135</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7139</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7143</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7147</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7151</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7155</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7159</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7163</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4856</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2202,59,-2202</points>
<connection>
<GID>7171</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2202,53,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2186.5,53,-2186.5</points>
<connection>
<GID>7169</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4857</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2202,82,-2202</points>
<connection>
<GID>7175</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2202,76,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2186.5,76,-2186.5</points>
<connection>
<GID>7173</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4858</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2202,107,-2202</points>
<connection>
<GID>7179</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2202,101,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2186.5,101,-2186.5</points>
<connection>
<GID>7177</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4859</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2202,130,-2202</points>
<connection>
<GID>7183</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2202,124,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2186.5,124,-2186.5</points>
<connection>
<GID>7181</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4860</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2202,153,-2202</points>
<connection>
<GID>7187</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2202,147,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2186.5,147,-2186.5</points>
<connection>
<GID>7185</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4861</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2202,176,-2202</points>
<connection>
<GID>7191</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2202,170,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2186.5,170,-2186.5</points>
<connection>
<GID>7189</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4862</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2202,201,-2202</points>
<connection>
<GID>7195</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2202,195,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2186.5,195,-2186.5</points>
<connection>
<GID>7193</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4863</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2202,224,-2202</points>
<connection>
<GID>7199</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2202,218,-2186.5</points>
<intersection>-2202 1</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2186.5,218,-2186.5</points>
<connection>
<GID>7197</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4864</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2189.5,211,-2189.5</points>
<connection>
<GID>7165</GID>
<name>OUT</name></connection>
<connection>
<GID>7169</GID>
<name>clock</name></connection>
<connection>
<GID>7173</GID>
<name>clock</name></connection>
<connection>
<GID>7177</GID>
<name>clock</name></connection>
<connection>
<GID>7181</GID>
<name>clock</name></connection>
<connection>
<GID>7185</GID>
<name>clock</name></connection>
<connection>
<GID>7189</GID>
<name>clock</name></connection>
<connection>
<GID>7193</GID>
<name>clock</name></connection>
<connection>
<GID>7197</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4865</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2199,222,-2199</points>
<connection>
<GID>7167</GID>
<name>OUT</name></connection>
<connection>
<GID>7171</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7175</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7179</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7183</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7187</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7191</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7195</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7199</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4866</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2336,59,-2336</points>
<connection>
<GID>7207</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2336,53,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2320.5,53,-2320.5</points>
<connection>
<GID>7205</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4867</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2336,82,-2336</points>
<connection>
<GID>7211</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2336,76,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2320.5,76,-2320.5</points>
<connection>
<GID>7209</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4868</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2336,107,-2336</points>
<connection>
<GID>7215</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2336,101,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2320.5,101,-2320.5</points>
<connection>
<GID>7213</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4869</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2336,130,-2336</points>
<connection>
<GID>6856</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2336,124,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2320.5,124,-2320.5</points>
<connection>
<GID>6854</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4870</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2336,153,-2336</points>
<connection>
<GID>6860</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2336,147,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2320.5,147,-2320.5</points>
<connection>
<GID>6858</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4871</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2336,176,-2336</points>
<connection>
<GID>6864</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2336,170,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2320.5,170,-2320.5</points>
<connection>
<GID>6862</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4872</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2336,201,-2336</points>
<connection>
<GID>6868</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2336,195,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2320.5,195,-2320.5</points>
<connection>
<GID>6866</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4873</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2336,224,-2336</points>
<connection>
<GID>6872</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2336,218,-2320.5</points>
<intersection>-2336 1</intersection>
<intersection>-2320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2320.5,218,-2320.5</points>
<connection>
<GID>6870</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4874</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2323.5,211,-2323.5</points>
<connection>
<GID>7213</GID>
<name>clock</name></connection>
<connection>
<GID>7209</GID>
<name>clock</name></connection>
<connection>
<GID>7205</GID>
<name>clock</name></connection>
<connection>
<GID>7201</GID>
<name>OUT</name></connection>
<connection>
<GID>6870</GID>
<name>clock</name></connection>
<connection>
<GID>6866</GID>
<name>clock</name></connection>
<connection>
<GID>6862</GID>
<name>clock</name></connection>
<connection>
<GID>6858</GID>
<name>clock</name></connection>
<connection>
<GID>6854</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4875</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2333,222,-2333</points>
<connection>
<GID>7215</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7211</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7207</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7203</GID>
<name>OUT</name></connection>
<connection>
<GID>6872</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6868</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6864</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6860</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6856</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4876</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2317.5,59,-2317.5</points>
<connection>
<GID>6880</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2317.5,53,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2302,53,-2302</points>
<connection>
<GID>6878</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4877</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2317.5,82,-2317.5</points>
<connection>
<GID>6884</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2317.5,76,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2302,76,-2302</points>
<connection>
<GID>6882</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4878</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2317.5,107,-2317.5</points>
<connection>
<GID>6888</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2317.5,101,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2302,101,-2302</points>
<connection>
<GID>6886</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4879</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2317.5,130,-2317.5</points>
<connection>
<GID>6892</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2317.5,124,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2302,124,-2302</points>
<connection>
<GID>6890</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4880</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2317.5,153,-2317.5</points>
<connection>
<GID>6896</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2317.5,147,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2302,147,-2302</points>
<connection>
<GID>6894</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4881</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2317.5,176,-2317.5</points>
<connection>
<GID>6900</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2317.5,170,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2302,170,-2302</points>
<connection>
<GID>6898</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4882</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2317.5,201,-2317.5</points>
<connection>
<GID>6904</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2317.5,195,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2302,195,-2302</points>
<connection>
<GID>6902</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4883</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2317.5,224,-2317.5</points>
<connection>
<GID>6908</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2317.5,218,-2302</points>
<intersection>-2317.5 1</intersection>
<intersection>-2302 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2302,218,-2302</points>
<connection>
<GID>6906</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4884</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2305,211,-2305</points>
<connection>
<GID>6874</GID>
<name>OUT</name></connection>
<connection>
<GID>6878</GID>
<name>clock</name></connection>
<connection>
<GID>6882</GID>
<name>clock</name></connection>
<connection>
<GID>6886</GID>
<name>clock</name></connection>
<connection>
<GID>6890</GID>
<name>clock</name></connection>
<connection>
<GID>6894</GID>
<name>clock</name></connection>
<connection>
<GID>6898</GID>
<name>clock</name></connection>
<connection>
<GID>6902</GID>
<name>clock</name></connection>
<connection>
<GID>6906</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4885</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2314.5,222,-2314.5</points>
<connection>
<GID>6876</GID>
<name>OUT</name></connection>
<connection>
<GID>6880</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6884</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6888</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6892</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6896</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6900</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6904</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6908</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4886</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2298.5,59,-2298.5</points>
<connection>
<GID>6918</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2298.5,53,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2283,53,-2283</points>
<connection>
<GID>6916</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4887</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2298.5,82,-2298.5</points>
<connection>
<GID>6923</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2298.5,76,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2283,76,-2283</points>
<connection>
<GID>6921</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4888</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2298.5,107,-2298.5</points>
<connection>
<GID>6928</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2298.5,101,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2283,101,-2283</points>
<connection>
<GID>6926</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4889</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2298.5,130,-2298.5</points>
<connection>
<GID>6933</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2298.5,124,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2283,124,-2283</points>
<connection>
<GID>6931</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4890</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2298.5,153,-2298.5</points>
<connection>
<GID>6938</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2298.5,147,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2283,147,-2283</points>
<connection>
<GID>6936</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4891</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2298.5,176,-2298.5</points>
<connection>
<GID>6941</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2298.5,170,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2283,170,-2283</points>
<connection>
<GID>6940</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4892</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2298.5,201,-2298.5</points>
<connection>
<GID>6944</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2298.5,195,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2283,195,-2283</points>
<connection>
<GID>6943</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4893</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2298.5,224,-2298.5</points>
<connection>
<GID>6946</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2298.5,218,-2283</points>
<intersection>-2298.5 1</intersection>
<intersection>-2283 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2283,218,-2283</points>
<connection>
<GID>6945</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4894</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2286,211,-2286</points>
<connection>
<GID>6911</GID>
<name>OUT</name></connection>
<connection>
<GID>6916</GID>
<name>clock</name></connection>
<connection>
<GID>6921</GID>
<name>clock</name></connection>
<connection>
<GID>6926</GID>
<name>clock</name></connection>
<connection>
<GID>6931</GID>
<name>clock</name></connection>
<connection>
<GID>6936</GID>
<name>clock</name></connection>
<connection>
<GID>6940</GID>
<name>clock</name></connection>
<connection>
<GID>6943</GID>
<name>clock</name></connection>
<connection>
<GID>6945</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4895</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2295.5,222,-2295.5</points>
<connection>
<GID>6913</GID>
<name>OUT</name></connection>
<connection>
<GID>6918</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6923</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6928</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6933</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6938</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6941</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6944</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6946</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4896</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2280,59,-2280</points>
<connection>
<GID>6950</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2280,53,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2264.5,53,-2264.5</points>
<connection>
<GID>6949</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4897</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2280,82,-2280</points>
<connection>
<GID>6952</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2280,76,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2264.5,76,-2264.5</points>
<connection>
<GID>6951</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4898</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2280,107,-2280</points>
<connection>
<GID>6954</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2280,101,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2264.5,101,-2264.5</points>
<connection>
<GID>6953</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4899</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2280,130,-2280</points>
<connection>
<GID>6956</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2280,124,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2264.5,124,-2264.5</points>
<connection>
<GID>6955</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4900</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2280,153,-2280</points>
<connection>
<GID>6958</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2280,147,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2264.5,147,-2264.5</points>
<connection>
<GID>6957</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4901</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2280,176,-2280</points>
<connection>
<GID>6960</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2280,170,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2264.5,170,-2264.5</points>
<connection>
<GID>6959</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4902</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2280,201,-2280</points>
<connection>
<GID>6962</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2280,195,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2264.5,195,-2264.5</points>
<connection>
<GID>6961</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4903</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2280,224,-2280</points>
<connection>
<GID>6964</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2280,218,-2264.5</points>
<intersection>-2280 1</intersection>
<intersection>-2264.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2264.5,218,-2264.5</points>
<connection>
<GID>6963</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4904</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2267.5,211,-2267.5</points>
<connection>
<GID>6947</GID>
<name>OUT</name></connection>
<connection>
<GID>6949</GID>
<name>clock</name></connection>
<connection>
<GID>6951</GID>
<name>clock</name></connection>
<connection>
<GID>6953</GID>
<name>clock</name></connection>
<connection>
<GID>6955</GID>
<name>clock</name></connection>
<connection>
<GID>6957</GID>
<name>clock</name></connection>
<connection>
<GID>6959</GID>
<name>clock</name></connection>
<connection>
<GID>6961</GID>
<name>clock</name></connection>
<connection>
<GID>6963</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4905</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2277,222,-2277</points>
<connection>
<GID>6948</GID>
<name>OUT</name></connection>
<connection>
<GID>6950</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6952</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6954</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6956</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6958</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6960</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6962</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6964</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4906</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-2346,40.5,-2181</points>
<connection>
<GID>6980</GID>
<name>N_in1</name></connection>
<connection>
<GID>6965</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 12</intersection>
<intersection>-2302 11</intersection>
<intersection>-2283 10</intersection>
<intersection>-2264.5 9</intersection>
<intersection>-2242.5 8</intersection>
<intersection>-2224 7</intersection>
<intersection>-2205 6</intersection>
<intersection>-2186.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-2186.5,46,-2186.5</points>
<connection>
<GID>7169</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40.5,-2205,46,-2205</points>
<connection>
<GID>7133</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>40.5,-2224,46,-2224</points>
<connection>
<GID>7097</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>40.5,-2242.5,46,-2242.5</points>
<connection>
<GID>7043</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>40.5,-2264.5,46,-2264.5</points>
<connection>
<GID>6949</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>40.5,-2283,46,-2283</points>
<connection>
<GID>6916</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>40.5,-2302,46,-2302</points>
<connection>
<GID>6878</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>40.5,-2320.5,46,-2320.5</points>
<connection>
<GID>7205</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4907</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-2345.5,63.5,-2180.5</points>
<connection>
<GID>6981</GID>
<name>N_in1</name></connection>
<connection>
<GID>6966</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 4</intersection>
<intersection>-2311 5</intersection>
<intersection>-2292 6</intersection>
<intersection>-2273.5 7</intersection>
<intersection>-2251.5 8</intersection>
<intersection>-2233 9</intersection>
<intersection>-2214 10</intersection>
<intersection>-2195.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>59,-2329.5,63.5,-2329.5</points>
<intersection>59 12</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>59,-2311,63.5,-2311</points>
<intersection>59 13</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59,-2292,63.5,-2292</points>
<intersection>59 14</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59,-2273.5,63.5,-2273.5</points>
<intersection>59 15</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>59,-2251.5,63.5,-2251.5</points>
<intersection>59 18</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>59,-2233,63.5,-2233</points>
<intersection>59 19</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>59,-2214,63.5,-2214</points>
<intersection>59 20</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>59,-2195.5,63.5,-2195.5</points>
<intersection>59 21</intersection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>59,-2330.5,59,-2329.5</points>
<connection>
<GID>7207</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>59,-2312,59,-2311</points>
<connection>
<GID>6880</GID>
<name>OUT_0</name></connection>
<intersection>-2311 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>59,-2293,59,-2292</points>
<connection>
<GID>6918</GID>
<name>OUT_0</name></connection>
<intersection>-2292 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>59,-2274.5,59,-2273.5</points>
<connection>
<GID>6950</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>59,-2252.5,59,-2251.5</points>
<connection>
<GID>7049</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>59,-2234,59,-2233</points>
<connection>
<GID>7099</GID>
<name>OUT_0</name></connection>
<intersection>-2233 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>59,-2215,59,-2214</points>
<connection>
<GID>7135</GID>
<name>OUT_0</name></connection>
<intersection>-2214 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>59,-2196.5,59,-2195.5</points>
<connection>
<GID>7171</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>4908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-2345.5,66.5,-2181</points>
<connection>
<GID>6982</GID>
<name>N_in1</name></connection>
<connection>
<GID>6967</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 10</intersection>
<intersection>-2302 9</intersection>
<intersection>-2283 8</intersection>
<intersection>-2264.5 7</intersection>
<intersection>-2242.5 6</intersection>
<intersection>-2224 5</intersection>
<intersection>-2205 4</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>66.5,-2186.5,69,-2186.5</points>
<connection>
<GID>7173</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-2205,69,-2205</points>
<connection>
<GID>7137</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66.5,-2224,69,-2224</points>
<connection>
<GID>7101</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66.5,-2242.5,69,-2242.5</points>
<connection>
<GID>7065</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66.5,-2264.5,69,-2264.5</points>
<connection>
<GID>6951</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-2283,69,-2283</points>
<connection>
<GID>6921</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66.5,-2302,69,-2302</points>
<connection>
<GID>6882</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>66.5,-2320.5,69,-2320.5</points>
<connection>
<GID>7209</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4909</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-2345.5,86,-2180.5</points>
<connection>
<GID>6983</GID>
<name>N_in1</name></connection>
<connection>
<GID>6968</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 6</intersection>
<intersection>-2311 7</intersection>
<intersection>-2292 8</intersection>
<intersection>-2273.5 9</intersection>
<intersection>-2251.5 10</intersection>
<intersection>-2233 11</intersection>
<intersection>-2214 12</intersection>
<intersection>-2195.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>82,-2329.5,86,-2329.5</points>
<intersection>82 14</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82,-2311,86,-2311</points>
<intersection>82 15</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>82,-2292,86,-2292</points>
<intersection>82 16</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82,-2273.5,86,-2273.5</points>
<intersection>82 17</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>82,-2251.5,86,-2251.5</points>
<intersection>82 20</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>82,-2233,86,-2233</points>
<intersection>82 21</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>82,-2214,86,-2214</points>
<intersection>82 22</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>82,-2195.5,86,-2195.5</points>
<intersection>82 23</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>82,-2330.5,82,-2329.5</points>
<connection>
<GID>7211</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>82,-2312,82,-2311</points>
<connection>
<GID>6884</GID>
<name>OUT_0</name></connection>
<intersection>-2311 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>82,-2293,82,-2292</points>
<connection>
<GID>6923</GID>
<name>OUT_0</name></connection>
<intersection>-2292 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>82,-2274.5,82,-2273.5</points>
<connection>
<GID>6952</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>82,-2252.5,82,-2251.5</points>
<connection>
<GID>7067</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>82,-2234,82,-2233</points>
<connection>
<GID>7103</GID>
<name>OUT_0</name></connection>
<intersection>-2233 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>82,-2215,82,-2214</points>
<connection>
<GID>7139</GID>
<name>OUT_0</name></connection>
<intersection>-2214 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>82,-2196.5,82,-2195.5</points>
<connection>
<GID>7175</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-2345.5,89.5,-2180.5</points>
<connection>
<GID>6984</GID>
<name>N_in1</name></connection>
<connection>
<GID>6969</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 13</intersection>
<intersection>-2302 12</intersection>
<intersection>-2283 11</intersection>
<intersection>-2264.5 10</intersection>
<intersection>-2242.5 9</intersection>
<intersection>-2224 8</intersection>
<intersection>-2205 7</intersection>
<intersection>-2186.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-2186.5,94,-2186.5</points>
<connection>
<GID>7177</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-2205,94,-2205</points>
<connection>
<GID>7141</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89.5,-2224,94,-2224</points>
<connection>
<GID>7105</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-2242.5,94,-2242.5</points>
<connection>
<GID>7069</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>89.5,-2264.5,94,-2264.5</points>
<connection>
<GID>6953</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89.5,-2283,94,-2283</points>
<connection>
<GID>6926</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>89.5,-2302,94,-2302</points>
<connection>
<GID>6886</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>89.5,-2320.5,94,-2320.5</points>
<connection>
<GID>7213</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-2345.5,110.5,-2181</points>
<connection>
<GID>6985</GID>
<name>N_in1</name></connection>
<connection>
<GID>6970</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 6</intersection>
<intersection>-2311 7</intersection>
<intersection>-2292 8</intersection>
<intersection>-2273.5 9</intersection>
<intersection>-2251.5 10</intersection>
<intersection>-2233 11</intersection>
<intersection>-2214 12</intersection>
<intersection>-2195.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>107,-2329.5,110.5,-2329.5</points>
<intersection>107 14</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>107,-2311,110.5,-2311</points>
<intersection>107 15</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>107,-2292,110.5,-2292</points>
<intersection>107 16</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>107,-2273.5,110.5,-2273.5</points>
<intersection>107 17</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>107,-2251.5,110.5,-2251.5</points>
<intersection>107 20</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>107,-2233,110.5,-2233</points>
<intersection>107 21</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>107,-2214,110.5,-2214</points>
<intersection>107 22</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>107,-2195.5,110.5,-2195.5</points>
<intersection>107 23</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>107,-2330.5,107,-2329.5</points>
<connection>
<GID>7215</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>107,-2312,107,-2311</points>
<connection>
<GID>6888</GID>
<name>OUT_0</name></connection>
<intersection>-2311 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>107,-2293,107,-2292</points>
<connection>
<GID>6928</GID>
<name>OUT_0</name></connection>
<intersection>-2292 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>107,-2274.5,107,-2273.5</points>
<connection>
<GID>6954</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>107,-2252.5,107,-2251.5</points>
<connection>
<GID>7071</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>107,-2234,107,-2233</points>
<connection>
<GID>7107</GID>
<name>OUT_0</name></connection>
<intersection>-2233 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>107,-2215,107,-2214</points>
<connection>
<GID>7143</GID>
<name>OUT_0</name></connection>
<intersection>-2214 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>107,-2196.5,107,-2195.5</points>
<connection>
<GID>7179</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2345.5,114.5,-2180.5</points>
<connection>
<GID>6986</GID>
<name>N_in1</name></connection>
<connection>
<GID>6971</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 13</intersection>
<intersection>-2302 12</intersection>
<intersection>-2283 11</intersection>
<intersection>-2264.5 10</intersection>
<intersection>-2242.5 9</intersection>
<intersection>-2224 8</intersection>
<intersection>-2205 7</intersection>
<intersection>-2186.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>114.5,-2186.5,117,-2186.5</points>
<connection>
<GID>7181</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-2205,117,-2205</points>
<connection>
<GID>7145</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-2224,117,-2224</points>
<connection>
<GID>7109</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114.5,-2242.5,117,-2242.5</points>
<connection>
<GID>7073</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114.5,-2264.5,117,-2264.5</points>
<connection>
<GID>6955</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>114.5,-2283,117,-2283</points>
<connection>
<GID>6931</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114.5,-2302,117,-2302</points>
<connection>
<GID>6890</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>114.5,-2320.5,117,-2320.5</points>
<connection>
<GID>6854</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4913</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-2345.5,133,-2180.5</points>
<connection>
<GID>6987</GID>
<name>N_in1</name></connection>
<connection>
<GID>6972</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 6</intersection>
<intersection>-2311 7</intersection>
<intersection>-2292 8</intersection>
<intersection>-2273.5 9</intersection>
<intersection>-2251.5 10</intersection>
<intersection>-2233 11</intersection>
<intersection>-2214 12</intersection>
<intersection>-2195.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>130,-2329.5,133,-2329.5</points>
<intersection>130 14</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-2311,133,-2311</points>
<intersection>130 15</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>130,-2292,133,-2292</points>
<intersection>130 16</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>130,-2273.5,133,-2273.5</points>
<intersection>130 17</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>130,-2251.5,133,-2251.5</points>
<intersection>130 20</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>130,-2233,133,-2233</points>
<intersection>130 21</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>130,-2214,133,-2214</points>
<intersection>130 22</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>130,-2195.5,133,-2195.5</points>
<intersection>130 23</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>130,-2330.5,130,-2329.5</points>
<connection>
<GID>6856</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>130,-2312,130,-2311</points>
<connection>
<GID>6892</GID>
<name>OUT_0</name></connection>
<intersection>-2311 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>130,-2293,130,-2292</points>
<connection>
<GID>6933</GID>
<name>OUT_0</name></connection>
<intersection>-2292 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>130,-2274.5,130,-2273.5</points>
<connection>
<GID>6956</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>130,-2252.5,130,-2251.5</points>
<connection>
<GID>7075</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>130,-2234,130,-2233</points>
<connection>
<GID>7111</GID>
<name>OUT_0</name></connection>
<intersection>-2233 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>130,-2215,130,-2214</points>
<connection>
<GID>7147</GID>
<name>OUT_0</name></connection>
<intersection>-2214 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>130,-2196.5,130,-2195.5</points>
<connection>
<GID>7183</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4914</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2345.5,137,-2180.5</points>
<connection>
<GID>6988</GID>
<name>N_in1</name></connection>
<connection>
<GID>6973</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 13</intersection>
<intersection>-2302 12</intersection>
<intersection>-2283 11</intersection>
<intersection>-2264.5 10</intersection>
<intersection>-2242.5 9</intersection>
<intersection>-2224 8</intersection>
<intersection>-2205 7</intersection>
<intersection>-2186.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>137,-2186.5,140,-2186.5</points>
<connection>
<GID>7185</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137,-2205,140,-2205</points>
<connection>
<GID>7149</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-2224,140,-2224</points>
<connection>
<GID>7113</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137,-2242.5,140,-2242.5</points>
<connection>
<GID>7077</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-2264.5,140,-2264.5</points>
<connection>
<GID>6957</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>137,-2283,140,-2283</points>
<connection>
<GID>6936</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137,-2302,140,-2302</points>
<connection>
<GID>6894</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-2320.5,140,-2320.5</points>
<connection>
<GID>6858</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>4915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-2345,156,-2180.5</points>
<connection>
<GID>6989</GID>
<name>N_in1</name></connection>
<connection>
<GID>6974</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 6</intersection>
<intersection>-2311 7</intersection>
<intersection>-2292 8</intersection>
<intersection>-2273.5 9</intersection>
<intersection>-2251.5 10</intersection>
<intersection>-2233 11</intersection>
<intersection>-2214 12</intersection>
<intersection>-2195.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>153,-2329.5,156,-2329.5</points>
<intersection>153 14</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>153,-2311,156,-2311</points>
<intersection>153 15</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>153,-2292,156,-2292</points>
<intersection>153 16</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>153,-2273.5,156,-2273.5</points>
<intersection>153 17</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>153,-2251.5,156,-2251.5</points>
<intersection>153 20</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>153,-2233,156,-2233</points>
<intersection>153 21</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>153,-2214,156,-2214</points>
<intersection>153 22</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>153,-2195.5,156,-2195.5</points>
<intersection>153 23</intersection>
<intersection>156 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>153,-2330.5,153,-2329.5</points>
<connection>
<GID>6860</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>153,-2312,153,-2311</points>
<connection>
<GID>6896</GID>
<name>OUT_0</name></connection>
<intersection>-2311 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>153,-2293,153,-2292</points>
<connection>
<GID>6938</GID>
<name>OUT_0</name></connection>
<intersection>-2292 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>153,-2274.5,153,-2273.5</points>
<connection>
<GID>6958</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>153,-2252.5,153,-2251.5</points>
<connection>
<GID>7079</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>153,-2234,153,-2233</points>
<connection>
<GID>7115</GID>
<name>OUT_0</name></connection>
<intersection>-2233 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>153,-2215,153,-2214</points>
<connection>
<GID>7151</GID>
<name>OUT_0</name></connection>
<intersection>-2214 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>153,-2196.5,153,-2195.5</points>
<connection>
<GID>7187</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-2345,161,-2180.5</points>
<connection>
<GID>6990</GID>
<name>N_in1</name></connection>
<connection>
<GID>6975</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 13</intersection>
<intersection>-2302 12</intersection>
<intersection>-2283 11</intersection>
<intersection>-2264.5 10</intersection>
<intersection>-2242.5 9</intersection>
<intersection>-2224 8</intersection>
<intersection>-2205 7</intersection>
<intersection>-2186.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>161,-2186.5,163,-2186.5</points>
<connection>
<GID>7189</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>161,-2205,163,-2205</points>
<connection>
<GID>7153</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>161,-2224,163,-2224</points>
<connection>
<GID>7117</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>161,-2242.5,163,-2242.5</points>
<connection>
<GID>7081</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>161,-2264.5,163,-2264.5</points>
<connection>
<GID>6959</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>161,-2283,163,-2283</points>
<connection>
<GID>6940</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>161,-2302,163,-2302</points>
<connection>
<GID>6898</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>161,-2320.5,163,-2320.5</points>
<connection>
<GID>6862</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>4917</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-2344.5,179,-2180.5</points>
<connection>
<GID>6991</GID>
<name>N_in1</name></connection>
<connection>
<GID>6977</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 16</intersection>
<intersection>-2311 15</intersection>
<intersection>-2292 14</intersection>
<intersection>-2273.5 13</intersection>
<intersection>-2251.5 12</intersection>
<intersection>-2233 11</intersection>
<intersection>-2214 10</intersection>
<intersection>-2195.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>176,-2195.5,179,-2195.5</points>
<intersection>176 26</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>176,-2214,179,-2214</points>
<intersection>176 25</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>176,-2233,179,-2233</points>
<intersection>176 24</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>176,-2251.5,179,-2251.5</points>
<intersection>176 23</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>176,-2273.5,179,-2273.5</points>
<intersection>176 20</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>176,-2292,179,-2292</points>
<intersection>176 19</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>176,-2311,179,-2311</points>
<intersection>176 18</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>176,-2329.5,179,-2329.5</points>
<intersection>176 17</intersection>
<intersection>179 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>176,-2330.5,176,-2329.5</points>
<connection>
<GID>6864</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>176,-2312,176,-2311</points>
<connection>
<GID>6900</GID>
<name>OUT_0</name></connection>
<intersection>-2311 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>176,-2293,176,-2292</points>
<connection>
<GID>6941</GID>
<name>OUT_0</name></connection>
<intersection>-2292 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>176,-2274.5,176,-2273.5</points>
<connection>
<GID>6960</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>176,-2252.5,176,-2251.5</points>
<connection>
<GID>7083</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>176,-2234,176,-2233</points>
<connection>
<GID>7119</GID>
<name>OUT_0</name></connection>
<intersection>-2233 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>176,-2215,176,-2214</points>
<connection>
<GID>7155</GID>
<name>OUT_0</name></connection>
<intersection>-2214 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>176,-2196.5,176,-2195.5</points>
<connection>
<GID>7191</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>4918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2344.5,183.5,-2180.5</points>
<connection>
<GID>6992</GID>
<name>N_in1</name></connection>
<connection>
<GID>6976</GID>
<name>N_in0</name></connection>
<intersection>-2320.5 13</intersection>
<intersection>-2302 12</intersection>
<intersection>-2283 11</intersection>
<intersection>-2264.5 10</intersection>
<intersection>-2242.5 9</intersection>
<intersection>-2224 8</intersection>
<intersection>-2205 7</intersection>
<intersection>-2186.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>183.5,-2186.5,188,-2186.5</points>
<connection>
<GID>7193</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>183.5,-2205,188,-2205</points>
<connection>
<GID>7157</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>183.5,-2224,188,-2224</points>
<connection>
<GID>7121</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>183.5,-2242.5,188,-2242.5</points>
<connection>
<GID>7085</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183.5,-2264.5,188,-2264.5</points>
<connection>
<GID>6961</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183.5,-2283,188,-2283</points>
<connection>
<GID>6943</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183.5,-2302,188,-2302</points>
<connection>
<GID>6902</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183.5,-2320.5,188,-2320.5</points>
<connection>
<GID>6866</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-2344,204.5,-2181</points>
<connection>
<GID>6993</GID>
<name>N_in1</name></connection>
<connection>
<GID>6978</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 6</intersection>
<intersection>-2311 7</intersection>
<intersection>-2292 8</intersection>
<intersection>-2273.5 9</intersection>
<intersection>-2251.5 10</intersection>
<intersection>-2233 11</intersection>
<intersection>-2214 12</intersection>
<intersection>-2195.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>201,-2329.5,204.5,-2329.5</points>
<intersection>201 14</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>201,-2311,204.5,-2311</points>
<intersection>201 15</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>201,-2292,204.5,-2292</points>
<intersection>201 16</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>201,-2273.5,204.5,-2273.5</points>
<intersection>201 17</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>201,-2251.5,204.5,-2251.5</points>
<intersection>201 20</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>201,-2233,204.5,-2233</points>
<intersection>201 21</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>201,-2214,204.5,-2214</points>
<intersection>201 22</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>201,-2195.5,204.5,-2195.5</points>
<intersection>201 23</intersection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>201,-2330.5,201,-2329.5</points>
<connection>
<GID>6868</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201,-2312,201,-2311</points>
<connection>
<GID>6904</GID>
<name>OUT_0</name></connection>
<intersection>-2311 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>201,-2293,201,-2292</points>
<connection>
<GID>6944</GID>
<name>OUT_0</name></connection>
<intersection>-2292 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>201,-2274.5,201,-2273.5</points>
<connection>
<GID>6962</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>201,-2252.5,201,-2251.5</points>
<connection>
<GID>7087</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>201,-2234,201,-2233</points>
<connection>
<GID>7123</GID>
<name>OUT_0</name></connection>
<intersection>-2233 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>201,-2215,201,-2214</points>
<connection>
<GID>7159</GID>
<name>OUT_0</name></connection>
<intersection>-2214 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>201,-2196.5,201,-2195.5</points>
<connection>
<GID>7195</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>4920</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-2344,208,-2181</points>
<connection>
<GID>6995</GID>
<name>N_in0</name></connection>
<connection>
<GID>6994</GID>
<name>N_in1</name></connection>
<intersection>-2320.5 11</intersection>
<intersection>-2302 10</intersection>
<intersection>-2283 9</intersection>
<intersection>-2264.5 7</intersection>
<intersection>-2242.5 6</intersection>
<intersection>-2224 5</intersection>
<intersection>-2205 4</intersection>
<intersection>-2186.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208,-2186.5,211,-2186.5</points>
<connection>
<GID>7197</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208,-2205,211,-2205</points>
<connection>
<GID>7161</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>208,-2224,211,-2224</points>
<connection>
<GID>7125</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>208,-2242.5,211,-2242.5</points>
<connection>
<GID>7089</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>208,-2264.5,211,-2264.5</points>
<connection>
<GID>6963</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>208,-2283,211,-2283</points>
<connection>
<GID>6945</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>208,-2302,211,-2302</points>
<connection>
<GID>6906</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>208,-2320.5,211,-2320.5</points>
<connection>
<GID>6870</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>4921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-2344,229,-2182</points>
<connection>
<GID>6996</GID>
<name>N_in1</name></connection>
<connection>
<GID>6979</GID>
<name>N_in0</name></connection>
<intersection>-2329.5 11</intersection>
<intersection>-2311 10</intersection>
<intersection>-2292 9</intersection>
<intersection>-2273.5 8</intersection>
<intersection>-2251.5 7</intersection>
<intersection>-2233 6</intersection>
<intersection>-2214 5</intersection>
<intersection>-2195.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>224,-2195.5,229,-2195.5</points>
<intersection>224 21</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>224,-2214,229,-2214</points>
<intersection>224 20</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>224,-2233,229,-2233</points>
<intersection>224 19</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>224,-2251.5,229,-2251.5</points>
<intersection>224 18</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>224,-2273.5,229,-2273.5</points>
<intersection>224 15</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>224,-2292,229,-2292</points>
<intersection>224 14</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>224,-2311,229,-2311</points>
<intersection>224 13</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>224,-2329.5,229,-2329.5</points>
<intersection>224 12</intersection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>224,-2330.5,224,-2329.5</points>
<connection>
<GID>6872</GID>
<name>OUT_0</name></connection>
<intersection>-2329.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>224,-2312,224,-2311</points>
<connection>
<GID>6908</GID>
<name>OUT_0</name></connection>
<intersection>-2311 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>224,-2293,224,-2292</points>
<connection>
<GID>6946</GID>
<name>OUT_0</name></connection>
<intersection>-2292 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>224,-2274.5,224,-2273.5</points>
<connection>
<GID>6964</GID>
<name>OUT_0</name></connection>
<intersection>-2273.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>224,-2252.5,224,-2251.5</points>
<connection>
<GID>7091</GID>
<name>OUT_0</name></connection>
<intersection>-2251.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>224,-2234,224,-2233</points>
<connection>
<GID>7127</GID>
<name>OUT_0</name></connection>
<intersection>-2233 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>224,-2215,224,-2214</points>
<connection>
<GID>7163</GID>
<name>OUT_0</name></connection>
<intersection>-2214 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>224,-2196.5,224,-2195.5</points>
<connection>
<GID>7199</GID>
<name>OUT_0</name></connection>
<intersection>-2195.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>4922</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-128,-2188.5,18.5,-2188.5</points>
<connection>
<GID>7165</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-2340,-128,-2188.5</points>
<connection>
<GID>7002</GID>
<name>OUT_15</name></connection>
<intersection>-2198 4</intersection>
<intersection>-2188.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-2198,30,-2198</points>
<connection>
<GID>7167</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>4923</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-127,-2207,18.5,-2207</points>
<connection>
<GID>7129</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-127,-2341,-127,-2207</points>
<intersection>-2341 6</intersection>
<intersection>-2216.5 5</intersection>
<intersection>-2207 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-127,-2216.5,30,-2216.5</points>
<connection>
<GID>7131</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2341,-127,-2341</points>
<connection>
<GID>7002</GID>
<name>OUT_14</name></connection>
<intersection>-127 4</intersection></hsegment></shape></wire>
<wire>
<ID>4924</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-126,-2226,18.5,-2226</points>
<connection>
<GID>7093</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-2342,-126,-2226</points>
<intersection>-2342 6</intersection>
<intersection>-2235.5 4</intersection>
<intersection>-2226 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-2235.5,30,-2235.5</points>
<connection>
<GID>7095</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2342,-126,-2342</points>
<connection>
<GID>7002</GID>
<name>OUT_13</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>4925</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-125,-2244.5,18.5,-2244.5</points>
<connection>
<GID>7033</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-125,-2343,-125,-2244.5</points>
<intersection>-2343 5</intersection>
<intersection>-2254 4</intersection>
<intersection>-2244.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-125,-2254,30,-2254</points>
<connection>
<GID>7038</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2343,-125,-2343</points>
<connection>
<GID>7002</GID>
<name>OUT_12</name></connection>
<intersection>-125 3</intersection></hsegment></shape></wire>
<wire>
<ID>4926</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,-2266.5,18.5,-2266.5</points>
<connection>
<GID>6947</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-2344,-124,-2266.5</points>
<intersection>-2344 6</intersection>
<intersection>-2276 4</intersection>
<intersection>-2266.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-2276,29.5,-2276</points>
<connection>
<GID>6948</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2344,-124,-2344</points>
<connection>
<GID>7002</GID>
<name>OUT_11</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>4927</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123,-2285,18.5,-2285</points>
<connection>
<GID>6911</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-2345,-123,-2285</points>
<intersection>-2345 5</intersection>
<intersection>-2294.5 4</intersection>
<intersection>-2285 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-2294.5,29.5,-2294.5</points>
<connection>
<GID>6913</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2345,-123,-2345</points>
<connection>
<GID>7002</GID>
<name>OUT_10</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>4928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-2304,18.5,-2304</points>
<connection>
<GID>6874</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-2346,-122,-2304</points>
<intersection>-2346 5</intersection>
<intersection>-2313.5 4</intersection>
<intersection>-2304 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-2313.5,29.5,-2313.5</points>
<connection>
<GID>6876</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2346,-122,-2346</points>
<connection>
<GID>7002</GID>
<name>OUT_9</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>4929</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-2322.5,18.5,-2322.5</points>
<connection>
<GID>7201</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-2347,-121,-2322.5</points>
<intersection>-2347 5</intersection>
<intersection>-2332 4</intersection>
<intersection>-2322.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-2332,29.5,-2332</points>
<connection>
<GID>7203</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2347,-121,-2347</points>
<connection>
<GID>7002</GID>
<name>OUT_8</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>4930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-2346,17.5,-2181</points>
<connection>
<GID>7000</GID>
<name>N_in1</name></connection>
<connection>
<GID>6998</GID>
<name>N_in0</name></connection>
<intersection>-2324.5 10</intersection>
<intersection>-2306 9</intersection>
<intersection>-2287 8</intersection>
<intersection>-2268.5 7</intersection>
<intersection>-2246.5 6</intersection>
<intersection>-2228 5</intersection>
<intersection>-2209 4</intersection>
<intersection>-2190.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-2190.5,18.5,-2190.5</points>
<connection>
<GID>7165</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-2209,18.5,-2209</points>
<connection>
<GID>7129</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>17.5,-2228,18.5,-2228</points>
<connection>
<GID>7093</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>17.5,-2246.5,18.5,-2246.5</points>
<connection>
<GID>7033</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>17.5,-2268.5,18.5,-2268.5</points>
<connection>
<GID>6947</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>17.5,-2287,18.5,-2287</points>
<connection>
<GID>6911</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>17.5,-2306,18.5,-2306</points>
<connection>
<GID>6874</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>17.5,-2324.5,18.5,-2324.5</points>
<connection>
<GID>7201</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-2346,27.5,-2181</points>
<connection>
<GID>6999</GID>
<name>N_in1</name></connection>
<connection>
<GID>6997</GID>
<name>N_in0</name></connection>
<intersection>-2334 3</intersection>
<intersection>-2315.5 5</intersection>
<intersection>-2296.5 7</intersection>
<intersection>-2278 9</intersection>
<intersection>-2256 11</intersection>
<intersection>-2237.5 13</intersection>
<intersection>-2218.5 15</intersection>
<intersection>-2200 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-2334,29.5,-2334</points>
<connection>
<GID>7203</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-2315.5,29.5,-2315.5</points>
<connection>
<GID>6876</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-2296.5,29.5,-2296.5</points>
<connection>
<GID>6913</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>27.5,-2278,29.5,-2278</points>
<connection>
<GID>6948</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>27.5,-2256,30,-2256</points>
<connection>
<GID>7038</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>27.5,-2237.5,30,-2237.5</points>
<connection>
<GID>7095</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>27.5,-2218.5,30,-2218.5</points>
<connection>
<GID>7131</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>27.5,-2200,30,-2200</points>
<connection>
<GID>7167</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4932</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2433.5,59,-2433.5</points>
<connection>
<GID>7098</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2433.5,53,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2418,53,-2418</points>
<connection>
<GID>7086</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4933</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2433.5,82,-2433.5</points>
<connection>
<GID>7124</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2433.5,76,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2418,76,-2418</points>
<connection>
<GID>7122</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4934</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2433.5,107,-2433.5</points>
<connection>
<GID>7132</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2433.5,101,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2418,101,-2418</points>
<connection>
<GID>7128</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4935</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2433.5,130,-2433.5</points>
<connection>
<GID>7140</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2433.5,124,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2418,124,-2418</points>
<connection>
<GID>7136</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4936</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2433.5,153,-2433.5</points>
<connection>
<GID>7146</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2433.5,147,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2418,147,-2418</points>
<connection>
<GID>7142</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4937</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2433.5,176,-2433.5</points>
<connection>
<GID>7150</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2433.5,170,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2418,170,-2418</points>
<connection>
<GID>7148</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4938</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2433.5,201,-2433.5</points>
<connection>
<GID>7154</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2433.5,195,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2418,195,-2418</points>
<connection>
<GID>7152</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4939</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2433.5,224,-2433.5</points>
<connection>
<GID>7158</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2433.5,218,-2418</points>
<intersection>-2433.5 1</intersection>
<intersection>-2418 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2418,218,-2418</points>
<connection>
<GID>7156</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4940</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2421,211,-2421</points>
<connection>
<GID>7080</GID>
<name>OUT</name></connection>
<connection>
<GID>7086</GID>
<name>clock</name></connection>
<connection>
<GID>7122</GID>
<name>clock</name></connection>
<connection>
<GID>7128</GID>
<name>clock</name></connection>
<connection>
<GID>7136</GID>
<name>clock</name></connection>
<connection>
<GID>7142</GID>
<name>clock</name></connection>
<connection>
<GID>7148</GID>
<name>clock</name></connection>
<connection>
<GID>7152</GID>
<name>clock</name></connection>
<connection>
<GID>7156</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4941</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2430.5,222,-2430.5</points>
<connection>
<GID>7082</GID>
<name>OUT</name></connection>
<connection>
<GID>7098</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7124</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7132</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7140</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7146</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7150</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7154</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7158</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2415,59,-2415</points>
<connection>
<GID>7166</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2415,53,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2399.5,53,-2399.5</points>
<connection>
<GID>7164</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4943</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2415,82,-2415</points>
<connection>
<GID>7170</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2415,76,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2399.5,76,-2399.5</points>
<connection>
<GID>7168</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4944</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2415,107,-2415</points>
<connection>
<GID>7174</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2415,101,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2399.5,101,-2399.5</points>
<connection>
<GID>7172</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4945</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2415,130,-2415</points>
<connection>
<GID>7178</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2415,124,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2399.5,124,-2399.5</points>
<connection>
<GID>7176</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4946</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2415,153,-2415</points>
<connection>
<GID>7182</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2415,147,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2399.5,147,-2399.5</points>
<connection>
<GID>7180</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4947</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2415,176,-2415</points>
<connection>
<GID>7186</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2415,170,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2399.5,170,-2399.5</points>
<connection>
<GID>7184</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4948</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2415,201,-2415</points>
<connection>
<GID>7190</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2415,195,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2399.5,195,-2399.5</points>
<connection>
<GID>7188</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4949</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2415,224,-2415</points>
<connection>
<GID>7194</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2415,218,-2399.5</points>
<intersection>-2415 1</intersection>
<intersection>-2399.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2399.5,218,-2399.5</points>
<connection>
<GID>7192</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4950</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2402.5,211,-2402.5</points>
<connection>
<GID>7160</GID>
<name>OUT</name></connection>
<connection>
<GID>7164</GID>
<name>clock</name></connection>
<connection>
<GID>7168</GID>
<name>clock</name></connection>
<connection>
<GID>7172</GID>
<name>clock</name></connection>
<connection>
<GID>7176</GID>
<name>clock</name></connection>
<connection>
<GID>7180</GID>
<name>clock</name></connection>
<connection>
<GID>7184</GID>
<name>clock</name></connection>
<connection>
<GID>7188</GID>
<name>clock</name></connection>
<connection>
<GID>7192</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4951</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2412,222,-2412</points>
<connection>
<GID>7162</GID>
<name>OUT</name></connection>
<connection>
<GID>7166</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7170</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7174</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7178</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7182</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7186</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7190</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7194</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4952</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2396,59,-2396</points>
<connection>
<GID>7202</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2396,53,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2380.5,53,-2380.5</points>
<connection>
<GID>7200</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4953</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2396,82,-2396</points>
<connection>
<GID>7206</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2396,76,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2380.5,76,-2380.5</points>
<connection>
<GID>7204</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2396,107,-2396</points>
<connection>
<GID>7210</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2396,101,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2380.5,101,-2380.5</points>
<connection>
<GID>7208</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4955</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2396,130,-2396</points>
<connection>
<GID>7214</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2396,124,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2380.5,124,-2380.5</points>
<connection>
<GID>7212</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4956</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2396,153,-2396</points>
<connection>
<GID>6855</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2396,147,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2380.5,147,-2380.5</points>
<connection>
<GID>7216</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4957</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2396,176,-2396</points>
<connection>
<GID>6859</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2396,170,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2380.5,170,-2380.5</points>
<connection>
<GID>6857</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4958</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2396,201,-2396</points>
<connection>
<GID>6863</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2396,195,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2380.5,195,-2380.5</points>
<connection>
<GID>6861</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2396,224,-2396</points>
<connection>
<GID>6867</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2396,218,-2380.5</points>
<intersection>-2396 1</intersection>
<intersection>-2380.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2380.5,218,-2380.5</points>
<connection>
<GID>6865</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4960</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2383.5,211,-2383.5</points>
<connection>
<GID>7216</GID>
<name>clock</name></connection>
<connection>
<GID>7212</GID>
<name>clock</name></connection>
<connection>
<GID>7208</GID>
<name>clock</name></connection>
<connection>
<GID>7204</GID>
<name>clock</name></connection>
<connection>
<GID>7200</GID>
<name>clock</name></connection>
<connection>
<GID>7196</GID>
<name>OUT</name></connection>
<connection>
<GID>6865</GID>
<name>clock</name></connection>
<connection>
<GID>6861</GID>
<name>clock</name></connection>
<connection>
<GID>6857</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4961</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2393,222,-2393</points>
<connection>
<GID>7214</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7210</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7206</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7202</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7198</GID>
<name>OUT</name></connection>
<connection>
<GID>6867</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6863</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6859</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6855</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4962</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2377.5,59,-2377.5</points>
<connection>
<GID>6875</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2377.5,53,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2362,53,-2362</points>
<connection>
<GID>6873</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4963</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2377.5,82,-2377.5</points>
<connection>
<GID>6879</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2377.5,76,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2362,76,-2362</points>
<connection>
<GID>6877</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4964</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2377.5,107,-2377.5</points>
<connection>
<GID>6883</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2377.5,101,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2362,101,-2362</points>
<connection>
<GID>6881</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4965</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2377.5,130,-2377.5</points>
<connection>
<GID>6887</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2377.5,124,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2362,124,-2362</points>
<connection>
<GID>6885</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2377.5,153,-2377.5</points>
<connection>
<GID>6891</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2377.5,147,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2362,147,-2362</points>
<connection>
<GID>6889</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4967</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2377.5,176,-2377.5</points>
<connection>
<GID>6895</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2377.5,170,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2362,170,-2362</points>
<connection>
<GID>6893</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4968</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2377.5,201,-2377.5</points>
<connection>
<GID>6899</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2377.5,195,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2362,195,-2362</points>
<connection>
<GID>6897</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2377.5,224,-2377.5</points>
<connection>
<GID>6903</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2377.5,218,-2362</points>
<intersection>-2377.5 1</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2362,218,-2362</points>
<connection>
<GID>6901</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4970</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2365,211,-2365</points>
<connection>
<GID>6869</GID>
<name>OUT</name></connection>
<connection>
<GID>6873</GID>
<name>clock</name></connection>
<connection>
<GID>6877</GID>
<name>clock</name></connection>
<connection>
<GID>6881</GID>
<name>clock</name></connection>
<connection>
<GID>6885</GID>
<name>clock</name></connection>
<connection>
<GID>6889</GID>
<name>clock</name></connection>
<connection>
<GID>6893</GID>
<name>clock</name></connection>
<connection>
<GID>6897</GID>
<name>clock</name></connection>
<connection>
<GID>6901</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4971</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-2374.5,222,-2374.5</points>
<connection>
<GID>6871</GID>
<name>OUT</name></connection>
<connection>
<GID>6875</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6879</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6883</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6887</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6891</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6895</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6899</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6903</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4972</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2511.5,59,-2511.5</points>
<connection>
<GID>6912</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2511.5,53,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2496,53,-2496</points>
<connection>
<GID>6909</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2511.5,82,-2511.5</points>
<connection>
<GID>6917</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2511.5,76,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2496,76,-2496</points>
<connection>
<GID>6914</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2511.5,107,-2511.5</points>
<connection>
<GID>6922</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2511.5,101,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2496,101,-2496</points>
<connection>
<GID>6919</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4975</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2511.5,130,-2511.5</points>
<connection>
<GID>6927</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2511.5,124,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2496,124,-2496</points>
<connection>
<GID>6924</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4976</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2511.5,153,-2511.5</points>
<connection>
<GID>6932</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2511.5,147,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2496,147,-2496</points>
<connection>
<GID>6929</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4977</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2511.5,176,-2511.5</points>
<connection>
<GID>6937</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2511.5,170,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2496,170,-2496</points>
<connection>
<GID>6934</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4978</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2511.5,201,-2511.5</points>
<connection>
<GID>7004</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2511.5,195,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2496,195,-2496</points>
<connection>
<GID>7003</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4979</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2511.5,224,-2511.5</points>
<connection>
<GID>7006</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2511.5,218,-2496</points>
<intersection>-2511.5 1</intersection>
<intersection>-2496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2496,218,-2496</points>
<connection>
<GID>7005</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4980</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2499,211,-2499</points>
<connection>
<GID>6905</GID>
<name>OUT</name></connection>
<connection>
<GID>6909</GID>
<name>clock</name></connection>
<connection>
<GID>6914</GID>
<name>clock</name></connection>
<connection>
<GID>6919</GID>
<name>clock</name></connection>
<connection>
<GID>6924</GID>
<name>clock</name></connection>
<connection>
<GID>6929</GID>
<name>clock</name></connection>
<connection>
<GID>6934</GID>
<name>clock</name></connection>
<connection>
<GID>7003</GID>
<name>clock</name></connection>
<connection>
<GID>7005</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4981</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2508.5,222,-2508.5</points>
<connection>
<GID>6907</GID>
<name>OUT</name></connection>
<connection>
<GID>6912</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6917</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6922</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6927</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6932</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6937</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7004</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7006</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4982</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2493,59,-2493</points>
<connection>
<GID>7010</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2493,53,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2477.5,53,-2477.5</points>
<connection>
<GID>7009</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4983</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2493,82,-2493</points>
<connection>
<GID>7012</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2493,76,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2477.5,76,-2477.5</points>
<connection>
<GID>7011</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4984</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2493,107,-2493</points>
<connection>
<GID>7014</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2493,101,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2477.5,101,-2477.5</points>
<connection>
<GID>7013</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4985</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2493,130,-2493</points>
<connection>
<GID>7016</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2493,124,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2477.5,124,-2477.5</points>
<connection>
<GID>7015</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4986</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2493,153,-2493</points>
<connection>
<GID>7018</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2493,147,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2477.5,147,-2477.5</points>
<connection>
<GID>7017</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4987</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2493,176,-2493</points>
<connection>
<GID>7020</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2493,170,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2477.5,170,-2477.5</points>
<connection>
<GID>7019</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4988</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2493,201,-2493</points>
<connection>
<GID>7022</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2493,195,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2477.5,195,-2477.5</points>
<connection>
<GID>7021</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4989</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2493,224,-2493</points>
<connection>
<GID>7024</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2493,218,-2477.5</points>
<intersection>-2493 1</intersection>
<intersection>-2477.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2477.5,218,-2477.5</points>
<connection>
<GID>7023</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>4990</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2480.5,211,-2480.5</points>
<connection>
<GID>7007</GID>
<name>OUT</name></connection>
<connection>
<GID>7009</GID>
<name>clock</name></connection>
<connection>
<GID>7011</GID>
<name>clock</name></connection>
<connection>
<GID>7013</GID>
<name>clock</name></connection>
<connection>
<GID>7015</GID>
<name>clock</name></connection>
<connection>
<GID>7017</GID>
<name>clock</name></connection>
<connection>
<GID>7019</GID>
<name>clock</name></connection>
<connection>
<GID>7021</GID>
<name>clock</name></connection>
<connection>
<GID>7023</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4991</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2490,222,-2490</points>
<connection>
<GID>7008</GID>
<name>OUT</name></connection>
<connection>
<GID>7010</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7012</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7014</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7016</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7018</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7020</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7022</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7024</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4992</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2474,59,-2474</points>
<connection>
<GID>6920</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2474,53,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2458.5,53,-2458.5</points>
<connection>
<GID>6915</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>4993</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2474,82,-2474</points>
<connection>
<GID>6930</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2474,76,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2458.5,76,-2458.5</points>
<connection>
<GID>6925</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>4994</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2474,107,-2474</points>
<connection>
<GID>6939</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2474,101,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2458.5,101,-2458.5</points>
<connection>
<GID>6935</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>4995</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2474,130,-2474</points>
<connection>
<GID>7026</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2474,124,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2458.5,124,-2458.5</points>
<connection>
<GID>6942</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>4996</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2474,153,-2474</points>
<connection>
<GID>7028</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2474,147,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2458.5,147,-2458.5</points>
<connection>
<GID>7027</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>4997</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2474,176,-2474</points>
<connection>
<GID>7030</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2474,170,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2458.5,170,-2458.5</points>
<connection>
<GID>7029</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>4998</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2474,201,-2474</points>
<connection>
<GID>7032</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2474,195,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2458.5,195,-2458.5</points>
<connection>
<GID>7031</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>4999</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2474,224,-2474</points>
<connection>
<GID>7035</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2474,218,-2458.5</points>
<intersection>-2474 1</intersection>
<intersection>-2458.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2458.5,218,-2458.5</points>
<connection>
<GID>7034</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>5000</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2461.5,211,-2461.5</points>
<connection>
<GID>7034</GID>
<name>clock</name></connection>
<connection>
<GID>7031</GID>
<name>clock</name></connection>
<connection>
<GID>7029</GID>
<name>clock</name></connection>
<connection>
<GID>7027</GID>
<name>clock</name></connection>
<connection>
<GID>7025</GID>
<name>OUT</name></connection>
<connection>
<GID>6942</GID>
<name>clock</name></connection>
<connection>
<GID>6935</GID>
<name>clock</name></connection>
<connection>
<GID>6925</GID>
<name>clock</name></connection>
<connection>
<GID>6915</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5001</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2471,222,-2471</points>
<connection>
<GID>6910</GID>
<name>OUT</name></connection>
<connection>
<GID>6920</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6930</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>6939</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7026</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7028</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7030</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7032</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7035</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5002</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-2455.5,59,-2455.5</points>
<connection>
<GID>7040</GID>
<name>IN_0</name></connection>
<intersection>53 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53,-2455.5,53,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52,-2440,53,-2440</points>
<connection>
<GID>7039</GID>
<name>OUT_0</name></connection>
<intersection>53 2</intersection></hsegment></shape></wire>
<wire>
<ID>5003</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-2455.5,82,-2455.5</points>
<connection>
<GID>7042</GID>
<name>IN_0</name></connection>
<intersection>76 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76,-2455.5,76,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-2440,76,-2440</points>
<connection>
<GID>7041</GID>
<name>OUT_0</name></connection>
<intersection>76 2</intersection></hsegment></shape></wire>
<wire>
<ID>5004</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-2455.5,107,-2455.5</points>
<connection>
<GID>7045</GID>
<name>IN_0</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-2455.5,101,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-2440,101,-2440</points>
<connection>
<GID>7044</GID>
<name>OUT_0</name></connection>
<intersection>101 2</intersection></hsegment></shape></wire>
<wire>
<ID>5005</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-2455.5,130,-2455.5</points>
<connection>
<GID>7047</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-2455.5,124,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,-2440,124,-2440</points>
<connection>
<GID>7046</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>5006</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-2455.5,153,-2455.5</points>
<connection>
<GID>7050</GID>
<name>IN_0</name></connection>
<intersection>147 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>147,-2455.5,147,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>146,-2440,147,-2440</points>
<connection>
<GID>7048</GID>
<name>OUT_0</name></connection>
<intersection>147 2</intersection></hsegment></shape></wire>
<wire>
<ID>5007</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-2455.5,176,-2455.5</points>
<connection>
<GID>7052</GID>
<name>IN_0</name></connection>
<intersection>170 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>170,-2455.5,170,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169,-2440,170,-2440</points>
<connection>
<GID>7051</GID>
<name>OUT_0</name></connection>
<intersection>170 2</intersection></hsegment></shape></wire>
<wire>
<ID>5008</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2455.5,201,-2455.5</points>
<connection>
<GID>7054</GID>
<name>IN_0</name></connection>
<intersection>195 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195,-2455.5,195,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>194,-2440,195,-2440</points>
<connection>
<GID>7053</GID>
<name>OUT_0</name></connection>
<intersection>195 2</intersection></hsegment></shape></wire>
<wire>
<ID>5009</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,-2455.5,224,-2455.5</points>
<connection>
<GID>7056</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-2455.5,218,-2440</points>
<intersection>-2455.5 1</intersection>
<intersection>-2440 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-2440,218,-2440</points>
<connection>
<GID>7055</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>5010</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-2443,211,-2443</points>
<connection>
<GID>7036</GID>
<name>OUT</name></connection>
<connection>
<GID>7039</GID>
<name>clock</name></connection>
<connection>
<GID>7041</GID>
<name>clock</name></connection>
<connection>
<GID>7044</GID>
<name>clock</name></connection>
<connection>
<GID>7046</GID>
<name>clock</name></connection>
<connection>
<GID>7048</GID>
<name>clock</name></connection>
<connection>
<GID>7051</GID>
<name>clock</name></connection>
<connection>
<GID>7053</GID>
<name>clock</name></connection>
<connection>
<GID>7055</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5011</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-2452.5,222,-2452.5</points>
<connection>
<GID>7037</GID>
<name>OUT</name></connection>
<connection>
<GID>7040</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7042</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7045</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7047</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7050</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7052</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7054</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7056</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-2521.5,40.5,-2356.5</points>
<connection>
<GID>7084</GID>
<name>N_in1</name></connection>
<connection>
<GID>7057</GID>
<name>N_in0</name></connection>
<intersection>-2496 12</intersection>
<intersection>-2477.5 11</intersection>
<intersection>-2458.5 10</intersection>
<intersection>-2440 9</intersection>
<intersection>-2418 8</intersection>
<intersection>-2399.5 7</intersection>
<intersection>-2380.5 6</intersection>
<intersection>-2362 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-2362,46,-2362</points>
<connection>
<GID>6873</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40.5,-2380.5,46,-2380.5</points>
<connection>
<GID>7200</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>40.5,-2399.5,46,-2399.5</points>
<connection>
<GID>7164</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>40.5,-2418,46,-2418</points>
<connection>
<GID>7086</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>40.5,-2440,46,-2440</points>
<connection>
<GID>7039</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>40.5,-2458.5,46,-2458.5</points>
<connection>
<GID>6915</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>40.5,-2477.5,46,-2477.5</points>
<connection>
<GID>7009</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>40.5,-2496,46,-2496</points>
<connection>
<GID>6909</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-2521,63.5,-2356</points>
<connection>
<GID>7088</GID>
<name>N_in1</name></connection>
<connection>
<GID>7058</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 4</intersection>
<intersection>-2486 5</intersection>
<intersection>-2467 6</intersection>
<intersection>-2448.5 7</intersection>
<intersection>-2426.5 8</intersection>
<intersection>-2408 9</intersection>
<intersection>-2389 10</intersection>
<intersection>-2370.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>59,-2504.5,63.5,-2504.5</points>
<intersection>59 12</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>59,-2486,63.5,-2486</points>
<intersection>59 14</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59,-2467,63.5,-2467</points>
<intersection>59 13</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>59,-2448.5,63.5,-2448.5</points>
<intersection>59 15</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>59,-2426.5,63.5,-2426.5</points>
<intersection>59 18</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>59,-2408,63.5,-2408</points>
<intersection>59 19</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>59,-2389,63.5,-2389</points>
<intersection>59 20</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>59,-2370.5,63.5,-2370.5</points>
<intersection>59 21</intersection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>59,-2506,59,-2504.5</points>
<connection>
<GID>6912</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>59,-2468.5,59,-2467</points>
<connection>
<GID>6920</GID>
<name>OUT_0</name></connection>
<intersection>-2467 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>59,-2487.5,59,-2486</points>
<connection>
<GID>7010</GID>
<name>OUT_0</name></connection>
<intersection>-2486 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>59,-2450,59,-2448.5</points>
<connection>
<GID>7040</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>59,-2428,59,-2426.5</points>
<connection>
<GID>7098</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>59,-2409.5,59,-2408</points>
<connection>
<GID>7166</GID>
<name>OUT_0</name></connection>
<intersection>-2408 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>59,-2390.5,59,-2389</points>
<connection>
<GID>7202</GID>
<name>OUT_0</name></connection>
<intersection>-2389 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>59,-2372,59,-2370.5</points>
<connection>
<GID>6875</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-2521,66.5,-2356.5</points>
<connection>
<GID>7090</GID>
<name>N_in1</name></connection>
<connection>
<GID>7059</GID>
<name>N_in0</name></connection>
<intersection>-2496 10</intersection>
<intersection>-2477.5 9</intersection>
<intersection>-2458.5 8</intersection>
<intersection>-2440 7</intersection>
<intersection>-2418 6</intersection>
<intersection>-2399.5 5</intersection>
<intersection>-2380.5 4</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>66.5,-2362,69,-2362</points>
<connection>
<GID>6877</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-2380.5,69,-2380.5</points>
<connection>
<GID>7204</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66.5,-2399.5,69,-2399.5</points>
<connection>
<GID>7168</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>66.5,-2418,69,-2418</points>
<connection>
<GID>7122</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66.5,-2440,69,-2440</points>
<connection>
<GID>7041</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-2458.5,69,-2458.5</points>
<connection>
<GID>6925</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66.5,-2477.5,69,-2477.5</points>
<connection>
<GID>7011</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>66.5,-2496,69,-2496</points>
<connection>
<GID>6914</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-2521,86,-2356</points>
<connection>
<GID>7092</GID>
<name>N_in1</name></connection>
<connection>
<GID>7060</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 6</intersection>
<intersection>-2486 7</intersection>
<intersection>-2467 8</intersection>
<intersection>-2448.5 9</intersection>
<intersection>-2426.5 10</intersection>
<intersection>-2408 11</intersection>
<intersection>-2389 12</intersection>
<intersection>-2370.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>82,-2504.5,86,-2504.5</points>
<intersection>82 14</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82,-2486,86,-2486</points>
<intersection>82 16</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>82,-2467,86,-2467</points>
<intersection>82 15</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82,-2448.5,86,-2448.5</points>
<intersection>82 17</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>82,-2426.5,86,-2426.5</points>
<intersection>82 20</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>82,-2408,86,-2408</points>
<intersection>82 21</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>82,-2389,86,-2389</points>
<intersection>82 22</intersection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>82,-2370.5,86,-2370.5</points>
<intersection>82 23</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>82,-2506,82,-2504.5</points>
<connection>
<GID>6917</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>82,-2468.5,82,-2467</points>
<connection>
<GID>6930</GID>
<name>OUT_0</name></connection>
<intersection>-2467 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>82,-2487.5,82,-2486</points>
<connection>
<GID>7012</GID>
<name>OUT_0</name></connection>
<intersection>-2486 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>82,-2450,82,-2448.5</points>
<connection>
<GID>7042</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>82,-2428,82,-2426.5</points>
<connection>
<GID>7124</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>82,-2409.5,82,-2408</points>
<connection>
<GID>7170</GID>
<name>OUT_0</name></connection>
<intersection>-2408 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>82,-2390.5,82,-2389</points>
<connection>
<GID>7206</GID>
<name>OUT_0</name></connection>
<intersection>-2389 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>82,-2372,82,-2370.5</points>
<connection>
<GID>6879</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-2521,89.5,-2356</points>
<connection>
<GID>7094</GID>
<name>N_in1</name></connection>
<connection>
<GID>7061</GID>
<name>N_in0</name></connection>
<intersection>-2496 13</intersection>
<intersection>-2477.5 12</intersection>
<intersection>-2458.5 11</intersection>
<intersection>-2440 10</intersection>
<intersection>-2418 9</intersection>
<intersection>-2399.5 8</intersection>
<intersection>-2380.5 7</intersection>
<intersection>-2362 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-2362,94,-2362</points>
<connection>
<GID>6881</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-2380.5,94,-2380.5</points>
<connection>
<GID>7208</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89.5,-2399.5,94,-2399.5</points>
<connection>
<GID>7172</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-2418,94,-2418</points>
<connection>
<GID>7128</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>89.5,-2440,94,-2440</points>
<connection>
<GID>7044</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89.5,-2458.5,94,-2458.5</points>
<connection>
<GID>6935</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>89.5,-2477.5,94,-2477.5</points>
<connection>
<GID>7013</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>89.5,-2496,94,-2496</points>
<connection>
<GID>6919</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-2521,110.5,-2356.5</points>
<connection>
<GID>7096</GID>
<name>N_in1</name></connection>
<connection>
<GID>7062</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 6</intersection>
<intersection>-2486 7</intersection>
<intersection>-2467 8</intersection>
<intersection>-2448.5 9</intersection>
<intersection>-2426.5 10</intersection>
<intersection>-2408 11</intersection>
<intersection>-2389 12</intersection>
<intersection>-2370.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>107,-2504.5,110.5,-2504.5</points>
<intersection>107 14</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>107,-2486,110.5,-2486</points>
<intersection>107 16</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>107,-2467,110.5,-2467</points>
<intersection>107 15</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>107,-2448.5,110.5,-2448.5</points>
<intersection>107 17</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>107,-2426.5,110.5,-2426.5</points>
<intersection>107 20</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>107,-2408,110.5,-2408</points>
<intersection>107 21</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>107,-2389,110.5,-2389</points>
<intersection>107 22</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>107,-2370.5,110.5,-2370.5</points>
<intersection>107 23</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>107,-2506,107,-2504.5</points>
<connection>
<GID>6922</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>107,-2468.5,107,-2467</points>
<connection>
<GID>6939</GID>
<name>OUT_0</name></connection>
<intersection>-2467 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>107,-2487.5,107,-2486</points>
<connection>
<GID>7014</GID>
<name>OUT_0</name></connection>
<intersection>-2486 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>107,-2450,107,-2448.5</points>
<connection>
<GID>7045</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>107,-2428,107,-2426.5</points>
<connection>
<GID>7132</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>107,-2409.5,107,-2408</points>
<connection>
<GID>7174</GID>
<name>OUT_0</name></connection>
<intersection>-2408 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>107,-2390.5,107,-2389</points>
<connection>
<GID>7210</GID>
<name>OUT_0</name></connection>
<intersection>-2389 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>107,-2372,107,-2370.5</points>
<connection>
<GID>6883</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2521,114.5,-2356</points>
<connection>
<GID>7100</GID>
<name>N_in1</name></connection>
<connection>
<GID>7063</GID>
<name>N_in0</name></connection>
<intersection>-2496 13</intersection>
<intersection>-2477.5 12</intersection>
<intersection>-2458.5 11</intersection>
<intersection>-2440 10</intersection>
<intersection>-2418 9</intersection>
<intersection>-2399.5 8</intersection>
<intersection>-2380.5 7</intersection>
<intersection>-2362 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>114.5,-2362,117,-2362</points>
<connection>
<GID>6885</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-2380.5,117,-2380.5</points>
<connection>
<GID>7212</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-2399.5,117,-2399.5</points>
<connection>
<GID>7176</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114.5,-2418,117,-2418</points>
<connection>
<GID>7136</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114.5,-2440,117,-2440</points>
<connection>
<GID>7046</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>114.5,-2458.5,117,-2458.5</points>
<connection>
<GID>6942</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>114.5,-2477.5,117,-2477.5</points>
<connection>
<GID>7015</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>114.5,-2496,117,-2496</points>
<connection>
<GID>6924</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-2521,133,-2356</points>
<connection>
<GID>7102</GID>
<name>N_in1</name></connection>
<connection>
<GID>7064</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 6</intersection>
<intersection>-2486 7</intersection>
<intersection>-2467 8</intersection>
<intersection>-2448.5 9</intersection>
<intersection>-2426.5 10</intersection>
<intersection>-2408 11</intersection>
<intersection>-2389 12</intersection>
<intersection>-2370.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>130,-2504.5,133,-2504.5</points>
<intersection>130 14</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-2486,133,-2486</points>
<intersection>130 15</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>130,-2467,133,-2467</points>
<intersection>130 16</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>130,-2448.5,133,-2448.5</points>
<intersection>130 17</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>130,-2426.5,133,-2426.5</points>
<intersection>130 20</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>130,-2408,133,-2408</points>
<intersection>130 21</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>130,-2389,133,-2389</points>
<intersection>130 22</intersection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>130,-2370.5,133,-2370.5</points>
<intersection>130 23</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>130,-2506,130,-2504.5</points>
<connection>
<GID>6927</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>130,-2487.5,130,-2486</points>
<connection>
<GID>7016</GID>
<name>OUT_0</name></connection>
<intersection>-2486 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>130,-2468.5,130,-2467</points>
<connection>
<GID>7026</GID>
<name>OUT_0</name></connection>
<intersection>-2467 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>130,-2450,130,-2448.5</points>
<connection>
<GID>7047</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>130,-2428,130,-2426.5</points>
<connection>
<GID>7140</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>130,-2409.5,130,-2408</points>
<connection>
<GID>7178</GID>
<name>OUT_0</name></connection>
<intersection>-2408 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>130,-2390.5,130,-2389</points>
<connection>
<GID>7214</GID>
<name>OUT_0</name></connection>
<intersection>-2389 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>130,-2372,130,-2370.5</points>
<connection>
<GID>6887</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2521,137,-2356</points>
<connection>
<GID>7104</GID>
<name>N_in1</name></connection>
<connection>
<GID>7066</GID>
<name>N_in0</name></connection>
<intersection>-2496 13</intersection>
<intersection>-2477.5 12</intersection>
<intersection>-2458.5 11</intersection>
<intersection>-2440 10</intersection>
<intersection>-2418 9</intersection>
<intersection>-2399.5 8</intersection>
<intersection>-2380.5 7</intersection>
<intersection>-2362 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>137,-2362,140,-2362</points>
<connection>
<GID>6889</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137,-2380.5,140,-2380.5</points>
<connection>
<GID>7216</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-2399.5,140,-2399.5</points>
<connection>
<GID>7180</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137,-2418,140,-2418</points>
<connection>
<GID>7142</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-2440,140,-2440</points>
<connection>
<GID>7048</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>137,-2458.5,140,-2458.5</points>
<connection>
<GID>7027</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137,-2477.5,140,-2477.5</points>
<connection>
<GID>7017</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-2496,140,-2496</points>
<connection>
<GID>6929</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>5021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-2520.5,156,-2356</points>
<connection>
<GID>7106</GID>
<name>N_in1</name></connection>
<connection>
<GID>7068</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 6</intersection>
<intersection>-2486 7</intersection>
<intersection>-2467 8</intersection>
<intersection>-2448.5 9</intersection>
<intersection>-2426.5 10</intersection>
<intersection>-2408 11</intersection>
<intersection>-2389 12</intersection>
<intersection>-2370.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>153,-2504.5,156,-2504.5</points>
<intersection>153 15</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>153,-2486,156,-2486</points>
<intersection>153 16</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>153,-2467,156,-2467</points>
<intersection>153 17</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>153,-2448.5,156,-2448.5</points>
<intersection>153 18</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>153,-2426.5,156,-2426.5</points>
<intersection>153 21</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>153,-2408,156,-2408</points>
<intersection>153 22</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>153,-2389,156,-2389</points>
<intersection>153 23</intersection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>153,-2370.5,156,-2370.5</points>
<intersection>153 14</intersection>
<intersection>156 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>153,-2372,153,-2370.5</points>
<connection>
<GID>6891</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>153,-2506,153,-2504.5</points>
<connection>
<GID>6932</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>153,-2487.5,153,-2486</points>
<connection>
<GID>7018</GID>
<name>OUT_0</name></connection>
<intersection>-2486 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>153,-2468.5,153,-2467</points>
<connection>
<GID>7028</GID>
<name>OUT_0</name></connection>
<intersection>-2467 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>153,-2450,153,-2448.5</points>
<connection>
<GID>7050</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>153,-2428,153,-2426.5</points>
<connection>
<GID>7146</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>153,-2409.5,153,-2408</points>
<connection>
<GID>7182</GID>
<name>OUT_0</name></connection>
<intersection>-2408 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>153,-2390.5,153,-2389</points>
<connection>
<GID>6855</GID>
<name>OUT_0</name></connection>
<intersection>-2389 12</intersection></vsegment></shape></wire>
<wire>
<ID>5022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-2520.5,161,-2356</points>
<connection>
<GID>7108</GID>
<name>N_in1</name></connection>
<connection>
<GID>7070</GID>
<name>N_in0</name></connection>
<intersection>-2496 13</intersection>
<intersection>-2477.5 12</intersection>
<intersection>-2458.5 11</intersection>
<intersection>-2440 10</intersection>
<intersection>-2418 9</intersection>
<intersection>-2399.5 8</intersection>
<intersection>-2380.5 7</intersection>
<intersection>-2362 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>161,-2362,163,-2362</points>
<connection>
<GID>6893</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>161,-2380.5,163,-2380.5</points>
<connection>
<GID>6857</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>161,-2399.5,163,-2399.5</points>
<connection>
<GID>7184</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>161,-2418,163,-2418</points>
<connection>
<GID>7148</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>161,-2440,163,-2440</points>
<connection>
<GID>7051</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>161,-2458.5,163,-2458.5</points>
<connection>
<GID>7029</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>161,-2477.5,163,-2477.5</points>
<connection>
<GID>7019</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>161,-2496,163,-2496</points>
<connection>
<GID>6934</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>5023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-2520,179,-2356</points>
<connection>
<GID>7110</GID>
<name>N_in1</name></connection>
<connection>
<GID>7074</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 16</intersection>
<intersection>-2486 15</intersection>
<intersection>-2467 14</intersection>
<intersection>-2448.5 13</intersection>
<intersection>-2426.5 12</intersection>
<intersection>-2408 11</intersection>
<intersection>-2389 10</intersection>
<intersection>-2370.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>176,-2370.5,179,-2370.5</points>
<intersection>176 17</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>176,-2389,179,-2389</points>
<intersection>176 26</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>176,-2408,179,-2408</points>
<intersection>176 25</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>176,-2426.5,179,-2426.5</points>
<intersection>176 24</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>176,-2448.5,179,-2448.5</points>
<intersection>176 21</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>176,-2467,179,-2467</points>
<intersection>176 20</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>176,-2486,179,-2486</points>
<intersection>176 19</intersection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>176,-2504.5,179,-2504.5</points>
<intersection>176 18</intersection>
<intersection>179 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>176,-2372,176,-2370.5</points>
<connection>
<GID>6895</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>176,-2506,176,-2504.5</points>
<connection>
<GID>6937</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>176,-2487.5,176,-2486</points>
<connection>
<GID>7020</GID>
<name>OUT_0</name></connection>
<intersection>-2486 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>176,-2468.5,176,-2467</points>
<connection>
<GID>7030</GID>
<name>OUT_0</name></connection>
<intersection>-2467 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>176,-2450,176,-2448.5</points>
<connection>
<GID>7052</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>176,-2428,176,-2426.5</points>
<connection>
<GID>7150</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>176,-2409.5,176,-2408</points>
<connection>
<GID>7186</GID>
<name>OUT_0</name></connection>
<intersection>-2408 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>176,-2390.5,176,-2389</points>
<connection>
<GID>6859</GID>
<name>OUT_0</name></connection>
<intersection>-2389 10</intersection></vsegment></shape></wire>
<wire>
<ID>5024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2520,183.5,-2356</points>
<connection>
<GID>7112</GID>
<name>N_in1</name></connection>
<connection>
<GID>7072</GID>
<name>N_in0</name></connection>
<intersection>-2496 13</intersection>
<intersection>-2477.5 12</intersection>
<intersection>-2458.5 11</intersection>
<intersection>-2440 10</intersection>
<intersection>-2418 9</intersection>
<intersection>-2399.5 8</intersection>
<intersection>-2380.5 7</intersection>
<intersection>-2362 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>183.5,-2362,188,-2362</points>
<connection>
<GID>6897</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>183.5,-2380.5,188,-2380.5</points>
<connection>
<GID>6861</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>183.5,-2399.5,188,-2399.5</points>
<connection>
<GID>7188</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>183.5,-2418,188,-2418</points>
<connection>
<GID>7152</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>183.5,-2440,188,-2440</points>
<connection>
<GID>7053</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>183.5,-2458.5,188,-2458.5</points>
<connection>
<GID>7031</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>183.5,-2477.5,188,-2477.5</points>
<connection>
<GID>7021</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>183.5,-2496,188,-2496</points>
<connection>
<GID>7003</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5025</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-2519.5,204.5,-2356.5</points>
<connection>
<GID>7114</GID>
<name>N_in1</name></connection>
<connection>
<GID>7076</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 6</intersection>
<intersection>-2486 7</intersection>
<intersection>-2467 8</intersection>
<intersection>-2448.5 9</intersection>
<intersection>-2426.5 10</intersection>
<intersection>-2408 11</intersection>
<intersection>-2389 12</intersection>
<intersection>-2370.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>201,-2504.5,204.5,-2504.5</points>
<intersection>201 15</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>201,-2486,204.5,-2486</points>
<intersection>201 16</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>201,-2467,204.5,-2467</points>
<intersection>201 17</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>201,-2448.5,204.5,-2448.5</points>
<intersection>201 18</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>201,-2426.5,204.5,-2426.5</points>
<intersection>201 21</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>201,-2408,204.5,-2408</points>
<intersection>201 22</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>201,-2389,204.5,-2389</points>
<intersection>201 23</intersection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>201,-2370.5,204.5,-2370.5</points>
<intersection>201 14</intersection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>201,-2372,201,-2370.5</points>
<connection>
<GID>6899</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>201,-2506,201,-2504.5</points>
<connection>
<GID>7004</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>201,-2487.5,201,-2486</points>
<connection>
<GID>7022</GID>
<name>OUT_0</name></connection>
<intersection>-2486 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>201,-2468.5,201,-2467</points>
<connection>
<GID>7032</GID>
<name>OUT_0</name></connection>
<intersection>-2467 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>201,-2450,201,-2448.5</points>
<connection>
<GID>7054</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>201,-2428,201,-2426.5</points>
<connection>
<GID>7154</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>201,-2409.5,201,-2408</points>
<connection>
<GID>7190</GID>
<name>OUT_0</name></connection>
<intersection>-2408 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>201,-2390.5,201,-2389</points>
<connection>
<GID>6863</GID>
<name>OUT_0</name></connection>
<intersection>-2389 12</intersection></vsegment></shape></wire>
<wire>
<ID>5026</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-2519.5,208,-2356.5</points>
<connection>
<GID>7118</GID>
<name>N_in0</name></connection>
<connection>
<GID>7116</GID>
<name>N_in1</name></connection>
<intersection>-2496 11</intersection>
<intersection>-2477.5 10</intersection>
<intersection>-2458.5 9</intersection>
<intersection>-2440 7</intersection>
<intersection>-2418 6</intersection>
<intersection>-2399.5 5</intersection>
<intersection>-2380.5 4</intersection>
<intersection>-2362 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>208,-2362,211,-2362</points>
<connection>
<GID>6901</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>208,-2380.5,211,-2380.5</points>
<connection>
<GID>6865</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>208,-2399.5,211,-2399.5</points>
<connection>
<GID>7192</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>208,-2418,211,-2418</points>
<connection>
<GID>7156</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>208,-2440,211,-2440</points>
<connection>
<GID>7055</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>208,-2458.5,211,-2458.5</points>
<connection>
<GID>7034</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>208,-2477.5,211,-2477.5</points>
<connection>
<GID>7023</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>208,-2496,211,-2496</points>
<connection>
<GID>7005</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>5027</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-2519.5,229,-2357.5</points>
<connection>
<GID>7120</GID>
<name>N_in1</name></connection>
<connection>
<GID>7078</GID>
<name>N_in0</name></connection>
<intersection>-2504.5 11</intersection>
<intersection>-2486 10</intersection>
<intersection>-2467 9</intersection>
<intersection>-2448.5 8</intersection>
<intersection>-2426.5 7</intersection>
<intersection>-2408 6</intersection>
<intersection>-2389 5</intersection>
<intersection>-2370.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>224,-2370.5,229,-2370.5</points>
<intersection>224 12</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>224,-2389,229,-2389</points>
<intersection>224 21</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>224,-2408,229,-2408</points>
<intersection>224 20</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>224,-2426.5,229,-2426.5</points>
<intersection>224 19</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>224,-2448.5,229,-2448.5</points>
<intersection>224 16</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>224,-2467,229,-2467</points>
<intersection>224 15</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>224,-2486,229,-2486</points>
<intersection>224 14</intersection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>224,-2504.5,229,-2504.5</points>
<intersection>224 13</intersection>
<intersection>229 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>224,-2372,224,-2370.5</points>
<connection>
<GID>6903</GID>
<name>OUT_0</name></connection>
<intersection>-2370.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>224,-2506,224,-2504.5</points>
<connection>
<GID>7006</GID>
<name>OUT_0</name></connection>
<intersection>-2504.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>224,-2487.5,224,-2486</points>
<connection>
<GID>7024</GID>
<name>OUT_0</name></connection>
<intersection>-2486 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>224,-2468.5,224,-2467</points>
<connection>
<GID>7035</GID>
<name>OUT_0</name></connection>
<intersection>-2467 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>224,-2450,224,-2448.5</points>
<connection>
<GID>7056</GID>
<name>OUT_0</name></connection>
<intersection>-2448.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>224,-2428,224,-2426.5</points>
<connection>
<GID>7158</GID>
<name>OUT_0</name></connection>
<intersection>-2426.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>224,-2409.5,224,-2408</points>
<connection>
<GID>7194</GID>
<name>OUT_0</name></connection>
<intersection>-2408 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>224,-2390.5,224,-2389</points>
<connection>
<GID>6867</GID>
<name>OUT_0</name></connection>
<intersection>-2389 5</intersection></vsegment></shape></wire>
<wire>
<ID>5028</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-121,-2364,18.5,-2364</points>
<connection>
<GID>6869</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-2373.5,-121,-2348</points>
<intersection>-2373.5 4</intersection>
<intersection>-2364 2</intersection>
<intersection>-2348 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-2373.5,30,-2373.5</points>
<connection>
<GID>6871</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2348,-121,-2348</points>
<connection>
<GID>7002</GID>
<name>OUT_7</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>5029</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-122,-2382.5,18.5,-2382.5</points>
<connection>
<GID>7196</GID>
<name>IN_0</name></connection>
<intersection>-122 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-122,-2392,-122,-2349</points>
<intersection>-2392 5</intersection>
<intersection>-2382.5 2</intersection>
<intersection>-2349 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-122,-2392,30,-2392</points>
<connection>
<GID>7198</GID>
<name>IN_0</name></connection>
<intersection>-122 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2349,-122,-2349</points>
<connection>
<GID>7002</GID>
<name>OUT_6</name></connection>
<intersection>-122 4</intersection></hsegment></shape></wire>
<wire>
<ID>5030</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-123,-2401.5,18.5,-2401.5</points>
<connection>
<GID>7160</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-2411,-123,-2350</points>
<intersection>-2411 4</intersection>
<intersection>-2401.5 2</intersection>
<intersection>-2350 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-2411,30,-2411</points>
<connection>
<GID>7162</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2350,-123,-2350</points>
<connection>
<GID>7002</GID>
<name>OUT_5</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>5031</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-124,-2420,18.5,-2420</points>
<connection>
<GID>7080</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-2429.5,-124,-2351</points>
<intersection>-2429.5 4</intersection>
<intersection>-2420 2</intersection>
<intersection>-2351 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-2429.5,30,-2429.5</points>
<connection>
<GID>7082</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2351,-124,-2351</points>
<connection>
<GID>7002</GID>
<name>OUT_4</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>5032</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125,-2442,18.5,-2442</points>
<connection>
<GID>7036</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-125,-2451.5,-125,-2352</points>
<intersection>-2451.5 4</intersection>
<intersection>-2442 1</intersection>
<intersection>-2352 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-125,-2451.5,29.5,-2451.5</points>
<connection>
<GID>7037</GID>
<name>IN_0</name></connection>
<intersection>-125 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2352,-125,-2352</points>
<connection>
<GID>7002</GID>
<name>OUT_3</name></connection>
<intersection>-125 3</intersection></hsegment></shape></wire>
<wire>
<ID>5033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,-2460.5,18.5,-2460.5</points>
<connection>
<GID>7025</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-2470,-126,-2353</points>
<intersection>-2470 4</intersection>
<intersection>-2460.5 1</intersection>
<intersection>-2353 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-2470,29.5,-2470</points>
<connection>
<GID>6910</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2353,-126,-2353</points>
<connection>
<GID>7002</GID>
<name>OUT_2</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>5034</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127,-2479.5,18.5,-2479.5</points>
<connection>
<GID>7007</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-127,-2489,-127,-2354</points>
<intersection>-2489 4</intersection>
<intersection>-2479.5 1</intersection>
<intersection>-2354 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-127,-2489,29.5,-2489</points>
<connection>
<GID>7008</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-2354,-127,-2354</points>
<connection>
<GID>7002</GID>
<name>OUT_1</name></connection>
<intersection>-127 3</intersection></hsegment></shape></wire>
<wire>
<ID>5035</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-128,-2498,18.5,-2498</points>
<connection>
<GID>6905</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-2507.5,-128,-2355</points>
<connection>
<GID>7002</GID>
<name>OUT_0</name></connection>
<intersection>-2507.5 4</intersection>
<intersection>-2498 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-2507.5,29.5,-2507.5</points>
<connection>
<GID>6907</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>5036</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-2521.5,17.5,-2356.5</points>
<connection>
<GID>7138</GID>
<name>N_in1</name></connection>
<connection>
<GID>7130</GID>
<name>N_in0</name></connection>
<intersection>-2500 10</intersection>
<intersection>-2481.5 9</intersection>
<intersection>-2462.5 8</intersection>
<intersection>-2444 7</intersection>
<intersection>-2422 6</intersection>
<intersection>-2403.5 5</intersection>
<intersection>-2384.5 4</intersection>
<intersection>-2366 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-2366,18.5,-2366</points>
<connection>
<GID>6869</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-2384.5,18.5,-2384.5</points>
<connection>
<GID>7196</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>17.5,-2403.5,18.5,-2403.5</points>
<connection>
<GID>7160</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>17.5,-2422,18.5,-2422</points>
<connection>
<GID>7080</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>17.5,-2444,18.5,-2444</points>
<connection>
<GID>7036</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>17.5,-2462.5,18.5,-2462.5</points>
<connection>
<GID>7025</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>17.5,-2481.5,18.5,-2481.5</points>
<connection>
<GID>7007</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>17.5,-2500,18.5,-2500</points>
<connection>
<GID>6905</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5037</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-2521.5,27.5,-2356.5</points>
<connection>
<GID>7134</GID>
<name>N_in1</name></connection>
<connection>
<GID>7126</GID>
<name>N_in0</name></connection>
<intersection>-2509.5 3</intersection>
<intersection>-2491 5</intersection>
<intersection>-2472 7</intersection>
<intersection>-2453.5 9</intersection>
<intersection>-2431.5 11</intersection>
<intersection>-2413 13</intersection>
<intersection>-2394 15</intersection>
<intersection>-2375.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-2509.5,29.5,-2509.5</points>
<connection>
<GID>6907</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-2491,29.5,-2491</points>
<connection>
<GID>7008</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-2472,29.5,-2472</points>
<connection>
<GID>6910</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>27.5,-2453.5,29.5,-2453.5</points>
<connection>
<GID>7037</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>27.5,-2431.5,30,-2431.5</points>
<connection>
<GID>7082</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>27.5,-2413,30,-2413</points>
<connection>
<GID>7162</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>27.5,-2394,30,-2394</points>
<connection>
<GID>7198</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>27.5,-2375.5,30,-2375.5</points>
<connection>
<GID>6871</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5038</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-2354.5,17.5,-2348</points>
<connection>
<GID>7130</GID>
<name>N_in1</name></connection>
<connection>
<GID>7000</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-2354.5,27.5,-2348</points>
<connection>
<GID>7126</GID>
<name>N_in1</name></connection>
<connection>
<GID>6999</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5040</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-2354.5,40.5,-2348</points>
<connection>
<GID>7057</GID>
<name>N_in1</name></connection>
<connection>
<GID>6980</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-2354,63.5,-2347.5</points>
<connection>
<GID>7058</GID>
<name>N_in1</name></connection>
<connection>
<GID>6981</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-2354.5,66.5,-2347.5</points>
<connection>
<GID>7059</GID>
<name>N_in1</name></connection>
<connection>
<GID>6982</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-2354,86,-2347.5</points>
<connection>
<GID>7060</GID>
<name>N_in1</name></connection>
<connection>
<GID>6983</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5044</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-2354,89.5,-2347.5</points>
<connection>
<GID>7061</GID>
<name>N_in1</name></connection>
<connection>
<GID>6984</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5045</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-2354.5,110.5,-2347.5</points>
<connection>
<GID>7062</GID>
<name>N_in1</name></connection>
<connection>
<GID>6985</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5046</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2354,114.5,-2347.5</points>
<connection>
<GID>7063</GID>
<name>N_in1</name></connection>
<connection>
<GID>6986</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-2354,133,-2347.5</points>
<connection>
<GID>7064</GID>
<name>N_in1</name></connection>
<connection>
<GID>6987</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5048</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2354,137,-2347.5</points>
<connection>
<GID>7066</GID>
<name>N_in1</name></connection>
<connection>
<GID>6988</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-2354,156,-2347</points>
<connection>
<GID>7068</GID>
<name>N_in1</name></connection>
<connection>
<GID>6989</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-2354,161,-2347</points>
<connection>
<GID>7070</GID>
<name>N_in1</name></connection>
<connection>
<GID>6990</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-2354,179,-2346.5</points>
<connection>
<GID>7074</GID>
<name>N_in1</name></connection>
<connection>
<GID>6991</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2354,183.5,-2346.5</points>
<connection>
<GID>7072</GID>
<name>N_in1</name></connection>
<connection>
<GID>6992</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5053</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-2354.5,204.5,-2346</points>
<connection>
<GID>7076</GID>
<name>N_in1</name></connection>
<connection>
<GID>6993</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5054</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-2354.5,208,-2346</points>
<connection>
<GID>7118</GID>
<name>N_in1</name></connection>
<connection>
<GID>6994</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-2355.5,229,-2346</points>
<connection>
<GID>7078</GID>
<name>N_in1</name></connection>
<connection>
<GID>6996</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5056</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2648,63,-2648</points>
<connection>
<GID>7414</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2648,57,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2632.5,57,-2632.5</points>
<connection>
<GID>7408</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2648,86,-2648</points>
<connection>
<GID>7432</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2648,80,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2632.5,80,-2632.5</points>
<connection>
<GID>7430</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5058</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2648,111,-2648</points>
<connection>
<GID>7436</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2648,105,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2632.5,105,-2632.5</points>
<connection>
<GID>7434</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5059</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2648,134,-2648</points>
<connection>
<GID>7440</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2648,128,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2632.5,128,-2632.5</points>
<connection>
<GID>7438</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2648,157,-2648</points>
<connection>
<GID>7444</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2648,151,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2632.5,151,-2632.5</points>
<connection>
<GID>7442</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2648,180,-2648</points>
<connection>
<GID>7448</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2648,174,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2632.5,174,-2632.5</points>
<connection>
<GID>7446</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2648,205,-2648</points>
<connection>
<GID>7452</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2648,199,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2632.5,199,-2632.5</points>
<connection>
<GID>7450</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2648,228,-2648</points>
<connection>
<GID>7456</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2648,222,-2632.5</points>
<intersection>-2648 1</intersection>
<intersection>-2632.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2632.5,222,-2632.5</points>
<connection>
<GID>7454</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2635.5,215,-2635.5</points>
<connection>
<GID>7454</GID>
<name>clock</name></connection>
<connection>
<GID>7450</GID>
<name>clock</name></connection>
<connection>
<GID>7446</GID>
<name>clock</name></connection>
<connection>
<GID>7442</GID>
<name>clock</name></connection>
<connection>
<GID>7438</GID>
<name>clock</name></connection>
<connection>
<GID>7434</GID>
<name>clock</name></connection>
<connection>
<GID>7430</GID>
<name>clock</name></connection>
<connection>
<GID>7408</GID>
<name>clock</name></connection>
<connection>
<GID>7398</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2645,226,-2645</points>
<connection>
<GID>7456</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7452</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7448</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7444</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7440</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7436</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7432</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7414</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7403</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2629.5,63,-2629.5</points>
<connection>
<GID>7464</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2629.5,57,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2614,57,-2614</points>
<connection>
<GID>7462</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2629.5,86,-2629.5</points>
<connection>
<GID>7468</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2629.5,80,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2614,80,-2614</points>
<connection>
<GID>7466</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2629.5,111,-2629.5</points>
<connection>
<GID>7472</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2629.5,105,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2614,105,-2614</points>
<connection>
<GID>7470</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2629.5,134,-2629.5</points>
<connection>
<GID>7476</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2629.5,128,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2614,128,-2614</points>
<connection>
<GID>7474</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5070</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2629.5,157,-2629.5</points>
<connection>
<GID>7480</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2629.5,151,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2614,151,-2614</points>
<connection>
<GID>7478</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5071</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2629.5,180,-2629.5</points>
<connection>
<GID>7484</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2629.5,174,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2614,174,-2614</points>
<connection>
<GID>7482</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2629.5,205,-2629.5</points>
<connection>
<GID>7488</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2629.5,199,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2614,199,-2614</points>
<connection>
<GID>7486</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2629.5,228,-2629.5</points>
<connection>
<GID>7492</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2629.5,222,-2614</points>
<intersection>-2629.5 1</intersection>
<intersection>-2614 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2614,222,-2614</points>
<connection>
<GID>7490</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5074</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2617,215,-2617</points>
<connection>
<GID>7490</GID>
<name>clock</name></connection>
<connection>
<GID>7486</GID>
<name>clock</name></connection>
<connection>
<GID>7482</GID>
<name>clock</name></connection>
<connection>
<GID>7478</GID>
<name>clock</name></connection>
<connection>
<GID>7474</GID>
<name>clock</name></connection>
<connection>
<GID>7470</GID>
<name>clock</name></connection>
<connection>
<GID>7466</GID>
<name>clock</name></connection>
<connection>
<GID>7462</GID>
<name>clock</name></connection>
<connection>
<GID>7458</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5075</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2626.5,226,-2626.5</points>
<connection>
<GID>7492</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7488</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7484</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7480</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7476</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7472</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7468</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7464</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7460</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2610.5,63,-2610.5</points>
<connection>
<GID>7500</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2610.5,57,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2595,57,-2595</points>
<connection>
<GID>7498</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2610.5,86,-2610.5</points>
<connection>
<GID>7504</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2610.5,80,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2595,80,-2595</points>
<connection>
<GID>7502</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5078</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2610.5,111,-2610.5</points>
<connection>
<GID>7508</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2610.5,105,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2595,105,-2595</points>
<connection>
<GID>7506</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5079</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2610.5,134,-2610.5</points>
<connection>
<GID>7512</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2610.5,128,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2595,128,-2595</points>
<connection>
<GID>7510</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2610.5,157,-2610.5</points>
<connection>
<GID>7516</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2610.5,151,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2595,151,-2595</points>
<connection>
<GID>7514</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5081</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2610.5,180,-2610.5</points>
<connection>
<GID>7520</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2610.5,174,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2595,174,-2595</points>
<connection>
<GID>7518</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2610.5,205,-2610.5</points>
<connection>
<GID>7524</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2610.5,199,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2595,199,-2595</points>
<connection>
<GID>7522</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5083</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2610.5,228,-2610.5</points>
<connection>
<GID>7528</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2610.5,222,-2595</points>
<intersection>-2610.5 1</intersection>
<intersection>-2595 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2595,222,-2595</points>
<connection>
<GID>7526</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5084</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2598,215,-2598</points>
<connection>
<GID>7526</GID>
<name>clock</name></connection>
<connection>
<GID>7522</GID>
<name>clock</name></connection>
<connection>
<GID>7518</GID>
<name>clock</name></connection>
<connection>
<GID>7514</GID>
<name>clock</name></connection>
<connection>
<GID>7510</GID>
<name>clock</name></connection>
<connection>
<GID>7506</GID>
<name>clock</name></connection>
<connection>
<GID>7502</GID>
<name>clock</name></connection>
<connection>
<GID>7498</GID>
<name>clock</name></connection>
<connection>
<GID>7494</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5085</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2607.5,226,-2607.5</points>
<connection>
<GID>7528</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7524</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7520</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7516</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7512</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7508</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7504</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7500</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7496</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5086</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2592,63,-2592</points>
<connection>
<GID>7536</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2592,57,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2576.5,57,-2576.5</points>
<connection>
<GID>7534</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5087</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2592,86,-2592</points>
<connection>
<GID>7540</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2592,80,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2576.5,80,-2576.5</points>
<connection>
<GID>7538</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5088</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2592,111,-2592</points>
<connection>
<GID>7544</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2592,105,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2576.5,105,-2576.5</points>
<connection>
<GID>7542</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2592,134,-2592</points>
<connection>
<GID>7548</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2592,128,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2576.5,128,-2576.5</points>
<connection>
<GID>7546</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5090</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2592,157,-2592</points>
<connection>
<GID>7552</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2592,151,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2576.5,151,-2576.5</points>
<connection>
<GID>7550</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5091</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2592,180,-2592</points>
<connection>
<GID>7556</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2592,174,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2576.5,174,-2576.5</points>
<connection>
<GID>7554</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5092</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2592,205,-2592</points>
<connection>
<GID>7560</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2592,199,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2576.5,199,-2576.5</points>
<connection>
<GID>7558</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5093</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2592,228,-2592</points>
<connection>
<GID>7564</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2592,222,-2576.5</points>
<intersection>-2592 1</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2576.5,222,-2576.5</points>
<connection>
<GID>7562</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5094</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2579.5,215,-2579.5</points>
<connection>
<GID>7562</GID>
<name>clock</name></connection>
<connection>
<GID>7558</GID>
<name>clock</name></connection>
<connection>
<GID>7554</GID>
<name>clock</name></connection>
<connection>
<GID>7550</GID>
<name>clock</name></connection>
<connection>
<GID>7546</GID>
<name>clock</name></connection>
<connection>
<GID>7542</GID>
<name>clock</name></connection>
<connection>
<GID>7538</GID>
<name>clock</name></connection>
<connection>
<GID>7534</GID>
<name>clock</name></connection>
<connection>
<GID>7530</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5095</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2589,226,-2589</points>
<connection>
<GID>7564</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7560</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7556</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7552</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7548</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7544</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7540</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7536</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7532</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5096</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2726,63,-2726</points>
<connection>
<GID>7572</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2726,57,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2710.5,57,-2710.5</points>
<connection>
<GID>7570</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5097</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2726,86,-2726</points>
<connection>
<GID>7576</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2726,80,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2710.5,80,-2710.5</points>
<connection>
<GID>7574</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5098</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2726,111,-2726</points>
<connection>
<GID>7580</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2726,105,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2710.5,105,-2710.5</points>
<connection>
<GID>7578</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5099</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2726,134,-2726</points>
<connection>
<GID>7221</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2726,128,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2710.5,128,-2710.5</points>
<connection>
<GID>7219</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2726,157,-2726</points>
<connection>
<GID>7225</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2726,151,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2710.5,151,-2710.5</points>
<connection>
<GID>7223</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2726,180,-2726</points>
<connection>
<GID>7229</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2726,174,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2710.5,174,-2710.5</points>
<connection>
<GID>7227</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2726,205,-2726</points>
<connection>
<GID>7233</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2726,199,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2710.5,199,-2710.5</points>
<connection>
<GID>7231</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2726,228,-2726</points>
<connection>
<GID>7237</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2726,222,-2710.5</points>
<intersection>-2726 1</intersection>
<intersection>-2710.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2710.5,222,-2710.5</points>
<connection>
<GID>7235</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2713.5,215,-2713.5</points>
<connection>
<GID>7578</GID>
<name>clock</name></connection>
<connection>
<GID>7574</GID>
<name>clock</name></connection>
<connection>
<GID>7570</GID>
<name>clock</name></connection>
<connection>
<GID>7566</GID>
<name>OUT</name></connection>
<connection>
<GID>7235</GID>
<name>clock</name></connection>
<connection>
<GID>7231</GID>
<name>clock</name></connection>
<connection>
<GID>7227</GID>
<name>clock</name></connection>
<connection>
<GID>7223</GID>
<name>clock</name></connection>
<connection>
<GID>7219</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2723,226,-2723</points>
<connection>
<GID>7580</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7576</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7572</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7568</GID>
<name>OUT</name></connection>
<connection>
<GID>7237</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7233</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7229</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7225</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7221</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2707.5,63,-2707.5</points>
<connection>
<GID>7245</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2707.5,57,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2692,57,-2692</points>
<connection>
<GID>7243</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2707.5,86,-2707.5</points>
<connection>
<GID>7249</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2707.5,80,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2692,80,-2692</points>
<connection>
<GID>7247</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2707.5,111,-2707.5</points>
<connection>
<GID>7253</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2707.5,105,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2692,105,-2692</points>
<connection>
<GID>7251</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2707.5,134,-2707.5</points>
<connection>
<GID>7257</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2707.5,128,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2692,128,-2692</points>
<connection>
<GID>7255</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2707.5,157,-2707.5</points>
<connection>
<GID>7261</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2707.5,151,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2692,151,-2692</points>
<connection>
<GID>7259</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2707.5,180,-2707.5</points>
<connection>
<GID>7265</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2707.5,174,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2692,174,-2692</points>
<connection>
<GID>7263</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2707.5,205,-2707.5</points>
<connection>
<GID>7269</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2707.5,199,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2692,199,-2692</points>
<connection>
<GID>7267</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2707.5,228,-2707.5</points>
<connection>
<GID>7273</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2707.5,222,-2692</points>
<intersection>-2707.5 1</intersection>
<intersection>-2692 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2692,222,-2692</points>
<connection>
<GID>7271</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2695,215,-2695</points>
<connection>
<GID>7271</GID>
<name>clock</name></connection>
<connection>
<GID>7267</GID>
<name>clock</name></connection>
<connection>
<GID>7263</GID>
<name>clock</name></connection>
<connection>
<GID>7259</GID>
<name>clock</name></connection>
<connection>
<GID>7255</GID>
<name>clock</name></connection>
<connection>
<GID>7251</GID>
<name>clock</name></connection>
<connection>
<GID>7247</GID>
<name>clock</name></connection>
<connection>
<GID>7243</GID>
<name>clock</name></connection>
<connection>
<GID>7239</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2704.5,226,-2704.5</points>
<connection>
<GID>7273</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7269</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7265</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7261</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7257</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7253</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7249</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7245</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7241</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2688.5,63,-2688.5</points>
<connection>
<GID>7283</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2688.5,57,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2673,57,-2673</points>
<connection>
<GID>7281</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2688.5,86,-2688.5</points>
<connection>
<GID>7288</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2688.5,80,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2673,80,-2673</points>
<connection>
<GID>7286</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2688.5,111,-2688.5</points>
<connection>
<GID>7293</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2688.5,105,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2673,105,-2673</points>
<connection>
<GID>7291</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2688.5,134,-2688.5</points>
<connection>
<GID>7298</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2688.5,128,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2673,128,-2673</points>
<connection>
<GID>7296</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2688.5,157,-2688.5</points>
<connection>
<GID>7303</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2688.5,151,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2673,151,-2673</points>
<connection>
<GID>7301</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2688.5,180,-2688.5</points>
<connection>
<GID>7306</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2688.5,174,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2673,174,-2673</points>
<connection>
<GID>7305</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2688.5,205,-2688.5</points>
<connection>
<GID>7309</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2688.5,199,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2673,199,-2673</points>
<connection>
<GID>7308</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2688.5,228,-2688.5</points>
<connection>
<GID>7311</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2688.5,222,-2673</points>
<intersection>-2688.5 1</intersection>
<intersection>-2673 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2673,222,-2673</points>
<connection>
<GID>7310</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2676,215,-2676</points>
<connection>
<GID>7310</GID>
<name>clock</name></connection>
<connection>
<GID>7308</GID>
<name>clock</name></connection>
<connection>
<GID>7305</GID>
<name>clock</name></connection>
<connection>
<GID>7301</GID>
<name>clock</name></connection>
<connection>
<GID>7296</GID>
<name>clock</name></connection>
<connection>
<GID>7291</GID>
<name>clock</name></connection>
<connection>
<GID>7286</GID>
<name>clock</name></connection>
<connection>
<GID>7281</GID>
<name>clock</name></connection>
<connection>
<GID>7276</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2685.5,226,-2685.5</points>
<connection>
<GID>7311</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7309</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7306</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7303</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7298</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7293</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7288</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7283</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7278</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2670,63,-2670</points>
<connection>
<GID>7315</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2670,57,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2654.5,57,-2654.5</points>
<connection>
<GID>7314</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2670,86,-2670</points>
<connection>
<GID>7317</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2670,80,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2654.5,80,-2654.5</points>
<connection>
<GID>7316</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2670,111,-2670</points>
<connection>
<GID>7319</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2670,105,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2654.5,105,-2654.5</points>
<connection>
<GID>7318</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2670,134,-2670</points>
<connection>
<GID>7321</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2670,128,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2654.5,128,-2654.5</points>
<connection>
<GID>7320</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2670,157,-2670</points>
<connection>
<GID>7323</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2670,151,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2654.5,151,-2654.5</points>
<connection>
<GID>7322</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2670,180,-2670</points>
<connection>
<GID>7325</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2670,174,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2654.5,174,-2654.5</points>
<connection>
<GID>7324</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2670,205,-2670</points>
<connection>
<GID>7327</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2670,199,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2654.5,199,-2654.5</points>
<connection>
<GID>7326</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2670,228,-2670</points>
<connection>
<GID>7329</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2670,222,-2654.5</points>
<intersection>-2670 1</intersection>
<intersection>-2654.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2654.5,222,-2654.5</points>
<connection>
<GID>7328</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2657.5,215,-2657.5</points>
<connection>
<GID>7328</GID>
<name>clock</name></connection>
<connection>
<GID>7326</GID>
<name>clock</name></connection>
<connection>
<GID>7324</GID>
<name>clock</name></connection>
<connection>
<GID>7322</GID>
<name>clock</name></connection>
<connection>
<GID>7320</GID>
<name>clock</name></connection>
<connection>
<GID>7318</GID>
<name>clock</name></connection>
<connection>
<GID>7316</GID>
<name>clock</name></connection>
<connection>
<GID>7314</GID>
<name>clock</name></connection>
<connection>
<GID>7312</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2667,226,-2667</points>
<connection>
<GID>7329</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7327</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7325</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7323</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7321</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7319</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7317</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7315</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7313</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-2736,44.5,-2571</points>
<connection>
<GID>7345</GID>
<name>N_in1</name></connection>
<connection>
<GID>7330</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 12</intersection>
<intersection>-2692 11</intersection>
<intersection>-2673 10</intersection>
<intersection>-2654.5 9</intersection>
<intersection>-2632.5 8</intersection>
<intersection>-2614 7</intersection>
<intersection>-2595 6</intersection>
<intersection>-2576.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-2576.5,50,-2576.5</points>
<connection>
<GID>7534</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>44.5,-2595,50,-2595</points>
<connection>
<GID>7498</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-2614,50,-2614</points>
<connection>
<GID>7462</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>44.5,-2632.5,50,-2632.5</points>
<connection>
<GID>7408</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>44.5,-2654.5,50,-2654.5</points>
<connection>
<GID>7314</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>44.5,-2673,50,-2673</points>
<connection>
<GID>7281</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>44.5,-2692,50,-2692</points>
<connection>
<GID>7243</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>44.5,-2710.5,50,-2710.5</points>
<connection>
<GID>7570</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-2735.5,67.5,-2570.5</points>
<connection>
<GID>7346</GID>
<name>N_in1</name></connection>
<connection>
<GID>7331</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 4</intersection>
<intersection>-2700 5</intersection>
<intersection>-2681 6</intersection>
<intersection>-2662.5 7</intersection>
<intersection>-2640.5 8</intersection>
<intersection>-2622 9</intersection>
<intersection>-2603 10</intersection>
<intersection>-2584.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63,-2718.5,67.5,-2718.5</points>
<intersection>63 12</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-2700,67.5,-2700</points>
<intersection>63 13</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>63,-2681,67.5,-2681</points>
<intersection>63 14</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>63,-2662.5,67.5,-2662.5</points>
<intersection>63 15</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>63,-2640.5,67.5,-2640.5</points>
<intersection>63 18</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-2622,67.5,-2622</points>
<intersection>63 19</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>63,-2603,67.5,-2603</points>
<intersection>63 20</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>63,-2584.5,67.5,-2584.5</points>
<intersection>63 21</intersection>
<intersection>67.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>63,-2720.5,63,-2718.5</points>
<connection>
<GID>7572</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>63,-2702,63,-2700</points>
<connection>
<GID>7245</GID>
<name>OUT_0</name></connection>
<intersection>-2700 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>63,-2683,63,-2681</points>
<connection>
<GID>7283</GID>
<name>OUT_0</name></connection>
<intersection>-2681 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>63,-2664.5,63,-2662.5</points>
<connection>
<GID>7315</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>63,-2642.5,63,-2640.5</points>
<connection>
<GID>7414</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>63,-2624,63,-2622</points>
<connection>
<GID>7464</GID>
<name>OUT_0</name></connection>
<intersection>-2622 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>63,-2605,63,-2603</points>
<connection>
<GID>7500</GID>
<name>OUT_0</name></connection>
<intersection>-2603 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>63,-2586.5,63,-2584.5</points>
<connection>
<GID>7536</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-2735.5,70.5,-2571</points>
<connection>
<GID>7347</GID>
<name>N_in1</name></connection>
<connection>
<GID>7332</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 10</intersection>
<intersection>-2692 9</intersection>
<intersection>-2673 8</intersection>
<intersection>-2654.5 7</intersection>
<intersection>-2632.5 6</intersection>
<intersection>-2614 5</intersection>
<intersection>-2595 4</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70.5,-2576.5,73,-2576.5</points>
<connection>
<GID>7538</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-2595,73,-2595</points>
<connection>
<GID>7502</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-2614,73,-2614</points>
<connection>
<GID>7466</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>70.5,-2632.5,73,-2632.5</points>
<connection>
<GID>7430</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>70.5,-2654.5,73,-2654.5</points>
<connection>
<GID>7316</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>70.5,-2673,73,-2673</points>
<connection>
<GID>7286</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>70.5,-2692,73,-2692</points>
<connection>
<GID>7247</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>70.5,-2710.5,73,-2710.5</points>
<connection>
<GID>7574</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-2735.5,90,-2570.5</points>
<connection>
<GID>7348</GID>
<name>N_in1</name></connection>
<connection>
<GID>7333</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 6</intersection>
<intersection>-2700 7</intersection>
<intersection>-2681 8</intersection>
<intersection>-2662.5 9</intersection>
<intersection>-2640.5 10</intersection>
<intersection>-2622 11</intersection>
<intersection>-2603 12</intersection>
<intersection>-2584.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-2718.5,90,-2718.5</points>
<intersection>86 14</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>86,-2700,90,-2700</points>
<intersection>86 15</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>86,-2681,90,-2681</points>
<intersection>86 16</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>86,-2662.5,90,-2662.5</points>
<intersection>86 17</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>86,-2640.5,90,-2640.5</points>
<intersection>86 20</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>86,-2622,90,-2622</points>
<intersection>86 21</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>86,-2603,90,-2603</points>
<intersection>86 22</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>86,-2584.5,90,-2584.5</points>
<intersection>86 23</intersection>
<intersection>90 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>86,-2720.5,86,-2718.5</points>
<connection>
<GID>7576</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>86,-2702,86,-2700</points>
<connection>
<GID>7249</GID>
<name>OUT_0</name></connection>
<intersection>-2700 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>86,-2683,86,-2681</points>
<connection>
<GID>7288</GID>
<name>OUT_0</name></connection>
<intersection>-2681 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>86,-2664.5,86,-2662.5</points>
<connection>
<GID>7317</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>86,-2642.5,86,-2640.5</points>
<connection>
<GID>7432</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>86,-2624,86,-2622</points>
<connection>
<GID>7468</GID>
<name>OUT_0</name></connection>
<intersection>-2622 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>86,-2605,86,-2603</points>
<connection>
<GID>7504</GID>
<name>OUT_0</name></connection>
<intersection>-2603 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>86,-2586.5,86,-2584.5</points>
<connection>
<GID>7540</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-2735.5,93.5,-2570.5</points>
<connection>
<GID>7349</GID>
<name>N_in1</name></connection>
<connection>
<GID>7334</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 13</intersection>
<intersection>-2692 12</intersection>
<intersection>-2673 11</intersection>
<intersection>-2654.5 10</intersection>
<intersection>-2632.5 9</intersection>
<intersection>-2614 8</intersection>
<intersection>-2595 7</intersection>
<intersection>-2576.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>93.5,-2576.5,98,-2576.5</points>
<connection>
<GID>7542</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>93.5,-2595,98,-2595</points>
<connection>
<GID>7506</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>93.5,-2614,98,-2614</points>
<connection>
<GID>7470</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-2632.5,98,-2632.5</points>
<connection>
<GID>7434</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>93.5,-2654.5,98,-2654.5</points>
<connection>
<GID>7318</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>93.5,-2673,98,-2673</points>
<connection>
<GID>7291</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>93.5,-2692,98,-2692</points>
<connection>
<GID>7251</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>93.5,-2710.5,98,-2710.5</points>
<connection>
<GID>7578</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2735.5,114.5,-2571</points>
<connection>
<GID>7350</GID>
<name>N_in1</name></connection>
<connection>
<GID>7335</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 6</intersection>
<intersection>-2700 7</intersection>
<intersection>-2681 8</intersection>
<intersection>-2662.5 9</intersection>
<intersection>-2640.5 10</intersection>
<intersection>-2622 11</intersection>
<intersection>-2603 12</intersection>
<intersection>-2584.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>111,-2718.5,114.5,-2718.5</points>
<intersection>111 14</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111,-2700,114.5,-2700</points>
<intersection>111 15</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111,-2681,114.5,-2681</points>
<intersection>111 16</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111,-2662.5,114.5,-2662.5</points>
<intersection>111 17</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,-2640.5,114.5,-2640.5</points>
<intersection>111 20</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>111,-2622,114.5,-2622</points>
<intersection>111 21</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>111,-2603,114.5,-2603</points>
<intersection>111 22</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111,-2584.5,114.5,-2584.5</points>
<intersection>111 23</intersection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>111,-2720.5,111,-2718.5</points>
<connection>
<GID>7580</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>111,-2702,111,-2700</points>
<connection>
<GID>7253</GID>
<name>OUT_0</name></connection>
<intersection>-2700 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>111,-2683,111,-2681</points>
<connection>
<GID>7293</GID>
<name>OUT_0</name></connection>
<intersection>-2681 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>111,-2664.5,111,-2662.5</points>
<connection>
<GID>7319</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>111,-2642.5,111,-2640.5</points>
<connection>
<GID>7436</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>111,-2624,111,-2622</points>
<connection>
<GID>7472</GID>
<name>OUT_0</name></connection>
<intersection>-2622 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>111,-2605,111,-2603</points>
<connection>
<GID>7508</GID>
<name>OUT_0</name></connection>
<intersection>-2603 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>111,-2586.5,111,-2584.5</points>
<connection>
<GID>7544</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-2735.5,118.5,-2570.5</points>
<connection>
<GID>7351</GID>
<name>N_in1</name></connection>
<connection>
<GID>7336</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 13</intersection>
<intersection>-2692 12</intersection>
<intersection>-2673 11</intersection>
<intersection>-2654.5 10</intersection>
<intersection>-2632.5 9</intersection>
<intersection>-2614 8</intersection>
<intersection>-2595 7</intersection>
<intersection>-2576.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>118.5,-2576.5,121,-2576.5</points>
<connection>
<GID>7546</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>118.5,-2595,121,-2595</points>
<connection>
<GID>7510</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118.5,-2614,121,-2614</points>
<connection>
<GID>7474</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>118.5,-2632.5,121,-2632.5</points>
<connection>
<GID>7438</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>118.5,-2654.5,121,-2654.5</points>
<connection>
<GID>7320</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>118.5,-2673,121,-2673</points>
<connection>
<GID>7296</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>118.5,-2692,121,-2692</points>
<connection>
<GID>7255</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>118.5,-2710.5,121,-2710.5</points>
<connection>
<GID>7219</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2735.5,137,-2570.5</points>
<connection>
<GID>7352</GID>
<name>N_in1</name></connection>
<connection>
<GID>7337</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 6</intersection>
<intersection>-2700 7</intersection>
<intersection>-2681 8</intersection>
<intersection>-2662.5 9</intersection>
<intersection>-2640.5 10</intersection>
<intersection>-2622 11</intersection>
<intersection>-2603 12</intersection>
<intersection>-2584.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>134,-2718.5,137,-2718.5</points>
<intersection>134 14</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>134,-2700,137,-2700</points>
<intersection>134 15</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>134,-2681,137,-2681</points>
<intersection>134 16</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>134,-2662.5,137,-2662.5</points>
<intersection>134 17</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>134,-2640.5,137,-2640.5</points>
<intersection>134 20</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>134,-2622,137,-2622</points>
<intersection>134 21</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>134,-2603,137,-2603</points>
<intersection>134 22</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>134,-2584.5,137,-2584.5</points>
<intersection>134 23</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>134,-2720.5,134,-2718.5</points>
<connection>
<GID>7221</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>134,-2702,134,-2700</points>
<connection>
<GID>7257</GID>
<name>OUT_0</name></connection>
<intersection>-2700 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>134,-2683,134,-2681</points>
<connection>
<GID>7298</GID>
<name>OUT_0</name></connection>
<intersection>-2681 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>134,-2664.5,134,-2662.5</points>
<connection>
<GID>7321</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>134,-2642.5,134,-2640.5</points>
<connection>
<GID>7440</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>134,-2624,134,-2622</points>
<connection>
<GID>7476</GID>
<name>OUT_0</name></connection>
<intersection>-2622 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>134,-2605,134,-2603</points>
<connection>
<GID>7512</GID>
<name>OUT_0</name></connection>
<intersection>-2603 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>134,-2586.5,134,-2584.5</points>
<connection>
<GID>7548</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-2735.5,141,-2570.5</points>
<connection>
<GID>7353</GID>
<name>N_in1</name></connection>
<connection>
<GID>7338</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 13</intersection>
<intersection>-2692 12</intersection>
<intersection>-2673 11</intersection>
<intersection>-2654.5 10</intersection>
<intersection>-2632.5 9</intersection>
<intersection>-2614 8</intersection>
<intersection>-2595 7</intersection>
<intersection>-2576.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>141,-2576.5,144,-2576.5</points>
<connection>
<GID>7550</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>141,-2595,144,-2595</points>
<connection>
<GID>7514</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>141,-2614,144,-2614</points>
<connection>
<GID>7478</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>141,-2632.5,144,-2632.5</points>
<connection>
<GID>7442</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>141,-2654.5,144,-2654.5</points>
<connection>
<GID>7322</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>141,-2673,144,-2673</points>
<connection>
<GID>7301</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>141,-2692,144,-2692</points>
<connection>
<GID>7259</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>141,-2710.5,144,-2710.5</points>
<connection>
<GID>7223</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>5145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-2735,160,-2570.5</points>
<connection>
<GID>7354</GID>
<name>N_in1</name></connection>
<connection>
<GID>7339</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 6</intersection>
<intersection>-2700 7</intersection>
<intersection>-2681 8</intersection>
<intersection>-2662.5 9</intersection>
<intersection>-2640.5 10</intersection>
<intersection>-2622 11</intersection>
<intersection>-2603 12</intersection>
<intersection>-2584.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>157,-2718.5,160,-2718.5</points>
<intersection>157 14</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>157,-2700,160,-2700</points>
<intersection>157 15</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>157,-2681,160,-2681</points>
<intersection>157 16</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,-2662.5,160,-2662.5</points>
<intersection>157 17</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>157,-2640.5,160,-2640.5</points>
<intersection>157 20</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>157,-2622,160,-2622</points>
<intersection>157 21</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>157,-2603,160,-2603</points>
<intersection>157 22</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>157,-2584.5,160,-2584.5</points>
<intersection>157 23</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>157,-2720.5,157,-2718.5</points>
<connection>
<GID>7225</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>157,-2702,157,-2700</points>
<connection>
<GID>7261</GID>
<name>OUT_0</name></connection>
<intersection>-2700 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>157,-2683,157,-2681</points>
<connection>
<GID>7303</GID>
<name>OUT_0</name></connection>
<intersection>-2681 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>157,-2664.5,157,-2662.5</points>
<connection>
<GID>7323</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>157,-2642.5,157,-2640.5</points>
<connection>
<GID>7444</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>157,-2624,157,-2622</points>
<connection>
<GID>7480</GID>
<name>OUT_0</name></connection>
<intersection>-2622 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>157,-2605,157,-2603</points>
<connection>
<GID>7516</GID>
<name>OUT_0</name></connection>
<intersection>-2603 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>157,-2586.5,157,-2584.5</points>
<connection>
<GID>7552</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-2735,165,-2570.5</points>
<connection>
<GID>7355</GID>
<name>N_in1</name></connection>
<connection>
<GID>7340</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 13</intersection>
<intersection>-2692 12</intersection>
<intersection>-2673 11</intersection>
<intersection>-2654.5 10</intersection>
<intersection>-2632.5 9</intersection>
<intersection>-2614 8</intersection>
<intersection>-2595 7</intersection>
<intersection>-2576.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>165,-2576.5,167,-2576.5</points>
<connection>
<GID>7554</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>165,-2595,167,-2595</points>
<connection>
<GID>7518</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>165,-2614,167,-2614</points>
<connection>
<GID>7482</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>165,-2632.5,167,-2632.5</points>
<connection>
<GID>7446</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>165,-2654.5,167,-2654.5</points>
<connection>
<GID>7324</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>165,-2673,167,-2673</points>
<connection>
<GID>7305</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>165,-2692,167,-2692</points>
<connection>
<GID>7263</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>165,-2710.5,167,-2710.5</points>
<connection>
<GID>7227</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>5147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-2734.5,183,-2570.5</points>
<connection>
<GID>7356</GID>
<name>N_in1</name></connection>
<connection>
<GID>7342</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 16</intersection>
<intersection>-2700 15</intersection>
<intersection>-2681 14</intersection>
<intersection>-2662.5 13</intersection>
<intersection>-2640.5 12</intersection>
<intersection>-2622 11</intersection>
<intersection>-2603 10</intersection>
<intersection>-2584.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>180,-2584.5,183,-2584.5</points>
<intersection>180 26</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>180,-2603,183,-2603</points>
<intersection>180 25</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>180,-2622,183,-2622</points>
<intersection>180 24</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>180,-2640.5,183,-2640.5</points>
<intersection>180 23</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>180,-2662.5,183,-2662.5</points>
<intersection>180 20</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>180,-2681,183,-2681</points>
<intersection>180 19</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>180,-2700,183,-2700</points>
<intersection>180 18</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>180,-2718.5,183,-2718.5</points>
<intersection>180 17</intersection>
<intersection>183 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>180,-2720.5,180,-2718.5</points>
<connection>
<GID>7229</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>180,-2702,180,-2700</points>
<connection>
<GID>7265</GID>
<name>OUT_0</name></connection>
<intersection>-2700 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>180,-2683,180,-2681</points>
<connection>
<GID>7306</GID>
<name>OUT_0</name></connection>
<intersection>-2681 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>180,-2664.5,180,-2662.5</points>
<connection>
<GID>7325</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>180,-2642.5,180,-2640.5</points>
<connection>
<GID>7448</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>180,-2624,180,-2622</points>
<connection>
<GID>7484</GID>
<name>OUT_0</name></connection>
<intersection>-2622 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>180,-2605,180,-2603</points>
<connection>
<GID>7520</GID>
<name>OUT_0</name></connection>
<intersection>-2603 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>180,-2586.5,180,-2584.5</points>
<connection>
<GID>7556</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>5148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-2734.5,187.5,-2570.5</points>
<connection>
<GID>7357</GID>
<name>N_in1</name></connection>
<connection>
<GID>7341</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 13</intersection>
<intersection>-2692 12</intersection>
<intersection>-2673 11</intersection>
<intersection>-2654.5 10</intersection>
<intersection>-2632.5 9</intersection>
<intersection>-2614 8</intersection>
<intersection>-2595 7</intersection>
<intersection>-2576.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>187.5,-2576.5,192,-2576.5</points>
<connection>
<GID>7558</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>187.5,-2595,192,-2595</points>
<connection>
<GID>7522</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187.5,-2614,192,-2614</points>
<connection>
<GID>7486</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>187.5,-2632.5,192,-2632.5</points>
<connection>
<GID>7450</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>187.5,-2654.5,192,-2654.5</points>
<connection>
<GID>7326</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>187.5,-2673,192,-2673</points>
<connection>
<GID>7308</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>187.5,-2692,192,-2692</points>
<connection>
<GID>7267</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>187.5,-2710.5,192,-2710.5</points>
<connection>
<GID>7231</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-2734,208.5,-2571</points>
<connection>
<GID>7358</GID>
<name>N_in1</name></connection>
<connection>
<GID>7343</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 6</intersection>
<intersection>-2700 7</intersection>
<intersection>-2681 8</intersection>
<intersection>-2662.5 9</intersection>
<intersection>-2640.5 10</intersection>
<intersection>-2622 11</intersection>
<intersection>-2603 12</intersection>
<intersection>-2584.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>205,-2718.5,208.5,-2718.5</points>
<intersection>205 14</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205,-2700,208.5,-2700</points>
<intersection>205 15</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>205,-2681,208.5,-2681</points>
<intersection>205 16</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>205,-2662.5,208.5,-2662.5</points>
<intersection>205 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>205,-2640.5,208.5,-2640.5</points>
<intersection>205 20</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205,-2622,208.5,-2622</points>
<intersection>205 21</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>205,-2603,208.5,-2603</points>
<intersection>205 22</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>205,-2584.5,208.5,-2584.5</points>
<intersection>205 23</intersection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>205,-2720.5,205,-2718.5</points>
<connection>
<GID>7233</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>205,-2702,205,-2700</points>
<connection>
<GID>7269</GID>
<name>OUT_0</name></connection>
<intersection>-2700 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>205,-2683,205,-2681</points>
<connection>
<GID>7309</GID>
<name>OUT_0</name></connection>
<intersection>-2681 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>205,-2664.5,205,-2662.5</points>
<connection>
<GID>7327</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>205,-2642.5,205,-2640.5</points>
<connection>
<GID>7452</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>205,-2624,205,-2622</points>
<connection>
<GID>7488</GID>
<name>OUT_0</name></connection>
<intersection>-2622 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>205,-2605,205,-2603</points>
<connection>
<GID>7524</GID>
<name>OUT_0</name></connection>
<intersection>-2603 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>205,-2586.5,205,-2584.5</points>
<connection>
<GID>7560</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-2734,212,-2571</points>
<connection>
<GID>7359</GID>
<name>N_in1</name></connection>
<connection>
<GID>7360</GID>
<name>N_in0</name></connection>
<intersection>-2710.5 11</intersection>
<intersection>-2692 10</intersection>
<intersection>-2673 9</intersection>
<intersection>-2654.5 7</intersection>
<intersection>-2632.5 6</intersection>
<intersection>-2614 5</intersection>
<intersection>-2595 4</intersection>
<intersection>-2576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-2576.5,215,-2576.5</points>
<connection>
<GID>7562</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>212,-2595,215,-2595</points>
<connection>
<GID>7526</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>212,-2614,215,-2614</points>
<connection>
<GID>7490</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>212,-2632.5,215,-2632.5</points>
<connection>
<GID>7454</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>212,-2654.5,215,-2654.5</points>
<connection>
<GID>7328</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>212,-2673,215,-2673</points>
<connection>
<GID>7310</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>212,-2692,215,-2692</points>
<connection>
<GID>7271</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>212,-2710.5,215,-2710.5</points>
<connection>
<GID>7235</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>5151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-2734,233,-2572</points>
<connection>
<GID>7361</GID>
<name>N_in1</name></connection>
<connection>
<GID>7344</GID>
<name>N_in0</name></connection>
<intersection>-2718.5 11</intersection>
<intersection>-2700 10</intersection>
<intersection>-2681 9</intersection>
<intersection>-2662.5 8</intersection>
<intersection>-2640.5 7</intersection>
<intersection>-2622 6</intersection>
<intersection>-2603 5</intersection>
<intersection>-2584.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>228,-2584.5,233,-2584.5</points>
<intersection>228 21</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-2603,233,-2603</points>
<intersection>228 20</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>228,-2622,233,-2622</points>
<intersection>228 19</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>228,-2640.5,233,-2640.5</points>
<intersection>228 18</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>228,-2662.5,233,-2662.5</points>
<intersection>228 15</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>228,-2681,233,-2681</points>
<intersection>228 14</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>228,-2700,233,-2700</points>
<intersection>228 13</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>228,-2718.5,233,-2718.5</points>
<intersection>228 12</intersection>
<intersection>233 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>228,-2720.5,228,-2718.5</points>
<connection>
<GID>7237</GID>
<name>OUT_0</name></connection>
<intersection>-2718.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>228,-2702,228,-2700</points>
<connection>
<GID>7273</GID>
<name>OUT_0</name></connection>
<intersection>-2700 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>228,-2683,228,-2681</points>
<connection>
<GID>7311</GID>
<name>OUT_0</name></connection>
<intersection>-2681 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>228,-2664.5,228,-2662.5</points>
<connection>
<GID>7329</GID>
<name>OUT_0</name></connection>
<intersection>-2662.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>228,-2642.5,228,-2640.5</points>
<connection>
<GID>7456</GID>
<name>OUT_0</name></connection>
<intersection>-2640.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>228,-2624,228,-2622</points>
<connection>
<GID>7492</GID>
<name>OUT_0</name></connection>
<intersection>-2622 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>228,-2605,228,-2603</points>
<connection>
<GID>7528</GID>
<name>OUT_0</name></connection>
<intersection>-2603 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>228,-2586.5,228,-2584.5</points>
<connection>
<GID>7564</GID>
<name>OUT_0</name></connection>
<intersection>-2584.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>5152</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-124,-2578.5,22.5,-2578.5</points>
<connection>
<GID>7530</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-2730,-124,-2578.5</points>
<connection>
<GID>7367</GID>
<name>OUT_15</name></connection>
<intersection>-2588 4</intersection>
<intersection>-2578.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-2588,34,-2588</points>
<connection>
<GID>7532</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>5153</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-123,-2597,22.5,-2597</points>
<connection>
<GID>7494</GID>
<name>IN_0</name></connection>
<intersection>-123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-123,-2731,-123,-2597</points>
<intersection>-2731 6</intersection>
<intersection>-2606.5 5</intersection>
<intersection>-2597 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-123,-2606.5,34,-2606.5</points>
<connection>
<GID>7496</GID>
<name>IN_0</name></connection>
<intersection>-123 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-2731,-123,-2731</points>
<connection>
<GID>7367</GID>
<name>OUT_14</name></connection>
<intersection>-123 4</intersection></hsegment></shape></wire>
<wire>
<ID>5154</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-122,-2616,22.5,-2616</points>
<connection>
<GID>7458</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-2732,-122,-2616</points>
<intersection>-2732 6</intersection>
<intersection>-2625.5 4</intersection>
<intersection>-2616 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-2625.5,34,-2625.5</points>
<connection>
<GID>7460</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-2732,-122,-2732</points>
<connection>
<GID>7367</GID>
<name>OUT_13</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>5155</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-121,-2634.5,22.5,-2634.5</points>
<connection>
<GID>7398</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-2733,-121,-2634.5</points>
<intersection>-2733 5</intersection>
<intersection>-2644 4</intersection>
<intersection>-2634.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-2644,34,-2644</points>
<connection>
<GID>7403</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2733,-121,-2733</points>
<connection>
<GID>7367</GID>
<name>OUT_12</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>5156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-2656.5,22.5,-2656.5</points>
<connection>
<GID>7312</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-2734,-120,-2656.5</points>
<intersection>-2734 6</intersection>
<intersection>-2666 4</intersection>
<intersection>-2656.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-120,-2666,33.5,-2666</points>
<connection>
<GID>7313</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-2734,-120,-2734</points>
<connection>
<GID>7367</GID>
<name>OUT_11</name></connection>
<intersection>-120 3</intersection></hsegment></shape></wire>
<wire>
<ID>5157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,-2675,22.5,-2675</points>
<connection>
<GID>7276</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-2735,-119,-2675</points>
<intersection>-2735 5</intersection>
<intersection>-2684.5 4</intersection>
<intersection>-2675 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-2684.5,33.5,-2684.5</points>
<connection>
<GID>7278</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2735,-119,-2735</points>
<connection>
<GID>7367</GID>
<name>OUT_10</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>5158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118,-2694,22.5,-2694</points>
<connection>
<GID>7239</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-118,-2736,-118,-2694</points>
<intersection>-2736 5</intersection>
<intersection>-2703.5 4</intersection>
<intersection>-2694 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-118,-2703.5,33.5,-2703.5</points>
<connection>
<GID>7241</GID>
<name>IN_0</name></connection>
<intersection>-118 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2736,-118,-2736</points>
<connection>
<GID>7367</GID>
<name>OUT_9</name></connection>
<intersection>-118 3</intersection></hsegment></shape></wire>
<wire>
<ID>5159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-117,-2712.5,22.5,-2712.5</points>
<connection>
<GID>7566</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-2737,-117,-2712.5</points>
<intersection>-2737 5</intersection>
<intersection>-2722 4</intersection>
<intersection>-2712.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-2722,33.5,-2722</points>
<connection>
<GID>7568</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2737,-117,-2737</points>
<connection>
<GID>7367</GID>
<name>OUT_8</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>5160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-2736,21.5,-2571</points>
<connection>
<GID>7365</GID>
<name>N_in1</name></connection>
<connection>
<GID>7363</GID>
<name>N_in0</name></connection>
<intersection>-2714.5 10</intersection>
<intersection>-2696 9</intersection>
<intersection>-2677 8</intersection>
<intersection>-2658.5 7</intersection>
<intersection>-2636.5 6</intersection>
<intersection>-2618 5</intersection>
<intersection>-2599 4</intersection>
<intersection>-2580.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-2580.5,22.5,-2580.5</points>
<connection>
<GID>7530</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-2599,22.5,-2599</points>
<connection>
<GID>7494</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>21.5,-2618,22.5,-2618</points>
<connection>
<GID>7458</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-2636.5,22.5,-2636.5</points>
<connection>
<GID>7398</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21.5,-2658.5,22.5,-2658.5</points>
<connection>
<GID>7312</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>21.5,-2677,22.5,-2677</points>
<connection>
<GID>7276</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>21.5,-2696,22.5,-2696</points>
<connection>
<GID>7239</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>21.5,-2714.5,22.5,-2714.5</points>
<connection>
<GID>7566</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-2736,31.5,-2571</points>
<connection>
<GID>7364</GID>
<name>N_in1</name></connection>
<connection>
<GID>7362</GID>
<name>N_in0</name></connection>
<intersection>-2724 3</intersection>
<intersection>-2705.5 5</intersection>
<intersection>-2686.5 7</intersection>
<intersection>-2668 9</intersection>
<intersection>-2646 11</intersection>
<intersection>-2627.5 13</intersection>
<intersection>-2608.5 15</intersection>
<intersection>-2590 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-2724,33.5,-2724</points>
<connection>
<GID>7568</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-2705.5,33.5,-2705.5</points>
<connection>
<GID>7241</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31.5,-2686.5,33.5,-2686.5</points>
<connection>
<GID>7278</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>31.5,-2668,33.5,-2668</points>
<connection>
<GID>7313</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>31.5,-2646,34,-2646</points>
<connection>
<GID>7403</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>31.5,-2627.5,34,-2627.5</points>
<connection>
<GID>7460</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>31.5,-2608.5,34,-2608.5</points>
<connection>
<GID>7496</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>31.5,-2590,34,-2590</points>
<connection>
<GID>7532</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2823.5,63,-2823.5</points>
<connection>
<GID>7463</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2823.5,57,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2808,57,-2808</points>
<connection>
<GID>7451</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2823.5,86,-2823.5</points>
<connection>
<GID>7489</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2823.5,80,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2808,80,-2808</points>
<connection>
<GID>7487</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2823.5,111,-2823.5</points>
<connection>
<GID>7497</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2823.5,105,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2808,105,-2808</points>
<connection>
<GID>7493</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2823.5,134,-2823.5</points>
<connection>
<GID>7505</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2823.5,128,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2808,128,-2808</points>
<connection>
<GID>7501</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2823.5,157,-2823.5</points>
<connection>
<GID>7511</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2823.5,151,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2808,151,-2808</points>
<connection>
<GID>7507</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2823.5,180,-2823.5</points>
<connection>
<GID>7515</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2823.5,174,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2808,174,-2808</points>
<connection>
<GID>7513</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2823.5,205,-2823.5</points>
<connection>
<GID>7519</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2823.5,199,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2808,199,-2808</points>
<connection>
<GID>7517</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2823.5,228,-2823.5</points>
<connection>
<GID>7523</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2823.5,222,-2808</points>
<intersection>-2823.5 1</intersection>
<intersection>-2808 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2808,222,-2808</points>
<connection>
<GID>7521</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2811,215,-2811</points>
<connection>
<GID>7521</GID>
<name>clock</name></connection>
<connection>
<GID>7517</GID>
<name>clock</name></connection>
<connection>
<GID>7513</GID>
<name>clock</name></connection>
<connection>
<GID>7507</GID>
<name>clock</name></connection>
<connection>
<GID>7501</GID>
<name>clock</name></connection>
<connection>
<GID>7493</GID>
<name>clock</name></connection>
<connection>
<GID>7487</GID>
<name>clock</name></connection>
<connection>
<GID>7451</GID>
<name>clock</name></connection>
<connection>
<GID>7445</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2820.5,226,-2820.5</points>
<connection>
<GID>7523</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7519</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7515</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7511</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7505</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7497</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7489</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7463</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7447</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2805,63,-2805</points>
<connection>
<GID>7531</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2805,57,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2789.5,57,-2789.5</points>
<connection>
<GID>7529</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2805,86,-2805</points>
<connection>
<GID>7535</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2805,80,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2789.5,80,-2789.5</points>
<connection>
<GID>7533</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2805,111,-2805</points>
<connection>
<GID>7539</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2805,105,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2789.5,105,-2789.5</points>
<connection>
<GID>7537</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2805,134,-2805</points>
<connection>
<GID>7543</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2805,128,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2789.5,128,-2789.5</points>
<connection>
<GID>7541</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2805,157,-2805</points>
<connection>
<GID>7547</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2805,151,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2789.5,151,-2789.5</points>
<connection>
<GID>7545</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2805,180,-2805</points>
<connection>
<GID>7551</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2805,174,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2789.5,174,-2789.5</points>
<connection>
<GID>7549</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2805,205,-2805</points>
<connection>
<GID>7555</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2805,199,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2789.5,199,-2789.5</points>
<connection>
<GID>7553</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2805,228,-2805</points>
<connection>
<GID>7559</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2805,222,-2789.5</points>
<intersection>-2805 1</intersection>
<intersection>-2789.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2789.5,222,-2789.5</points>
<connection>
<GID>7557</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2792.5,215,-2792.5</points>
<connection>
<GID>7557</GID>
<name>clock</name></connection>
<connection>
<GID>7553</GID>
<name>clock</name></connection>
<connection>
<GID>7549</GID>
<name>clock</name></connection>
<connection>
<GID>7545</GID>
<name>clock</name></connection>
<connection>
<GID>7541</GID>
<name>clock</name></connection>
<connection>
<GID>7537</GID>
<name>clock</name></connection>
<connection>
<GID>7533</GID>
<name>clock</name></connection>
<connection>
<GID>7529</GID>
<name>clock</name></connection>
<connection>
<GID>7525</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2802,226,-2802</points>
<connection>
<GID>7559</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7555</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7551</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7547</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7543</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7539</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7535</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7531</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7527</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2786,63,-2786</points>
<connection>
<GID>7567</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2786,57,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2770.5,57,-2770.5</points>
<connection>
<GID>7565</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2786,86,-2786</points>
<connection>
<GID>7571</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2786,80,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2770.5,80,-2770.5</points>
<connection>
<GID>7569</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2786,111,-2786</points>
<connection>
<GID>7575</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2786,105,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2770.5,105,-2770.5</points>
<connection>
<GID>7573</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2786,134,-2786</points>
<connection>
<GID>7579</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2786,128,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2770.5,128,-2770.5</points>
<connection>
<GID>7577</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2786,157,-2786</points>
<connection>
<GID>7220</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2786,151,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2770.5,151,-2770.5</points>
<connection>
<GID>7581</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2786,180,-2786</points>
<connection>
<GID>7224</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2786,174,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2770.5,174,-2770.5</points>
<connection>
<GID>7222</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2786,205,-2786</points>
<connection>
<GID>7228</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2786,199,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2770.5,199,-2770.5</points>
<connection>
<GID>7226</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2786,228,-2786</points>
<connection>
<GID>7232</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2786,222,-2770.5</points>
<intersection>-2786 1</intersection>
<intersection>-2770.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2770.5,222,-2770.5</points>
<connection>
<GID>7230</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2773.5,215,-2773.5</points>
<connection>
<GID>7581</GID>
<name>clock</name></connection>
<connection>
<GID>7577</GID>
<name>clock</name></connection>
<connection>
<GID>7573</GID>
<name>clock</name></connection>
<connection>
<GID>7569</GID>
<name>clock</name></connection>
<connection>
<GID>7565</GID>
<name>clock</name></connection>
<connection>
<GID>7561</GID>
<name>OUT</name></connection>
<connection>
<GID>7230</GID>
<name>clock</name></connection>
<connection>
<GID>7226</GID>
<name>clock</name></connection>
<connection>
<GID>7222</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2783,226,-2783</points>
<connection>
<GID>7579</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7575</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7571</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7567</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7563</GID>
<name>OUT</name></connection>
<connection>
<GID>7232</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7228</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7224</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7220</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2767.5,63,-2767.5</points>
<connection>
<GID>7240</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2767.5,57,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2752,57,-2752</points>
<connection>
<GID>7238</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2767.5,86,-2767.5</points>
<connection>
<GID>7244</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2767.5,80,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2752,80,-2752</points>
<connection>
<GID>7242</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2767.5,111,-2767.5</points>
<connection>
<GID>7248</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2767.5,105,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2752,105,-2752</points>
<connection>
<GID>7246</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2767.5,134,-2767.5</points>
<connection>
<GID>7252</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2767.5,128,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2752,128,-2752</points>
<connection>
<GID>7250</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2767.5,157,-2767.5</points>
<connection>
<GID>7256</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2767.5,151,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2752,151,-2752</points>
<connection>
<GID>7254</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2767.5,180,-2767.5</points>
<connection>
<GID>7260</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2767.5,174,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2752,174,-2752</points>
<connection>
<GID>7258</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2767.5,205,-2767.5</points>
<connection>
<GID>7264</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2767.5,199,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2752,199,-2752</points>
<connection>
<GID>7262</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2767.5,228,-2767.5</points>
<connection>
<GID>7268</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2767.5,222,-2752</points>
<intersection>-2767.5 1</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2752,222,-2752</points>
<connection>
<GID>7266</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2755,215,-2755</points>
<connection>
<GID>7266</GID>
<name>clock</name></connection>
<connection>
<GID>7262</GID>
<name>clock</name></connection>
<connection>
<GID>7258</GID>
<name>clock</name></connection>
<connection>
<GID>7254</GID>
<name>clock</name></connection>
<connection>
<GID>7250</GID>
<name>clock</name></connection>
<connection>
<GID>7246</GID>
<name>clock</name></connection>
<connection>
<GID>7242</GID>
<name>clock</name></connection>
<connection>
<GID>7238</GID>
<name>clock</name></connection>
<connection>
<GID>7234</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2764.5,226,-2764.5</points>
<connection>
<GID>7268</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7264</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7260</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7256</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7252</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7248</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7244</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7240</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7236</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2901.5,63,-2901.5</points>
<connection>
<GID>7277</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2901.5,57,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2886,57,-2886</points>
<connection>
<GID>7274</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2901.5,86,-2901.5</points>
<connection>
<GID>7282</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2901.5,80,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2886,80,-2886</points>
<connection>
<GID>7279</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2901.5,111,-2901.5</points>
<connection>
<GID>7287</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2901.5,105,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2886,105,-2886</points>
<connection>
<GID>7284</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2901.5,134,-2901.5</points>
<connection>
<GID>7292</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2901.5,128,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2886,128,-2886</points>
<connection>
<GID>7289</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2901.5,157,-2901.5</points>
<connection>
<GID>7297</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2901.5,151,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2886,151,-2886</points>
<connection>
<GID>7294</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2901.5,180,-2901.5</points>
<connection>
<GID>7302</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2901.5,174,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2886,174,-2886</points>
<connection>
<GID>7299</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2901.5,205,-2901.5</points>
<connection>
<GID>7369</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2901.5,199,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2886,199,-2886</points>
<connection>
<GID>7368</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2901.5,228,-2901.5</points>
<connection>
<GID>7371</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2901.5,222,-2886</points>
<intersection>-2901.5 1</intersection>
<intersection>-2886 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2886,222,-2886</points>
<connection>
<GID>7370</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2889,215,-2889</points>
<connection>
<GID>7370</GID>
<name>clock</name></connection>
<connection>
<GID>7368</GID>
<name>clock</name></connection>
<connection>
<GID>7299</GID>
<name>clock</name></connection>
<connection>
<GID>7294</GID>
<name>clock</name></connection>
<connection>
<GID>7289</GID>
<name>clock</name></connection>
<connection>
<GID>7284</GID>
<name>clock</name></connection>
<connection>
<GID>7279</GID>
<name>clock</name></connection>
<connection>
<GID>7274</GID>
<name>clock</name></connection>
<connection>
<GID>7270</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2898.5,226,-2898.5</points>
<connection>
<GID>7371</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7369</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7302</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7297</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7292</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7287</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7282</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7277</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7272</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2883,63,-2883</points>
<connection>
<GID>7375</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2883,57,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2867.5,57,-2867.5</points>
<connection>
<GID>7374</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2883,86,-2883</points>
<connection>
<GID>7377</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2883,80,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2867.5,80,-2867.5</points>
<connection>
<GID>7376</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2883,111,-2883</points>
<connection>
<GID>7379</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2883,105,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2867.5,105,-2867.5</points>
<connection>
<GID>7378</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2883,134,-2883</points>
<connection>
<GID>7381</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2883,128,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2867.5,128,-2867.5</points>
<connection>
<GID>7380</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2883,157,-2883</points>
<connection>
<GID>7383</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2883,151,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2867.5,151,-2867.5</points>
<connection>
<GID>7382</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2883,180,-2883</points>
<connection>
<GID>7385</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2883,174,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2867.5,174,-2867.5</points>
<connection>
<GID>7384</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2883,205,-2883</points>
<connection>
<GID>7387</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2883,199,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2867.5,199,-2867.5</points>
<connection>
<GID>7386</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2883,228,-2883</points>
<connection>
<GID>7389</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2883,222,-2867.5</points>
<intersection>-2883 1</intersection>
<intersection>-2867.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2867.5,222,-2867.5</points>
<connection>
<GID>7388</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2870.5,215,-2870.5</points>
<connection>
<GID>7388</GID>
<name>clock</name></connection>
<connection>
<GID>7386</GID>
<name>clock</name></connection>
<connection>
<GID>7384</GID>
<name>clock</name></connection>
<connection>
<GID>7382</GID>
<name>clock</name></connection>
<connection>
<GID>7380</GID>
<name>clock</name></connection>
<connection>
<GID>7378</GID>
<name>clock</name></connection>
<connection>
<GID>7376</GID>
<name>clock</name></connection>
<connection>
<GID>7374</GID>
<name>clock</name></connection>
<connection>
<GID>7372</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2880,226,-2880</points>
<connection>
<GID>7389</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7387</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7385</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7383</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7381</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7379</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7377</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7375</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7373</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2864,63,-2864</points>
<connection>
<GID>7285</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2864,57,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2848.5,57,-2848.5</points>
<connection>
<GID>7280</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2864,86,-2864</points>
<connection>
<GID>7295</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2864,80,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2848.5,80,-2848.5</points>
<connection>
<GID>7290</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2864,111,-2864</points>
<connection>
<GID>7304</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2864,105,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2848.5,105,-2848.5</points>
<connection>
<GID>7300</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2864,134,-2864</points>
<connection>
<GID>7391</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2864,128,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2848.5,128,-2848.5</points>
<connection>
<GID>7307</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2864,157,-2864</points>
<connection>
<GID>7393</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2864,151,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2848.5,151,-2848.5</points>
<connection>
<GID>7392</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2864,180,-2864</points>
<connection>
<GID>7395</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2864,174,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2848.5,174,-2848.5</points>
<connection>
<GID>7394</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2864,205,-2864</points>
<connection>
<GID>7397</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2864,199,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2848.5,199,-2848.5</points>
<connection>
<GID>7396</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2864,228,-2864</points>
<connection>
<GID>7400</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2864,222,-2848.5</points>
<intersection>-2864 1</intersection>
<intersection>-2848.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2848.5,222,-2848.5</points>
<connection>
<GID>7399</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2851.5,215,-2851.5</points>
<connection>
<GID>7399</GID>
<name>clock</name></connection>
<connection>
<GID>7396</GID>
<name>clock</name></connection>
<connection>
<GID>7394</GID>
<name>clock</name></connection>
<connection>
<GID>7392</GID>
<name>clock</name></connection>
<connection>
<GID>7390</GID>
<name>OUT</name></connection>
<connection>
<GID>7307</GID>
<name>clock</name></connection>
<connection>
<GID>7300</GID>
<name>clock</name></connection>
<connection>
<GID>7290</GID>
<name>clock</name></connection>
<connection>
<GID>7280</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2861,226,-2861</points>
<connection>
<GID>7400</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7397</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7395</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7393</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7391</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7304</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7295</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7285</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7275</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-2845.5,63,-2845.5</points>
<connection>
<GID>7405</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-2845.5,57,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56,-2830,57,-2830</points>
<connection>
<GID>7404</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire>
<wire>
<ID>5233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-2845.5,86,-2845.5</points>
<connection>
<GID>7407</GID>
<name>IN_0</name></connection>
<intersection>80 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>80,-2845.5,80,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-2830,80,-2830</points>
<connection>
<GID>7406</GID>
<name>OUT_0</name></connection>
<intersection>80 2</intersection></hsegment></shape></wire>
<wire>
<ID>5234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-2845.5,111,-2845.5</points>
<connection>
<GID>7410</GID>
<name>IN_0</name></connection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,-2845.5,105,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,-2830,105,-2830</points>
<connection>
<GID>7409</GID>
<name>OUT_0</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>5235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-2845.5,134,-2845.5</points>
<connection>
<GID>7412</GID>
<name>IN_0</name></connection>
<intersection>128 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>128,-2845.5,128,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127,-2830,128,-2830</points>
<connection>
<GID>7411</GID>
<name>OUT_0</name></connection>
<intersection>128 2</intersection></hsegment></shape></wire>
<wire>
<ID>5236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-2845.5,157,-2845.5</points>
<connection>
<GID>7415</GID>
<name>IN_0</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-2845.5,151,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150,-2830,151,-2830</points>
<connection>
<GID>7413</GID>
<name>OUT_0</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>5237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-2845.5,180,-2845.5</points>
<connection>
<GID>7417</GID>
<name>IN_0</name></connection>
<intersection>174 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174,-2845.5,174,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>173,-2830,174,-2830</points>
<connection>
<GID>7416</GID>
<name>OUT_0</name></connection>
<intersection>174 2</intersection></hsegment></shape></wire>
<wire>
<ID>5238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2845.5,205,-2845.5</points>
<connection>
<GID>7419</GID>
<name>IN_0</name></connection>
<intersection>199 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>199,-2845.5,199,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-2830,199,-2830</points>
<connection>
<GID>7418</GID>
<name>OUT_0</name></connection>
<intersection>199 2</intersection></hsegment></shape></wire>
<wire>
<ID>5239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-2845.5,228,-2845.5</points>
<connection>
<GID>7421</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-2845.5,222,-2830</points>
<intersection>-2845.5 1</intersection>
<intersection>-2830 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-2830,222,-2830</points>
<connection>
<GID>7420</GID>
<name>OUT_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>5240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-2833,215,-2833</points>
<connection>
<GID>7420</GID>
<name>clock</name></connection>
<connection>
<GID>7418</GID>
<name>clock</name></connection>
<connection>
<GID>7416</GID>
<name>clock</name></connection>
<connection>
<GID>7413</GID>
<name>clock</name></connection>
<connection>
<GID>7411</GID>
<name>clock</name></connection>
<connection>
<GID>7409</GID>
<name>clock</name></connection>
<connection>
<GID>7406</GID>
<name>clock</name></connection>
<connection>
<GID>7404</GID>
<name>clock</name></connection>
<connection>
<GID>7401</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-2842.5,226,-2842.5</points>
<connection>
<GID>7421</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7419</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7417</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7415</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7412</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7410</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7407</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7405</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7402</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-2911.5,44.5,-2746.5</points>
<connection>
<GID>7449</GID>
<name>N_in1</name></connection>
<connection>
<GID>7422</GID>
<name>N_in0</name></connection>
<intersection>-2886 12</intersection>
<intersection>-2867.5 11</intersection>
<intersection>-2848.5 10</intersection>
<intersection>-2830 9</intersection>
<intersection>-2808 8</intersection>
<intersection>-2789.5 7</intersection>
<intersection>-2770.5 6</intersection>
<intersection>-2752 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-2752,50,-2752</points>
<connection>
<GID>7238</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>44.5,-2770.5,50,-2770.5</points>
<connection>
<GID>7565</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-2789.5,50,-2789.5</points>
<connection>
<GID>7529</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>44.5,-2808,50,-2808</points>
<connection>
<GID>7451</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>44.5,-2830,50,-2830</points>
<connection>
<GID>7404</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>44.5,-2848.5,50,-2848.5</points>
<connection>
<GID>7280</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>44.5,-2867.5,50,-2867.5</points>
<connection>
<GID>7374</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>44.5,-2886,50,-2886</points>
<connection>
<GID>7274</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-2911,67.5,-2746</points>
<connection>
<GID>7453</GID>
<name>N_in1</name></connection>
<connection>
<GID>7423</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 4</intersection>
<intersection>-2875 5</intersection>
<intersection>-2856 6</intersection>
<intersection>-2837.5 7</intersection>
<intersection>-2815.5 8</intersection>
<intersection>-2797 9</intersection>
<intersection>-2778 10</intersection>
<intersection>-2759.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63,-2893.5,67.5,-2893.5</points>
<intersection>63 12</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-2875,67.5,-2875</points>
<intersection>63 14</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>63,-2856,67.5,-2856</points>
<intersection>63 13</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>63,-2837.5,67.5,-2837.5</points>
<intersection>63 15</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>63,-2815.5,67.5,-2815.5</points>
<intersection>63 18</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-2797,67.5,-2797</points>
<intersection>63 19</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>63,-2778,67.5,-2778</points>
<intersection>63 20</intersection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>63,-2759.5,67.5,-2759.5</points>
<intersection>63 21</intersection>
<intersection>67.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>63,-2896,63,-2893.5</points>
<connection>
<GID>7277</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>63,-2858.5,63,-2856</points>
<connection>
<GID>7285</GID>
<name>OUT_0</name></connection>
<intersection>-2856 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>63,-2877.5,63,-2875</points>
<connection>
<GID>7375</GID>
<name>OUT_0</name></connection>
<intersection>-2875 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>63,-2840,63,-2837.5</points>
<connection>
<GID>7405</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>63,-2818,63,-2815.5</points>
<connection>
<GID>7463</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>63,-2799.5,63,-2797</points>
<connection>
<GID>7531</GID>
<name>OUT_0</name></connection>
<intersection>-2797 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>63,-2780.5,63,-2778</points>
<connection>
<GID>7567</GID>
<name>OUT_0</name></connection>
<intersection>-2778 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>63,-2762,63,-2759.5</points>
<connection>
<GID>7240</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-2911,70.5,-2746.5</points>
<connection>
<GID>7455</GID>
<name>N_in1</name></connection>
<connection>
<GID>7424</GID>
<name>N_in0</name></connection>
<intersection>-2886 10</intersection>
<intersection>-2867.5 9</intersection>
<intersection>-2848.5 8</intersection>
<intersection>-2830 7</intersection>
<intersection>-2808 6</intersection>
<intersection>-2789.5 5</intersection>
<intersection>-2770.5 4</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70.5,-2752,73,-2752</points>
<connection>
<GID>7242</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-2770.5,73,-2770.5</points>
<connection>
<GID>7569</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-2789.5,73,-2789.5</points>
<connection>
<GID>7533</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>70.5,-2808,73,-2808</points>
<connection>
<GID>7487</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>70.5,-2830,73,-2830</points>
<connection>
<GID>7406</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>70.5,-2848.5,73,-2848.5</points>
<connection>
<GID>7290</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>70.5,-2867.5,73,-2867.5</points>
<connection>
<GID>7376</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>70.5,-2886,73,-2886</points>
<connection>
<GID>7279</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-2911,90,-2746</points>
<connection>
<GID>7457</GID>
<name>N_in1</name></connection>
<connection>
<GID>7425</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 6</intersection>
<intersection>-2875 7</intersection>
<intersection>-2856 8</intersection>
<intersection>-2837.5 9</intersection>
<intersection>-2815.5 10</intersection>
<intersection>-2797 11</intersection>
<intersection>-2778 12</intersection>
<intersection>-2759.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86,-2893.5,90,-2893.5</points>
<intersection>86 14</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>86,-2875,90,-2875</points>
<intersection>86 16</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>86,-2856,90,-2856</points>
<intersection>86 15</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>86,-2837.5,90,-2837.5</points>
<intersection>86 17</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>86,-2815.5,90,-2815.5</points>
<intersection>86 20</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>86,-2797,90,-2797</points>
<intersection>86 21</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>86,-2778,90,-2778</points>
<intersection>86 22</intersection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>86,-2759.5,90,-2759.5</points>
<intersection>86 23</intersection>
<intersection>90 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>86,-2896,86,-2893.5</points>
<connection>
<GID>7282</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>86,-2858.5,86,-2856</points>
<connection>
<GID>7295</GID>
<name>OUT_0</name></connection>
<intersection>-2856 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>86,-2877.5,86,-2875</points>
<connection>
<GID>7377</GID>
<name>OUT_0</name></connection>
<intersection>-2875 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>86,-2840,86,-2837.5</points>
<connection>
<GID>7407</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>86,-2818,86,-2815.5</points>
<connection>
<GID>7489</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>86,-2799.5,86,-2797</points>
<connection>
<GID>7535</GID>
<name>OUT_0</name></connection>
<intersection>-2797 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>86,-2780.5,86,-2778</points>
<connection>
<GID>7571</GID>
<name>OUT_0</name></connection>
<intersection>-2778 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>86,-2762,86,-2759.5</points>
<connection>
<GID>7244</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-2911,93.5,-2746</points>
<connection>
<GID>7459</GID>
<name>N_in1</name></connection>
<connection>
<GID>7426</GID>
<name>N_in0</name></connection>
<intersection>-2886 13</intersection>
<intersection>-2867.5 12</intersection>
<intersection>-2848.5 11</intersection>
<intersection>-2830 10</intersection>
<intersection>-2808 9</intersection>
<intersection>-2789.5 8</intersection>
<intersection>-2770.5 7</intersection>
<intersection>-2752 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>93.5,-2752,98,-2752</points>
<connection>
<GID>7246</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>93.5,-2770.5,98,-2770.5</points>
<connection>
<GID>7573</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>93.5,-2789.5,98,-2789.5</points>
<connection>
<GID>7537</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>93.5,-2808,98,-2808</points>
<connection>
<GID>7493</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>93.5,-2830,98,-2830</points>
<connection>
<GID>7409</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>93.5,-2848.5,98,-2848.5</points>
<connection>
<GID>7300</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>93.5,-2867.5,98,-2867.5</points>
<connection>
<GID>7378</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>93.5,-2886,98,-2886</points>
<connection>
<GID>7284</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2911,114.5,-2746.5</points>
<connection>
<GID>7461</GID>
<name>N_in1</name></connection>
<connection>
<GID>7427</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 6</intersection>
<intersection>-2875 7</intersection>
<intersection>-2856 8</intersection>
<intersection>-2837.5 9</intersection>
<intersection>-2815.5 10</intersection>
<intersection>-2797 11</intersection>
<intersection>-2778 12</intersection>
<intersection>-2759.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>111,-2893.5,114.5,-2893.5</points>
<intersection>111 14</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111,-2875,114.5,-2875</points>
<intersection>111 16</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111,-2856,114.5,-2856</points>
<intersection>111 15</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111,-2837.5,114.5,-2837.5</points>
<intersection>111 17</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,-2815.5,114.5,-2815.5</points>
<intersection>111 20</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>111,-2797,114.5,-2797</points>
<intersection>111 21</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>111,-2778,114.5,-2778</points>
<intersection>111 22</intersection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111,-2759.5,114.5,-2759.5</points>
<intersection>111 23</intersection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>111,-2896,111,-2893.5</points>
<connection>
<GID>7287</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>111,-2858.5,111,-2856</points>
<connection>
<GID>7304</GID>
<name>OUT_0</name></connection>
<intersection>-2856 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>111,-2877.5,111,-2875</points>
<connection>
<GID>7379</GID>
<name>OUT_0</name></connection>
<intersection>-2875 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>111,-2840,111,-2837.5</points>
<connection>
<GID>7410</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>111,-2818,111,-2815.5</points>
<connection>
<GID>7497</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>111,-2799.5,111,-2797</points>
<connection>
<GID>7539</GID>
<name>OUT_0</name></connection>
<intersection>-2797 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>111,-2780.5,111,-2778</points>
<connection>
<GID>7575</GID>
<name>OUT_0</name></connection>
<intersection>-2778 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>111,-2762,111,-2759.5</points>
<connection>
<GID>7248</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-2911,118.5,-2746</points>
<connection>
<GID>7465</GID>
<name>N_in1</name></connection>
<connection>
<GID>7428</GID>
<name>N_in0</name></connection>
<intersection>-2886 13</intersection>
<intersection>-2867.5 12</intersection>
<intersection>-2848.5 11</intersection>
<intersection>-2830 10</intersection>
<intersection>-2808 9</intersection>
<intersection>-2789.5 8</intersection>
<intersection>-2770.5 7</intersection>
<intersection>-2752 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>118.5,-2752,121,-2752</points>
<connection>
<GID>7250</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>118.5,-2770.5,121,-2770.5</points>
<connection>
<GID>7577</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118.5,-2789.5,121,-2789.5</points>
<connection>
<GID>7541</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>118.5,-2808,121,-2808</points>
<connection>
<GID>7501</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>118.5,-2830,121,-2830</points>
<connection>
<GID>7411</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>118.5,-2848.5,121,-2848.5</points>
<connection>
<GID>7307</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>118.5,-2867.5,121,-2867.5</points>
<connection>
<GID>7380</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>118.5,-2886,121,-2886</points>
<connection>
<GID>7289</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2911,137,-2746</points>
<connection>
<GID>7467</GID>
<name>N_in1</name></connection>
<connection>
<GID>7429</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 6</intersection>
<intersection>-2875 7</intersection>
<intersection>-2856 8</intersection>
<intersection>-2837.5 9</intersection>
<intersection>-2815.5 10</intersection>
<intersection>-2797 11</intersection>
<intersection>-2778 12</intersection>
<intersection>-2759.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>134,-2893.5,137,-2893.5</points>
<intersection>134 14</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>134,-2875,137,-2875</points>
<intersection>134 15</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>134,-2856,137,-2856</points>
<intersection>134 16</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>134,-2837.5,137,-2837.5</points>
<intersection>134 17</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>134,-2815.5,137,-2815.5</points>
<intersection>134 20</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>134,-2797,137,-2797</points>
<intersection>134 21</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>134,-2778,137,-2778</points>
<intersection>134 22</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>134,-2759.5,137,-2759.5</points>
<intersection>134 23</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>134,-2896,134,-2893.5</points>
<connection>
<GID>7292</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>134,-2877.5,134,-2875</points>
<connection>
<GID>7381</GID>
<name>OUT_0</name></connection>
<intersection>-2875 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>134,-2858.5,134,-2856</points>
<connection>
<GID>7391</GID>
<name>OUT_0</name></connection>
<intersection>-2856 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>134,-2840,134,-2837.5</points>
<connection>
<GID>7412</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>134,-2818,134,-2815.5</points>
<connection>
<GID>7505</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>134,-2799.5,134,-2797</points>
<connection>
<GID>7543</GID>
<name>OUT_0</name></connection>
<intersection>-2797 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>134,-2780.5,134,-2778</points>
<connection>
<GID>7579</GID>
<name>OUT_0</name></connection>
<intersection>-2778 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>134,-2762,134,-2759.5</points>
<connection>
<GID>7252</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-2911,141,-2746</points>
<connection>
<GID>7469</GID>
<name>N_in1</name></connection>
<connection>
<GID>7431</GID>
<name>N_in0</name></connection>
<intersection>-2886 13</intersection>
<intersection>-2867.5 12</intersection>
<intersection>-2848.5 11</intersection>
<intersection>-2830 10</intersection>
<intersection>-2808 9</intersection>
<intersection>-2789.5 8</intersection>
<intersection>-2770.5 7</intersection>
<intersection>-2752 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>141,-2752,144,-2752</points>
<connection>
<GID>7254</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>141,-2770.5,144,-2770.5</points>
<connection>
<GID>7581</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>141,-2789.5,144,-2789.5</points>
<connection>
<GID>7545</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>141,-2808,144,-2808</points>
<connection>
<GID>7507</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>141,-2830,144,-2830</points>
<connection>
<GID>7413</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>141,-2848.5,144,-2848.5</points>
<connection>
<GID>7392</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>141,-2867.5,144,-2867.5</points>
<connection>
<GID>7382</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>141,-2886,144,-2886</points>
<connection>
<GID>7294</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>5251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-2910.5,160,-2746</points>
<connection>
<GID>7471</GID>
<name>N_in1</name></connection>
<connection>
<GID>7433</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 6</intersection>
<intersection>-2875 7</intersection>
<intersection>-2856 8</intersection>
<intersection>-2837.5 9</intersection>
<intersection>-2815.5 10</intersection>
<intersection>-2797 11</intersection>
<intersection>-2778 12</intersection>
<intersection>-2759.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>157,-2893.5,160,-2893.5</points>
<intersection>157 15</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>157,-2875,160,-2875</points>
<intersection>157 16</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>157,-2856,160,-2856</points>
<intersection>157 17</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,-2837.5,160,-2837.5</points>
<intersection>157 18</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>157,-2815.5,160,-2815.5</points>
<intersection>157 21</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>157,-2797,160,-2797</points>
<intersection>157 22</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>157,-2778,160,-2778</points>
<intersection>157 23</intersection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>157,-2759.5,160,-2759.5</points>
<intersection>157 14</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>157,-2762,157,-2759.5</points>
<connection>
<GID>7256</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>157,-2896,157,-2893.5</points>
<connection>
<GID>7297</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>157,-2877.5,157,-2875</points>
<connection>
<GID>7383</GID>
<name>OUT_0</name></connection>
<intersection>-2875 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>157,-2858.5,157,-2856</points>
<connection>
<GID>7393</GID>
<name>OUT_0</name></connection>
<intersection>-2856 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>157,-2840,157,-2837.5</points>
<connection>
<GID>7415</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>157,-2818,157,-2815.5</points>
<connection>
<GID>7511</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>157,-2799.5,157,-2797</points>
<connection>
<GID>7547</GID>
<name>OUT_0</name></connection>
<intersection>-2797 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>157,-2780.5,157,-2778</points>
<connection>
<GID>7220</GID>
<name>OUT_0</name></connection>
<intersection>-2778 12</intersection></vsegment></shape></wire>
<wire>
<ID>5252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-2910.5,165,-2746</points>
<connection>
<GID>7473</GID>
<name>N_in1</name></connection>
<connection>
<GID>7435</GID>
<name>N_in0</name></connection>
<intersection>-2886 13</intersection>
<intersection>-2867.5 12</intersection>
<intersection>-2848.5 11</intersection>
<intersection>-2830 10</intersection>
<intersection>-2808 9</intersection>
<intersection>-2789.5 8</intersection>
<intersection>-2770.5 7</intersection>
<intersection>-2752 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>165,-2752,167,-2752</points>
<connection>
<GID>7258</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>165,-2770.5,167,-2770.5</points>
<connection>
<GID>7222</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>165,-2789.5,167,-2789.5</points>
<connection>
<GID>7549</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>165,-2808,167,-2808</points>
<connection>
<GID>7513</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>165,-2830,167,-2830</points>
<connection>
<GID>7416</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>165,-2848.5,167,-2848.5</points>
<connection>
<GID>7394</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>165,-2867.5,167,-2867.5</points>
<connection>
<GID>7384</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>165,-2886,167,-2886</points>
<connection>
<GID>7299</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>5253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-2910,183,-2746</points>
<connection>
<GID>7475</GID>
<name>N_in1</name></connection>
<connection>
<GID>7439</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 16</intersection>
<intersection>-2875 15</intersection>
<intersection>-2856 14</intersection>
<intersection>-2837.5 13</intersection>
<intersection>-2815.5 12</intersection>
<intersection>-2797 11</intersection>
<intersection>-2778 10</intersection>
<intersection>-2759.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>180,-2759.5,183,-2759.5</points>
<intersection>180 17</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>180,-2778,183,-2778</points>
<intersection>180 26</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>180,-2797,183,-2797</points>
<intersection>180 25</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>180,-2815.5,183,-2815.5</points>
<intersection>180 24</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>180,-2837.5,183,-2837.5</points>
<intersection>180 21</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>180,-2856,183,-2856</points>
<intersection>180 20</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>180,-2875,183,-2875</points>
<intersection>180 19</intersection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>180,-2893.5,183,-2893.5</points>
<intersection>180 18</intersection>
<intersection>183 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>180,-2762,180,-2759.5</points>
<connection>
<GID>7260</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>180,-2896,180,-2893.5</points>
<connection>
<GID>7302</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>180,-2877.5,180,-2875</points>
<connection>
<GID>7385</GID>
<name>OUT_0</name></connection>
<intersection>-2875 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>180,-2858.5,180,-2856</points>
<connection>
<GID>7395</GID>
<name>OUT_0</name></connection>
<intersection>-2856 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>180,-2840,180,-2837.5</points>
<connection>
<GID>7417</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>180,-2818,180,-2815.5</points>
<connection>
<GID>7515</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>180,-2799.5,180,-2797</points>
<connection>
<GID>7551</GID>
<name>OUT_0</name></connection>
<intersection>-2797 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>180,-2780.5,180,-2778</points>
<connection>
<GID>7224</GID>
<name>OUT_0</name></connection>
<intersection>-2778 10</intersection></vsegment></shape></wire>
<wire>
<ID>5254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-2910,187.5,-2746</points>
<connection>
<GID>7477</GID>
<name>N_in1</name></connection>
<connection>
<GID>7437</GID>
<name>N_in0</name></connection>
<intersection>-2886 13</intersection>
<intersection>-2867.5 12</intersection>
<intersection>-2848.5 11</intersection>
<intersection>-2830 10</intersection>
<intersection>-2808 9</intersection>
<intersection>-2789.5 8</intersection>
<intersection>-2770.5 7</intersection>
<intersection>-2752 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>187.5,-2752,192,-2752</points>
<connection>
<GID>7262</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>187.5,-2770.5,192,-2770.5</points>
<connection>
<GID>7226</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187.5,-2789.5,192,-2789.5</points>
<connection>
<GID>7553</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>187.5,-2808,192,-2808</points>
<connection>
<GID>7517</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>187.5,-2830,192,-2830</points>
<connection>
<GID>7418</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>187.5,-2848.5,192,-2848.5</points>
<connection>
<GID>7396</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>187.5,-2867.5,192,-2867.5</points>
<connection>
<GID>7386</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>187.5,-2886,192,-2886</points>
<connection>
<GID>7368</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-2909.5,208.5,-2746.5</points>
<connection>
<GID>7479</GID>
<name>N_in1</name></connection>
<connection>
<GID>7441</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 6</intersection>
<intersection>-2875 7</intersection>
<intersection>-2856 8</intersection>
<intersection>-2837.5 9</intersection>
<intersection>-2815.5 10</intersection>
<intersection>-2797 11</intersection>
<intersection>-2778 12</intersection>
<intersection>-2759.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>205,-2893.5,208.5,-2893.5</points>
<intersection>205 15</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205,-2875,208.5,-2875</points>
<intersection>205 16</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>205,-2856,208.5,-2856</points>
<intersection>205 17</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>205,-2837.5,208.5,-2837.5</points>
<intersection>205 18</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>205,-2815.5,208.5,-2815.5</points>
<intersection>205 21</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205,-2797,208.5,-2797</points>
<intersection>205 22</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>205,-2778,208.5,-2778</points>
<intersection>205 23</intersection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>205,-2759.5,208.5,-2759.5</points>
<intersection>205 14</intersection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>205,-2762,205,-2759.5</points>
<connection>
<GID>7264</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>205,-2896,205,-2893.5</points>
<connection>
<GID>7369</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>205,-2877.5,205,-2875</points>
<connection>
<GID>7387</GID>
<name>OUT_0</name></connection>
<intersection>-2875 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>205,-2858.5,205,-2856</points>
<connection>
<GID>7397</GID>
<name>OUT_0</name></connection>
<intersection>-2856 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>205,-2840,205,-2837.5</points>
<connection>
<GID>7419</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>205,-2818,205,-2815.5</points>
<connection>
<GID>7519</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>205,-2799.5,205,-2797</points>
<connection>
<GID>7555</GID>
<name>OUT_0</name></connection>
<intersection>-2797 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>205,-2780.5,205,-2778</points>
<connection>
<GID>7228</GID>
<name>OUT_0</name></connection>
<intersection>-2778 12</intersection></vsegment></shape></wire>
<wire>
<ID>5256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-2909.5,212,-2746.5</points>
<connection>
<GID>7481</GID>
<name>N_in1</name></connection>
<connection>
<GID>7483</GID>
<name>N_in0</name></connection>
<intersection>-2886 11</intersection>
<intersection>-2867.5 10</intersection>
<intersection>-2848.5 9</intersection>
<intersection>-2830 7</intersection>
<intersection>-2808 6</intersection>
<intersection>-2789.5 5</intersection>
<intersection>-2770.5 4</intersection>
<intersection>-2752 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-2752,215,-2752</points>
<connection>
<GID>7266</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>212,-2770.5,215,-2770.5</points>
<connection>
<GID>7230</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>212,-2789.5,215,-2789.5</points>
<connection>
<GID>7557</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>212,-2808,215,-2808</points>
<connection>
<GID>7521</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>212,-2830,215,-2830</points>
<connection>
<GID>7420</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>212,-2848.5,215,-2848.5</points>
<connection>
<GID>7399</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>212,-2867.5,215,-2867.5</points>
<connection>
<GID>7388</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>212,-2886,215,-2886</points>
<connection>
<GID>7370</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>5257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-2909.5,233,-2747.5</points>
<connection>
<GID>7485</GID>
<name>N_in1</name></connection>
<connection>
<GID>7443</GID>
<name>N_in0</name></connection>
<intersection>-2893.5 11</intersection>
<intersection>-2875 10</intersection>
<intersection>-2856 9</intersection>
<intersection>-2837.5 8</intersection>
<intersection>-2815.5 7</intersection>
<intersection>-2797 6</intersection>
<intersection>-2778 5</intersection>
<intersection>-2759.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>228,-2759.5,233,-2759.5</points>
<intersection>228 12</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-2778,233,-2778</points>
<intersection>228 21</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>228,-2797,233,-2797</points>
<intersection>228 20</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>228,-2815.5,233,-2815.5</points>
<intersection>228 19</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>228,-2837.5,233,-2837.5</points>
<intersection>228 16</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>228,-2856,233,-2856</points>
<intersection>228 15</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>228,-2875,233,-2875</points>
<intersection>228 14</intersection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>228,-2893.5,233,-2893.5</points>
<intersection>228 13</intersection>
<intersection>233 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>228,-2762,228,-2759.5</points>
<connection>
<GID>7268</GID>
<name>OUT_0</name></connection>
<intersection>-2759.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>228,-2896,228,-2893.5</points>
<connection>
<GID>7371</GID>
<name>OUT_0</name></connection>
<intersection>-2893.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>228,-2877.5,228,-2875</points>
<connection>
<GID>7389</GID>
<name>OUT_0</name></connection>
<intersection>-2875 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>228,-2858.5,228,-2856</points>
<connection>
<GID>7400</GID>
<name>OUT_0</name></connection>
<intersection>-2856 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>228,-2840,228,-2837.5</points>
<connection>
<GID>7421</GID>
<name>OUT_0</name></connection>
<intersection>-2837.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>228,-2818,228,-2815.5</points>
<connection>
<GID>7523</GID>
<name>OUT_0</name></connection>
<intersection>-2815.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>228,-2799.5,228,-2797</points>
<connection>
<GID>7559</GID>
<name>OUT_0</name></connection>
<intersection>-2797 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>228,-2780.5,228,-2778</points>
<connection>
<GID>7232</GID>
<name>OUT_0</name></connection>
<intersection>-2778 5</intersection></vsegment></shape></wire>
<wire>
<ID>5258</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-117,-2754,22.5,-2754</points>
<connection>
<GID>7234</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-117,-2763.5,-117,-2738</points>
<intersection>-2763.5 4</intersection>
<intersection>-2754 2</intersection>
<intersection>-2738 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-117,-2763.5,34,-2763.5</points>
<connection>
<GID>7236</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-2738,-117,-2738</points>
<connection>
<GID>7367</GID>
<name>OUT_7</name></connection>
<intersection>-117 3</intersection></hsegment></shape></wire>
<wire>
<ID>5259</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-118,-2772.5,22.5,-2772.5</points>
<connection>
<GID>7561</GID>
<name>IN_0</name></connection>
<intersection>-118 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-118,-2782,-118,-2739</points>
<intersection>-2782 5</intersection>
<intersection>-2772.5 2</intersection>
<intersection>-2739 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-118,-2782,34,-2782</points>
<connection>
<GID>7563</GID>
<name>IN_0</name></connection>
<intersection>-118 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-2739,-118,-2739</points>
<connection>
<GID>7367</GID>
<name>OUT_6</name></connection>
<intersection>-118 4</intersection></hsegment></shape></wire>
<wire>
<ID>5260</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-119,-2791.5,22.5,-2791.5</points>
<connection>
<GID>7525</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119,-2801,-119,-2740</points>
<intersection>-2801 4</intersection>
<intersection>-2791.5 2</intersection>
<intersection>-2740 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-119,-2801,34,-2801</points>
<connection>
<GID>7527</GID>
<name>IN_0</name></connection>
<intersection>-119 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-124,-2740,-119,-2740</points>
<connection>
<GID>7367</GID>
<name>OUT_5</name></connection>
<intersection>-119 3</intersection></hsegment></shape></wire>
<wire>
<ID>5261</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-120,-2810,22.5,-2810</points>
<connection>
<GID>7445</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-2819.5,-120,-2741</points>
<intersection>-2819.5 4</intersection>
<intersection>-2810 2</intersection>
<intersection>-2741 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-120,-2819.5,34,-2819.5</points>
<connection>
<GID>7447</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2741,-120,-2741</points>
<connection>
<GID>7367</GID>
<name>OUT_4</name></connection>
<intersection>-120 3</intersection></hsegment></shape></wire>
<wire>
<ID>5262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-2832,22.5,-2832</points>
<connection>
<GID>7401</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-121,-2841.5,-121,-2742</points>
<intersection>-2841.5 4</intersection>
<intersection>-2832 1</intersection>
<intersection>-2742 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-121,-2841.5,33.5,-2841.5</points>
<connection>
<GID>7402</GID>
<name>IN_0</name></connection>
<intersection>-121 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2742,-121,-2742</points>
<connection>
<GID>7367</GID>
<name>OUT_3</name></connection>
<intersection>-121 3</intersection></hsegment></shape></wire>
<wire>
<ID>5263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-2850.5,22.5,-2850.5</points>
<connection>
<GID>7390</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122,-2860,-122,-2743</points>
<intersection>-2860 4</intersection>
<intersection>-2850.5 1</intersection>
<intersection>-2743 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-122,-2860,33.5,-2860</points>
<connection>
<GID>7275</GID>
<name>IN_0</name></connection>
<intersection>-122 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2743,-122,-2743</points>
<connection>
<GID>7367</GID>
<name>OUT_2</name></connection>
<intersection>-122 3</intersection></hsegment></shape></wire>
<wire>
<ID>5264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123,-2869.5,22.5,-2869.5</points>
<connection>
<GID>7372</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-123,-2879,-123,-2744</points>
<intersection>-2879 4</intersection>
<intersection>-2869.5 1</intersection>
<intersection>-2744 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-123,-2879,33.5,-2879</points>
<connection>
<GID>7373</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-124,-2744,-123,-2744</points>
<connection>
<GID>7367</GID>
<name>OUT_1</name></connection>
<intersection>-123 3</intersection></hsegment></shape></wire>
<wire>
<ID>5265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,-2888,22.5,-2888</points>
<connection>
<GID>7270</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-124,-2897.5,-124,-2745</points>
<connection>
<GID>7367</GID>
<name>OUT_0</name></connection>
<intersection>-2897.5 4</intersection>
<intersection>-2888 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-124,-2897.5,33.5,-2897.5</points>
<connection>
<GID>7272</GID>
<name>IN_0</name></connection>
<intersection>-124 3</intersection></hsegment></shape></wire>
<wire>
<ID>5266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-2911.5,21.5,-2746.5</points>
<connection>
<GID>7503</GID>
<name>N_in1</name></connection>
<connection>
<GID>7495</GID>
<name>N_in0</name></connection>
<intersection>-2890 10</intersection>
<intersection>-2871.5 9</intersection>
<intersection>-2852.5 8</intersection>
<intersection>-2834 7</intersection>
<intersection>-2812 6</intersection>
<intersection>-2793.5 5</intersection>
<intersection>-2774.5 4</intersection>
<intersection>-2756 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-2756,22.5,-2756</points>
<connection>
<GID>7234</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-2774.5,22.5,-2774.5</points>
<connection>
<GID>7561</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>21.5,-2793.5,22.5,-2793.5</points>
<connection>
<GID>7525</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-2812,22.5,-2812</points>
<connection>
<GID>7445</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21.5,-2834,22.5,-2834</points>
<connection>
<GID>7401</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>21.5,-2852.5,22.5,-2852.5</points>
<connection>
<GID>7390</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>21.5,-2871.5,22.5,-2871.5</points>
<connection>
<GID>7372</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>21.5,-2890,22.5,-2890</points>
<connection>
<GID>7270</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-2911.5,31.5,-2746.5</points>
<connection>
<GID>7499</GID>
<name>N_in1</name></connection>
<connection>
<GID>7491</GID>
<name>N_in0</name></connection>
<intersection>-2899.5 3</intersection>
<intersection>-2881 5</intersection>
<intersection>-2862 7</intersection>
<intersection>-2843.5 9</intersection>
<intersection>-2821.5 11</intersection>
<intersection>-2803 13</intersection>
<intersection>-2784 15</intersection>
<intersection>-2765.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-2899.5,33.5,-2899.5</points>
<connection>
<GID>7272</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-2881,33.5,-2881</points>
<connection>
<GID>7373</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31.5,-2862,33.5,-2862</points>
<connection>
<GID>7275</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>31.5,-2843.5,33.5,-2843.5</points>
<connection>
<GID>7402</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>31.5,-2821.5,34,-2821.5</points>
<connection>
<GID>7447</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>31.5,-2803,34,-2803</points>
<connection>
<GID>7527</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>31.5,-2784,34,-2784</points>
<connection>
<GID>7563</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>31.5,-2765.5,34,-2765.5</points>
<connection>
<GID>7236</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-2744.5,21.5,-2738</points>
<connection>
<GID>7495</GID>
<name>N_in1</name></connection>
<connection>
<GID>7365</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-2744.5,31.5,-2738</points>
<connection>
<GID>7491</GID>
<name>N_in1</name></connection>
<connection>
<GID>7364</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-2744.5,44.5,-2738</points>
<connection>
<GID>7422</GID>
<name>N_in1</name></connection>
<connection>
<GID>7345</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-2744,67.5,-2737.5</points>
<connection>
<GID>7423</GID>
<name>N_in1</name></connection>
<connection>
<GID>7346</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-2744.5,70.5,-2737.5</points>
<connection>
<GID>7424</GID>
<name>N_in1</name></connection>
<connection>
<GID>7347</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-2744,90,-2737.5</points>
<connection>
<GID>7425</GID>
<name>N_in1</name></connection>
<connection>
<GID>7348</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-2744,93.5,-2737.5</points>
<connection>
<GID>7426</GID>
<name>N_in1</name></connection>
<connection>
<GID>7349</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-2744.5,114.5,-2737.5</points>
<connection>
<GID>7427</GID>
<name>N_in1</name></connection>
<connection>
<GID>7350</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-2744,118.5,-2737.5</points>
<connection>
<GID>7428</GID>
<name>N_in1</name></connection>
<connection>
<GID>7351</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-2744,137,-2737.5</points>
<connection>
<GID>7429</GID>
<name>N_in1</name></connection>
<connection>
<GID>7352</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-2744,141,-2737.5</points>
<connection>
<GID>7431</GID>
<name>N_in1</name></connection>
<connection>
<GID>7353</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-2744,160,-2737</points>
<connection>
<GID>7433</GID>
<name>N_in1</name></connection>
<connection>
<GID>7354</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-2744,165,-2737</points>
<connection>
<GID>7435</GID>
<name>N_in1</name></connection>
<connection>
<GID>7355</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-2744,183,-2736.5</points>
<connection>
<GID>7439</GID>
<name>N_in1</name></connection>
<connection>
<GID>7356</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-2744,187.5,-2736.5</points>
<connection>
<GID>7437</GID>
<name>N_in1</name></connection>
<connection>
<GID>7357</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-2744.5,208.5,-2736</points>
<connection>
<GID>7441</GID>
<name>N_in1</name></connection>
<connection>
<GID>7358</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-2744.5,212,-2736</points>
<connection>
<GID>7483</GID>
<name>N_in1</name></connection>
<connection>
<GID>7359</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-2745.5,233,-2736</points>
<connection>
<GID>7443</GID>
<name>N_in1</name></connection>
<connection>
<GID>7361</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3040,54,-3040</points>
<connection>
<GID>7779</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3040,48,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3024.5,48,-3024.5</points>
<connection>
<GID>7773</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3040,77,-3040</points>
<connection>
<GID>7797</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3040,71,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3024.5,71,-3024.5</points>
<connection>
<GID>7795</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3040,102,-3040</points>
<connection>
<GID>7801</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3040,96,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3024.5,96,-3024.5</points>
<connection>
<GID>7799</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3040,125,-3040</points>
<connection>
<GID>7805</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3040,119,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3024.5,119,-3024.5</points>
<connection>
<GID>7803</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3040,148,-3040</points>
<connection>
<GID>7809</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3040,142,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3024.5,142,-3024.5</points>
<connection>
<GID>7807</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3040,171,-3040</points>
<connection>
<GID>7813</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3040,165,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3024.5,165,-3024.5</points>
<connection>
<GID>7811</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3040,196,-3040</points>
<connection>
<GID>7817</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3040,190,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3024.5,190,-3024.5</points>
<connection>
<GID>7815</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3040,219,-3040</points>
<connection>
<GID>7821</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3040,213,-3024.5</points>
<intersection>-3040 1</intersection>
<intersection>-3024.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3024.5,213,-3024.5</points>
<connection>
<GID>7819</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3027.5,206,-3027.5</points>
<connection>
<GID>7819</GID>
<name>clock</name></connection>
<connection>
<GID>7815</GID>
<name>clock</name></connection>
<connection>
<GID>7811</GID>
<name>clock</name></connection>
<connection>
<GID>7807</GID>
<name>clock</name></connection>
<connection>
<GID>7803</GID>
<name>clock</name></connection>
<connection>
<GID>7799</GID>
<name>clock</name></connection>
<connection>
<GID>7795</GID>
<name>clock</name></connection>
<connection>
<GID>7773</GID>
<name>clock</name></connection>
<connection>
<GID>7763</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3037,217,-3037</points>
<connection>
<GID>7821</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7817</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7813</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7809</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7805</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7801</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7797</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7779</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7768</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3021.5,54,-3021.5</points>
<connection>
<GID>7829</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3021.5,48,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3006,48,-3006</points>
<connection>
<GID>7827</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3021.5,77,-3021.5</points>
<connection>
<GID>7833</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3021.5,71,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3006,71,-3006</points>
<connection>
<GID>7831</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3021.5,102,-3021.5</points>
<connection>
<GID>7837</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3021.5,96,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3006,96,-3006</points>
<connection>
<GID>7835</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3021.5,125,-3021.5</points>
<connection>
<GID>7841</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3021.5,119,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3006,119,-3006</points>
<connection>
<GID>7839</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3021.5,148,-3021.5</points>
<connection>
<GID>7845</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3021.5,142,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3006,142,-3006</points>
<connection>
<GID>7843</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3021.5,171,-3021.5</points>
<connection>
<GID>7849</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3021.5,165,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3006,165,-3006</points>
<connection>
<GID>7847</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3021.5,196,-3021.5</points>
<connection>
<GID>7853</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3021.5,190,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3006,190,-3006</points>
<connection>
<GID>7851</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5303</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3021.5,219,-3021.5</points>
<connection>
<GID>7857</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3021.5,213,-3006</points>
<intersection>-3021.5 1</intersection>
<intersection>-3006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3006,213,-3006</points>
<connection>
<GID>7855</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3009,206,-3009</points>
<connection>
<GID>7855</GID>
<name>clock</name></connection>
<connection>
<GID>7851</GID>
<name>clock</name></connection>
<connection>
<GID>7847</GID>
<name>clock</name></connection>
<connection>
<GID>7843</GID>
<name>clock</name></connection>
<connection>
<GID>7839</GID>
<name>clock</name></connection>
<connection>
<GID>7835</GID>
<name>clock</name></connection>
<connection>
<GID>7831</GID>
<name>clock</name></connection>
<connection>
<GID>7827</GID>
<name>clock</name></connection>
<connection>
<GID>7823</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3018.5,217,-3018.5</points>
<connection>
<GID>7857</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7853</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7849</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7845</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7841</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7837</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7833</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7829</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7825</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3002.5,54,-3002.5</points>
<connection>
<GID>7865</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3002.5,48,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-2987,48,-2987</points>
<connection>
<GID>7863</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3002.5,77,-3002.5</points>
<connection>
<GID>7869</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3002.5,71,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-2987,71,-2987</points>
<connection>
<GID>7867</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3002.5,102,-3002.5</points>
<connection>
<GID>7873</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3002.5,96,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-2987,96,-2987</points>
<connection>
<GID>7871</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5309</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3002.5,125,-3002.5</points>
<connection>
<GID>7877</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3002.5,119,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-2987,119,-2987</points>
<connection>
<GID>7875</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3002.5,148,-3002.5</points>
<connection>
<GID>7881</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3002.5,142,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-2987,142,-2987</points>
<connection>
<GID>7879</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3002.5,171,-3002.5</points>
<connection>
<GID>7885</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3002.5,165,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-2987,165,-2987</points>
<connection>
<GID>7883</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3002.5,196,-3002.5</points>
<connection>
<GID>7889</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3002.5,190,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-2987,190,-2987</points>
<connection>
<GID>7887</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3002.5,219,-3002.5</points>
<connection>
<GID>7893</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3002.5,213,-2987</points>
<intersection>-3002.5 1</intersection>
<intersection>-2987 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-2987,213,-2987</points>
<connection>
<GID>7891</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-2990,206,-2990</points>
<connection>
<GID>7891</GID>
<name>clock</name></connection>
<connection>
<GID>7887</GID>
<name>clock</name></connection>
<connection>
<GID>7883</GID>
<name>clock</name></connection>
<connection>
<GID>7879</GID>
<name>clock</name></connection>
<connection>
<GID>7875</GID>
<name>clock</name></connection>
<connection>
<GID>7871</GID>
<name>clock</name></connection>
<connection>
<GID>7867</GID>
<name>clock</name></connection>
<connection>
<GID>7863</GID>
<name>clock</name></connection>
<connection>
<GID>7859</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-2999.5,217,-2999.5</points>
<connection>
<GID>7893</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7889</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7885</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7881</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7877</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7873</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7869</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7865</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7861</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-2984,54,-2984</points>
<connection>
<GID>7901</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-2984,48,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-2968.5,48,-2968.5</points>
<connection>
<GID>7899</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-2984,77,-2984</points>
<connection>
<GID>7905</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-2984,71,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-2968.5,71,-2968.5</points>
<connection>
<GID>7903</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-2984,102,-2984</points>
<connection>
<GID>7909</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-2984,96,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-2968.5,96,-2968.5</points>
<connection>
<GID>7907</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-2984,125,-2984</points>
<connection>
<GID>7913</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-2984,119,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-2968.5,119,-2968.5</points>
<connection>
<GID>7911</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-2984,148,-2984</points>
<connection>
<GID>7917</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-2984,142,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-2968.5,142,-2968.5</points>
<connection>
<GID>7915</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-2984,171,-2984</points>
<connection>
<GID>7921</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-2984,165,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-2968.5,165,-2968.5</points>
<connection>
<GID>7919</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-2984,196,-2984</points>
<connection>
<GID>7925</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-2984,190,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-2968.5,190,-2968.5</points>
<connection>
<GID>7923</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-2984,219,-2984</points>
<connection>
<GID>7929</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-2984,213,-2968.5</points>
<intersection>-2984 1</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-2968.5,213,-2968.5</points>
<connection>
<GID>7927</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-2971.5,206,-2971.5</points>
<connection>
<GID>7927</GID>
<name>clock</name></connection>
<connection>
<GID>7923</GID>
<name>clock</name></connection>
<connection>
<GID>7919</GID>
<name>clock</name></connection>
<connection>
<GID>7915</GID>
<name>clock</name></connection>
<connection>
<GID>7911</GID>
<name>clock</name></connection>
<connection>
<GID>7907</GID>
<name>clock</name></connection>
<connection>
<GID>7903</GID>
<name>clock</name></connection>
<connection>
<GID>7899</GID>
<name>clock</name></connection>
<connection>
<GID>7895</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-2981,217,-2981</points>
<connection>
<GID>7929</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7925</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7921</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7917</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7913</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7909</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7905</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7901</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7897</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5326</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3118,54,-3118</points>
<connection>
<GID>7937</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3118,48,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3102.5,48,-3102.5</points>
<connection>
<GID>7935</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3118,77,-3118</points>
<connection>
<GID>7941</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3118,71,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3102.5,71,-3102.5</points>
<connection>
<GID>7939</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3118,102,-3118</points>
<connection>
<GID>7945</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3118,96,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3102.5,96,-3102.5</points>
<connection>
<GID>7943</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3118,125,-3118</points>
<connection>
<GID>7586</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3118,119,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3102.5,119,-3102.5</points>
<connection>
<GID>7584</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3118,148,-3118</points>
<connection>
<GID>7590</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3118,142,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3102.5,142,-3102.5</points>
<connection>
<GID>7588</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3118,171,-3118</points>
<connection>
<GID>7594</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3118,165,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3102.5,165,-3102.5</points>
<connection>
<GID>7592</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3118,196,-3118</points>
<connection>
<GID>7598</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3118,190,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3102.5,190,-3102.5</points>
<connection>
<GID>7596</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3118,219,-3118</points>
<connection>
<GID>7602</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3118,213,-3102.5</points>
<intersection>-3118 1</intersection>
<intersection>-3102.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3102.5,213,-3102.5</points>
<connection>
<GID>7600</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3105.5,206,-3105.5</points>
<connection>
<GID>7943</GID>
<name>clock</name></connection>
<connection>
<GID>7939</GID>
<name>clock</name></connection>
<connection>
<GID>7935</GID>
<name>clock</name></connection>
<connection>
<GID>7931</GID>
<name>OUT</name></connection>
<connection>
<GID>7600</GID>
<name>clock</name></connection>
<connection>
<GID>7596</GID>
<name>clock</name></connection>
<connection>
<GID>7592</GID>
<name>clock</name></connection>
<connection>
<GID>7588</GID>
<name>clock</name></connection>
<connection>
<GID>7584</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3115,217,-3115</points>
<connection>
<GID>7945</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7941</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7937</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7933</GID>
<name>OUT</name></connection>
<connection>
<GID>7602</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7598</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7594</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7590</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7586</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3099.5,54,-3099.5</points>
<connection>
<GID>7610</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3099.5,48,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3084,48,-3084</points>
<connection>
<GID>7608</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5337</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3099.5,77,-3099.5</points>
<connection>
<GID>7614</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3099.5,71,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3084,71,-3084</points>
<connection>
<GID>7612</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3099.5,102,-3099.5</points>
<connection>
<GID>7618</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3099.5,96,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3084,96,-3084</points>
<connection>
<GID>7616</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3099.5,125,-3099.5</points>
<connection>
<GID>7622</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3099.5,119,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3084,119,-3084</points>
<connection>
<GID>7620</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5340</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3099.5,148,-3099.5</points>
<connection>
<GID>7626</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3099.5,142,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3084,142,-3084</points>
<connection>
<GID>7624</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3099.5,171,-3099.5</points>
<connection>
<GID>7630</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3099.5,165,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3084,165,-3084</points>
<connection>
<GID>7628</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3099.5,196,-3099.5</points>
<connection>
<GID>7634</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3099.5,190,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3084,190,-3084</points>
<connection>
<GID>7632</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3099.5,219,-3099.5</points>
<connection>
<GID>7638</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3099.5,213,-3084</points>
<intersection>-3099.5 1</intersection>
<intersection>-3084 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3084,213,-3084</points>
<connection>
<GID>7636</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3087,206,-3087</points>
<connection>
<GID>7636</GID>
<name>clock</name></connection>
<connection>
<GID>7632</GID>
<name>clock</name></connection>
<connection>
<GID>7628</GID>
<name>clock</name></connection>
<connection>
<GID>7624</GID>
<name>clock</name></connection>
<connection>
<GID>7620</GID>
<name>clock</name></connection>
<connection>
<GID>7616</GID>
<name>clock</name></connection>
<connection>
<GID>7612</GID>
<name>clock</name></connection>
<connection>
<GID>7608</GID>
<name>clock</name></connection>
<connection>
<GID>7604</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3096.5,217,-3096.5</points>
<connection>
<GID>7638</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7634</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7630</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7626</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7622</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7618</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7614</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7610</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7606</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3080.5,54,-3080.5</points>
<connection>
<GID>7648</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3080.5,48,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3065,48,-3065</points>
<connection>
<GID>7646</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3080.5,77,-3080.5</points>
<connection>
<GID>7653</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3080.5,71,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3065,71,-3065</points>
<connection>
<GID>7651</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3080.5,102,-3080.5</points>
<connection>
<GID>7658</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3080.5,96,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3065,96,-3065</points>
<connection>
<GID>7656</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3080.5,125,-3080.5</points>
<connection>
<GID>7663</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3080.5,119,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3065,119,-3065</points>
<connection>
<GID>7661</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3080.5,148,-3080.5</points>
<connection>
<GID>7668</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3080.5,142,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3065,142,-3065</points>
<connection>
<GID>7666</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3080.5,171,-3080.5</points>
<connection>
<GID>7671</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3080.5,165,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3065,165,-3065</points>
<connection>
<GID>7670</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3080.5,196,-3080.5</points>
<connection>
<GID>7674</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3080.5,190,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3065,190,-3065</points>
<connection>
<GID>7673</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3080.5,219,-3080.5</points>
<connection>
<GID>7676</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3080.5,213,-3065</points>
<intersection>-3080.5 1</intersection>
<intersection>-3065 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3065,213,-3065</points>
<connection>
<GID>7675</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3068,206,-3068</points>
<connection>
<GID>7675</GID>
<name>clock</name></connection>
<connection>
<GID>7673</GID>
<name>clock</name></connection>
<connection>
<GID>7670</GID>
<name>clock</name></connection>
<connection>
<GID>7666</GID>
<name>clock</name></connection>
<connection>
<GID>7661</GID>
<name>clock</name></connection>
<connection>
<GID>7656</GID>
<name>clock</name></connection>
<connection>
<GID>7651</GID>
<name>clock</name></connection>
<connection>
<GID>7646</GID>
<name>clock</name></connection>
<connection>
<GID>7641</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5355</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3077.5,217,-3077.5</points>
<connection>
<GID>7676</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7674</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7671</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7668</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7663</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7658</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7653</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7648</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7643</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5356</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3062,54,-3062</points>
<connection>
<GID>7680</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3062,48,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3046.5,48,-3046.5</points>
<connection>
<GID>7679</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3062,77,-3062</points>
<connection>
<GID>7682</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3062,71,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3046.5,71,-3046.5</points>
<connection>
<GID>7681</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5358</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3062,102,-3062</points>
<connection>
<GID>7684</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3062,96,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3046.5,96,-3046.5</points>
<connection>
<GID>7683</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5359</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3062,125,-3062</points>
<connection>
<GID>7686</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3062,119,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3046.5,119,-3046.5</points>
<connection>
<GID>7685</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3062,148,-3062</points>
<connection>
<GID>7688</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3062,142,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3046.5,142,-3046.5</points>
<connection>
<GID>7687</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5361</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3062,171,-3062</points>
<connection>
<GID>7690</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3062,165,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3046.5,165,-3046.5</points>
<connection>
<GID>7689</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5362</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3062,196,-3062</points>
<connection>
<GID>7692</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3062,190,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3046.5,190,-3046.5</points>
<connection>
<GID>7691</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3062,219,-3062</points>
<connection>
<GID>7694</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3062,213,-3046.5</points>
<intersection>-3062 1</intersection>
<intersection>-3046.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3046.5,213,-3046.5</points>
<connection>
<GID>7693</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3049.5,206,-3049.5</points>
<connection>
<GID>7693</GID>
<name>clock</name></connection>
<connection>
<GID>7691</GID>
<name>clock</name></connection>
<connection>
<GID>7689</GID>
<name>clock</name></connection>
<connection>
<GID>7687</GID>
<name>clock</name></connection>
<connection>
<GID>7685</GID>
<name>clock</name></connection>
<connection>
<GID>7683</GID>
<name>clock</name></connection>
<connection>
<GID>7681</GID>
<name>clock</name></connection>
<connection>
<GID>7679</GID>
<name>clock</name></connection>
<connection>
<GID>7677</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3059,217,-3059</points>
<connection>
<GID>7694</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7692</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7690</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7688</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7686</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7684</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7682</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7678</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-3128,35.5,-2963</points>
<connection>
<GID>7710</GID>
<name>N_in1</name></connection>
<connection>
<GID>7695</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 12</intersection>
<intersection>-3084 11</intersection>
<intersection>-3065 10</intersection>
<intersection>-3046.5 9</intersection>
<intersection>-3024.5 8</intersection>
<intersection>-3006 7</intersection>
<intersection>-2987 6</intersection>
<intersection>-2968.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-2968.5,41,-2968.5</points>
<connection>
<GID>7899</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-2987,41,-2987</points>
<connection>
<GID>7863</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-3006,41,-3006</points>
<connection>
<GID>7827</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-3024.5,41,-3024.5</points>
<connection>
<GID>7773</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>35.5,-3046.5,41,-3046.5</points>
<connection>
<GID>7679</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>35.5,-3065,41,-3065</points>
<connection>
<GID>7646</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>35.5,-3084,41,-3084</points>
<connection>
<GID>7608</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>35.5,-3102.5,41,-3102.5</points>
<connection>
<GID>7935</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-3127.5,58.5,-2962.5</points>
<connection>
<GID>7711</GID>
<name>N_in1</name></connection>
<connection>
<GID>7696</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 4</intersection>
<intersection>-3092 5</intersection>
<intersection>-3073 6</intersection>
<intersection>-3054.5 7</intersection>
<intersection>-3032.5 8</intersection>
<intersection>-3014 9</intersection>
<intersection>-2995 10</intersection>
<intersection>-2976.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-3110.5,58.5,-3110.5</points>
<intersection>54 12</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54,-3092,58.5,-3092</points>
<intersection>54 13</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54,-3073,58.5,-3073</points>
<intersection>54 14</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54,-3054.5,58.5,-3054.5</points>
<intersection>54 15</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-3032.5,58.5,-3032.5</points>
<intersection>54 18</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>54,-3014,58.5,-3014</points>
<intersection>54 19</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>54,-2995,58.5,-2995</points>
<intersection>54 20</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>54,-2976.5,58.5,-2976.5</points>
<intersection>54 21</intersection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>54,-3112.5,54,-3110.5</points>
<connection>
<GID>7937</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>54,-3094,54,-3092</points>
<connection>
<GID>7610</GID>
<name>OUT_0</name></connection>
<intersection>-3092 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>54,-3075,54,-3073</points>
<connection>
<GID>7648</GID>
<name>OUT_0</name></connection>
<intersection>-3073 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>54,-3056.5,54,-3054.5</points>
<connection>
<GID>7680</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>54,-3034.5,54,-3032.5</points>
<connection>
<GID>7779</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>54,-3016,54,-3014</points>
<connection>
<GID>7829</GID>
<name>OUT_0</name></connection>
<intersection>-3014 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>54,-2997,54,-2995</points>
<connection>
<GID>7865</GID>
<name>OUT_0</name></connection>
<intersection>-2995 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>54,-2978.5,54,-2976.5</points>
<connection>
<GID>7901</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-3127.5,61.5,-2963</points>
<connection>
<GID>7712</GID>
<name>N_in1</name></connection>
<connection>
<GID>7697</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 10</intersection>
<intersection>-3084 9</intersection>
<intersection>-3065 8</intersection>
<intersection>-3046.5 7</intersection>
<intersection>-3024.5 6</intersection>
<intersection>-3006 5</intersection>
<intersection>-2987 4</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-2968.5,64,-2968.5</points>
<connection>
<GID>7903</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-2987,64,-2987</points>
<connection>
<GID>7867</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61.5,-3006,64,-3006</points>
<connection>
<GID>7831</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61.5,-3024.5,64,-3024.5</points>
<connection>
<GID>7795</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61.5,-3046.5,64,-3046.5</points>
<connection>
<GID>7681</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61.5,-3065,64,-3065</points>
<connection>
<GID>7651</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61.5,-3084,64,-3084</points>
<connection>
<GID>7612</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61.5,-3102.5,64,-3102.5</points>
<connection>
<GID>7939</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-3127.5,81,-2962.5</points>
<connection>
<GID>7713</GID>
<name>N_in1</name></connection>
<connection>
<GID>7698</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 6</intersection>
<intersection>-3092 7</intersection>
<intersection>-3073 8</intersection>
<intersection>-3054.5 9</intersection>
<intersection>-3032.5 10</intersection>
<intersection>-3014 11</intersection>
<intersection>-2995 12</intersection>
<intersection>-2976.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-3110.5,81,-3110.5</points>
<intersection>77 14</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>77,-3092,81,-3092</points>
<intersection>77 15</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>77,-3073,81,-3073</points>
<intersection>77 16</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-3054.5,81,-3054.5</points>
<intersection>77 17</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>77,-3032.5,81,-3032.5</points>
<intersection>77 20</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>77,-3014,81,-3014</points>
<intersection>77 21</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>77,-2995,81,-2995</points>
<intersection>77 22</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>77,-2976.5,81,-2976.5</points>
<intersection>77 23</intersection>
<intersection>81 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>77,-3112.5,77,-3110.5</points>
<connection>
<GID>7941</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>77,-3094,77,-3092</points>
<connection>
<GID>7614</GID>
<name>OUT_0</name></connection>
<intersection>-3092 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>77,-3075,77,-3073</points>
<connection>
<GID>7653</GID>
<name>OUT_0</name></connection>
<intersection>-3073 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>77,-3056.5,77,-3054.5</points>
<connection>
<GID>7682</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>77,-3034.5,77,-3032.5</points>
<connection>
<GID>7797</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>77,-3016,77,-3014</points>
<connection>
<GID>7833</GID>
<name>OUT_0</name></connection>
<intersection>-3014 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>77,-2997,77,-2995</points>
<connection>
<GID>7869</GID>
<name>OUT_0</name></connection>
<intersection>-2995 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>77,-2978.5,77,-2976.5</points>
<connection>
<GID>7905</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-3127.5,84.5,-2962.5</points>
<connection>
<GID>7714</GID>
<name>N_in1</name></connection>
<connection>
<GID>7699</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 13</intersection>
<intersection>-3084 12</intersection>
<intersection>-3065 11</intersection>
<intersection>-3046.5 10</intersection>
<intersection>-3024.5 9</intersection>
<intersection>-3006 8</intersection>
<intersection>-2987 7</intersection>
<intersection>-2968.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-2968.5,89,-2968.5</points>
<connection>
<GID>7907</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-2987,89,-2987</points>
<connection>
<GID>7871</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>84.5,-3006,89,-3006</points>
<connection>
<GID>7835</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84.5,-3024.5,89,-3024.5</points>
<connection>
<GID>7799</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84.5,-3046.5,89,-3046.5</points>
<connection>
<GID>7683</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84.5,-3065,89,-3065</points>
<connection>
<GID>7656</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>84.5,-3084,89,-3084</points>
<connection>
<GID>7616</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>84.5,-3102.5,89,-3102.5</points>
<connection>
<GID>7943</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3127.5,105.5,-2963</points>
<connection>
<GID>7715</GID>
<name>N_in1</name></connection>
<connection>
<GID>7700</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 6</intersection>
<intersection>-3092 7</intersection>
<intersection>-3073 8</intersection>
<intersection>-3054.5 9</intersection>
<intersection>-3032.5 10</intersection>
<intersection>-3014 11</intersection>
<intersection>-2995 12</intersection>
<intersection>-2976.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>102,-3110.5,105.5,-3110.5</points>
<intersection>102 14</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>102,-3092,105.5,-3092</points>
<intersection>102 15</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>102,-3073,105.5,-3073</points>
<intersection>102 16</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>102,-3054.5,105.5,-3054.5</points>
<intersection>102 17</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>102,-3032.5,105.5,-3032.5</points>
<intersection>102 20</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>102,-3014,105.5,-3014</points>
<intersection>102 21</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>102,-2995,105.5,-2995</points>
<intersection>102 22</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>102,-2976.5,105.5,-2976.5</points>
<intersection>102 23</intersection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>102,-3112.5,102,-3110.5</points>
<connection>
<GID>7945</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>102,-3094,102,-3092</points>
<connection>
<GID>7618</GID>
<name>OUT_0</name></connection>
<intersection>-3092 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>102,-3075,102,-3073</points>
<connection>
<GID>7658</GID>
<name>OUT_0</name></connection>
<intersection>-3073 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>102,-3056.5,102,-3054.5</points>
<connection>
<GID>7684</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>102,-3034.5,102,-3032.5</points>
<connection>
<GID>7801</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>102,-3016,102,-3014</points>
<connection>
<GID>7837</GID>
<name>OUT_0</name></connection>
<intersection>-3014 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>102,-2997,102,-2995</points>
<connection>
<GID>7873</GID>
<name>OUT_0</name></connection>
<intersection>-2995 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>102,-2978.5,102,-2976.5</points>
<connection>
<GID>7909</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3127.5,109.5,-2962.5</points>
<connection>
<GID>7716</GID>
<name>N_in1</name></connection>
<connection>
<GID>7701</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 13</intersection>
<intersection>-3084 12</intersection>
<intersection>-3065 11</intersection>
<intersection>-3046.5 10</intersection>
<intersection>-3024.5 9</intersection>
<intersection>-3006 8</intersection>
<intersection>-2987 7</intersection>
<intersection>-2968.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109.5,-2968.5,112,-2968.5</points>
<connection>
<GID>7911</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>109.5,-2987,112,-2987</points>
<connection>
<GID>7875</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109.5,-3006,112,-3006</points>
<connection>
<GID>7839</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>109.5,-3024.5,112,-3024.5</points>
<connection>
<GID>7803</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>109.5,-3046.5,112,-3046.5</points>
<connection>
<GID>7685</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>109.5,-3065,112,-3065</points>
<connection>
<GID>7661</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109.5,-3084,112,-3084</points>
<connection>
<GID>7620</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>109.5,-3102.5,112,-3102.5</points>
<connection>
<GID>7584</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-3127.5,128,-2962.5</points>
<connection>
<GID>7717</GID>
<name>N_in1</name></connection>
<connection>
<GID>7702</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 6</intersection>
<intersection>-3092 7</intersection>
<intersection>-3073 8</intersection>
<intersection>-3054.5 9</intersection>
<intersection>-3032.5 10</intersection>
<intersection>-3014 11</intersection>
<intersection>-2995 12</intersection>
<intersection>-2976.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>125,-3110.5,128,-3110.5</points>
<intersection>125 14</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125,-3092,128,-3092</points>
<intersection>125 15</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>125,-3073,128,-3073</points>
<intersection>125 16</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>125,-3054.5,128,-3054.5</points>
<intersection>125 17</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125,-3032.5,128,-3032.5</points>
<intersection>125 20</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>125,-3014,128,-3014</points>
<intersection>125 21</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>125,-2995,128,-2995</points>
<intersection>125 22</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>125,-2976.5,128,-2976.5</points>
<intersection>125 23</intersection>
<intersection>128 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>125,-3112.5,125,-3110.5</points>
<connection>
<GID>7586</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>125,-3094,125,-3092</points>
<connection>
<GID>7622</GID>
<name>OUT_0</name></connection>
<intersection>-3092 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>125,-3075,125,-3073</points>
<connection>
<GID>7663</GID>
<name>OUT_0</name></connection>
<intersection>-3073 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>125,-3056.5,125,-3054.5</points>
<connection>
<GID>7686</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>125,-3034.5,125,-3032.5</points>
<connection>
<GID>7805</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>125,-3016,125,-3014</points>
<connection>
<GID>7841</GID>
<name>OUT_0</name></connection>
<intersection>-3014 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>125,-2997,125,-2995</points>
<connection>
<GID>7877</GID>
<name>OUT_0</name></connection>
<intersection>-2995 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>125,-2978.5,125,-2976.5</points>
<connection>
<GID>7913</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-3127.5,132,-2962.5</points>
<connection>
<GID>7718</GID>
<name>N_in1</name></connection>
<connection>
<GID>7703</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 13</intersection>
<intersection>-3084 12</intersection>
<intersection>-3065 11</intersection>
<intersection>-3046.5 10</intersection>
<intersection>-3024.5 9</intersection>
<intersection>-3006 8</intersection>
<intersection>-2987 7</intersection>
<intersection>-2968.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>132,-2968.5,135,-2968.5</points>
<connection>
<GID>7915</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>132,-2987,135,-2987</points>
<connection>
<GID>7879</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>132,-3006,135,-3006</points>
<connection>
<GID>7843</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>132,-3024.5,135,-3024.5</points>
<connection>
<GID>7807</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132,-3046.5,135,-3046.5</points>
<connection>
<GID>7687</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132,-3065,135,-3065</points>
<connection>
<GID>7666</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>132,-3084,135,-3084</points>
<connection>
<GID>7624</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132,-3102.5,135,-3102.5</points>
<connection>
<GID>7588</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>5375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-3127,151,-2962.5</points>
<connection>
<GID>7719</GID>
<name>N_in1</name></connection>
<connection>
<GID>7704</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 6</intersection>
<intersection>-3092 7</intersection>
<intersection>-3073 8</intersection>
<intersection>-3054.5 9</intersection>
<intersection>-3032.5 10</intersection>
<intersection>-3014 11</intersection>
<intersection>-2995 12</intersection>
<intersection>-2976.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>148,-3110.5,151,-3110.5</points>
<intersection>148 14</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>148,-3092,151,-3092</points>
<intersection>148 15</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>148,-3073,151,-3073</points>
<intersection>148 16</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>148,-3054.5,151,-3054.5</points>
<intersection>148 17</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>148,-3032.5,151,-3032.5</points>
<intersection>148 20</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>148,-3014,151,-3014</points>
<intersection>148 21</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>148,-2995,151,-2995</points>
<intersection>148 22</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>148,-2976.5,151,-2976.5</points>
<intersection>148 23</intersection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>148,-3112.5,148,-3110.5</points>
<connection>
<GID>7590</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>148,-3094,148,-3092</points>
<connection>
<GID>7626</GID>
<name>OUT_0</name></connection>
<intersection>-3092 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>148,-3075,148,-3073</points>
<connection>
<GID>7668</GID>
<name>OUT_0</name></connection>
<intersection>-3073 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>148,-3056.5,148,-3054.5</points>
<connection>
<GID>7688</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>148,-3034.5,148,-3032.5</points>
<connection>
<GID>7809</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>148,-3016,148,-3014</points>
<connection>
<GID>7845</GID>
<name>OUT_0</name></connection>
<intersection>-3014 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>148,-2997,148,-2995</points>
<connection>
<GID>7881</GID>
<name>OUT_0</name></connection>
<intersection>-2995 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>148,-2978.5,148,-2976.5</points>
<connection>
<GID>7917</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-3127,156,-2962.5</points>
<connection>
<GID>7720</GID>
<name>N_in1</name></connection>
<connection>
<GID>7705</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 13</intersection>
<intersection>-3084 12</intersection>
<intersection>-3065 11</intersection>
<intersection>-3046.5 10</intersection>
<intersection>-3024.5 9</intersection>
<intersection>-3006 8</intersection>
<intersection>-2987 7</intersection>
<intersection>-2968.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>156,-2968.5,158,-2968.5</points>
<connection>
<GID>7919</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>156,-2987,158,-2987</points>
<connection>
<GID>7883</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>156,-3006,158,-3006</points>
<connection>
<GID>7847</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>156,-3024.5,158,-3024.5</points>
<connection>
<GID>7811</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156,-3046.5,158,-3046.5</points>
<connection>
<GID>7689</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>156,-3065,158,-3065</points>
<connection>
<GID>7670</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>156,-3084,158,-3084</points>
<connection>
<GID>7628</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>156,-3102.5,158,-3102.5</points>
<connection>
<GID>7592</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>5377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-3126.5,174,-2962.5</points>
<connection>
<GID>7721</GID>
<name>N_in1</name></connection>
<connection>
<GID>7707</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 16</intersection>
<intersection>-3092 15</intersection>
<intersection>-3073 14</intersection>
<intersection>-3054.5 13</intersection>
<intersection>-3032.5 12</intersection>
<intersection>-3014 11</intersection>
<intersection>-2995 10</intersection>
<intersection>-2976.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>171,-2976.5,174,-2976.5</points>
<intersection>171 26</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>171,-2995,174,-2995</points>
<intersection>171 25</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>171,-3014,174,-3014</points>
<intersection>171 24</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>171,-3032.5,174,-3032.5</points>
<intersection>171 23</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>171,-3054.5,174,-3054.5</points>
<intersection>171 20</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>171,-3073,174,-3073</points>
<intersection>171 19</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>171,-3092,174,-3092</points>
<intersection>171 18</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>171,-3110.5,174,-3110.5</points>
<intersection>171 17</intersection>
<intersection>174 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>171,-3112.5,171,-3110.5</points>
<connection>
<GID>7594</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>171,-3094,171,-3092</points>
<connection>
<GID>7630</GID>
<name>OUT_0</name></connection>
<intersection>-3092 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>171,-3075,171,-3073</points>
<connection>
<GID>7671</GID>
<name>OUT_0</name></connection>
<intersection>-3073 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>171,-3056.5,171,-3054.5</points>
<connection>
<GID>7690</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>171,-3034.5,171,-3032.5</points>
<connection>
<GID>7813</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>171,-3016,171,-3014</points>
<connection>
<GID>7849</GID>
<name>OUT_0</name></connection>
<intersection>-3014 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>171,-2997,171,-2995</points>
<connection>
<GID>7885</GID>
<name>OUT_0</name></connection>
<intersection>-2995 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>171,-2978.5,171,-2976.5</points>
<connection>
<GID>7921</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>5378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-3126.5,178.5,-2962.5</points>
<connection>
<GID>7722</GID>
<name>N_in1</name></connection>
<connection>
<GID>7706</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 13</intersection>
<intersection>-3084 12</intersection>
<intersection>-3065 11</intersection>
<intersection>-3046.5 10</intersection>
<intersection>-3024.5 9</intersection>
<intersection>-3006 8</intersection>
<intersection>-2987 7</intersection>
<intersection>-2968.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>178.5,-2968.5,183,-2968.5</points>
<connection>
<GID>7923</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>178.5,-2987,183,-2987</points>
<connection>
<GID>7887</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178.5,-3006,183,-3006</points>
<connection>
<GID>7851</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>178.5,-3024.5,183,-3024.5</points>
<connection>
<GID>7815</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>178.5,-3046.5,183,-3046.5</points>
<connection>
<GID>7691</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>178.5,-3065,183,-3065</points>
<connection>
<GID>7673</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>178.5,-3084,183,-3084</points>
<connection>
<GID>7632</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>178.5,-3102.5,183,-3102.5</points>
<connection>
<GID>7596</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-3126,199.5,-2963</points>
<connection>
<GID>7723</GID>
<name>N_in1</name></connection>
<connection>
<GID>7708</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 6</intersection>
<intersection>-3092 7</intersection>
<intersection>-3073 8</intersection>
<intersection>-3054.5 9</intersection>
<intersection>-3032.5 10</intersection>
<intersection>-3014 11</intersection>
<intersection>-2995 12</intersection>
<intersection>-2976.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196,-3110.5,199.5,-3110.5</points>
<intersection>196 14</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>196,-3092,199.5,-3092</points>
<intersection>196 15</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>196,-3073,199.5,-3073</points>
<intersection>196 16</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>196,-3054.5,199.5,-3054.5</points>
<intersection>196 17</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>196,-3032.5,199.5,-3032.5</points>
<intersection>196 20</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>196,-3014,199.5,-3014</points>
<intersection>196 21</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>196,-2995,199.5,-2995</points>
<intersection>196 22</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>196,-2976.5,199.5,-2976.5</points>
<intersection>196 23</intersection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>196,-3112.5,196,-3110.5</points>
<connection>
<GID>7598</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>196,-3094,196,-3092</points>
<connection>
<GID>7634</GID>
<name>OUT_0</name></connection>
<intersection>-3092 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>196,-3075,196,-3073</points>
<connection>
<GID>7674</GID>
<name>OUT_0</name></connection>
<intersection>-3073 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>196,-3056.5,196,-3054.5</points>
<connection>
<GID>7692</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>196,-3034.5,196,-3032.5</points>
<connection>
<GID>7817</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>196,-3016,196,-3014</points>
<connection>
<GID>7853</GID>
<name>OUT_0</name></connection>
<intersection>-3014 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>196,-2997,196,-2995</points>
<connection>
<GID>7889</GID>
<name>OUT_0</name></connection>
<intersection>-2995 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>196,-2978.5,196,-2976.5</points>
<connection>
<GID>7925</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-3126,203,-2963</points>
<connection>
<GID>7724</GID>
<name>N_in1</name></connection>
<connection>
<GID>7725</GID>
<name>N_in0</name></connection>
<intersection>-3102.5 11</intersection>
<intersection>-3084 10</intersection>
<intersection>-3065 9</intersection>
<intersection>-3046.5 7</intersection>
<intersection>-3024.5 6</intersection>
<intersection>-3006 5</intersection>
<intersection>-2987 4</intersection>
<intersection>-2968.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-2968.5,206,-2968.5</points>
<connection>
<GID>7927</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>203,-2987,206,-2987</points>
<connection>
<GID>7891</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>203,-3006,206,-3006</points>
<connection>
<GID>7855</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>203,-3024.5,206,-3024.5</points>
<connection>
<GID>7819</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-3046.5,206,-3046.5</points>
<connection>
<GID>7693</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>203,-3065,206,-3065</points>
<connection>
<GID>7675</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>203,-3084,206,-3084</points>
<connection>
<GID>7636</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-3102.5,206,-3102.5</points>
<connection>
<GID>7600</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment></shape></wire>
<wire>
<ID>5381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-3126,224,-2964</points>
<connection>
<GID>7726</GID>
<name>N_in1</name></connection>
<connection>
<GID>7709</GID>
<name>N_in0</name></connection>
<intersection>-3110.5 11</intersection>
<intersection>-3092 10</intersection>
<intersection>-3073 9</intersection>
<intersection>-3054.5 8</intersection>
<intersection>-3032.5 7</intersection>
<intersection>-3014 6</intersection>
<intersection>-2995 5</intersection>
<intersection>-2976.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>219,-2976.5,224,-2976.5</points>
<intersection>219 21</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>219,-2995,224,-2995</points>
<intersection>219 20</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>219,-3014,224,-3014</points>
<intersection>219 19</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>219,-3032.5,224,-3032.5</points>
<intersection>219 18</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>219,-3054.5,224,-3054.5</points>
<intersection>219 15</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>219,-3073,224,-3073</points>
<intersection>219 14</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>219,-3092,224,-3092</points>
<intersection>219 13</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>219,-3110.5,224,-3110.5</points>
<intersection>219 12</intersection>
<intersection>224 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>219,-3112.5,219,-3110.5</points>
<connection>
<GID>7602</GID>
<name>OUT_0</name></connection>
<intersection>-3110.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>219,-3094,219,-3092</points>
<connection>
<GID>7638</GID>
<name>OUT_0</name></connection>
<intersection>-3092 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>219,-3075,219,-3073</points>
<connection>
<GID>7676</GID>
<name>OUT_0</name></connection>
<intersection>-3073 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>219,-3056.5,219,-3054.5</points>
<connection>
<GID>7694</GID>
<name>OUT_0</name></connection>
<intersection>-3054.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>219,-3034.5,219,-3032.5</points>
<connection>
<GID>7821</GID>
<name>OUT_0</name></connection>
<intersection>-3032.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>219,-3016,219,-3014</points>
<connection>
<GID>7857</GID>
<name>OUT_0</name></connection>
<intersection>-3014 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>219,-2997,219,-2995</points>
<connection>
<GID>7893</GID>
<name>OUT_0</name></connection>
<intersection>-2995 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>219,-2978.5,219,-2976.5</points>
<connection>
<GID>7929</GID>
<name>OUT_0</name></connection>
<intersection>-2976.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>5382</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-133,-2970.5,13.5,-2970.5</points>
<connection>
<GID>7895</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-133,-3122,-133,-2970.5</points>
<connection>
<GID>7732</GID>
<name>OUT_15</name></connection>
<intersection>-2980 4</intersection>
<intersection>-2970.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-133,-2980,25,-2980</points>
<connection>
<GID>7897</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment></shape></wire>
<wire>
<ID>5383</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-132,-2989,13.5,-2989</points>
<connection>
<GID>7859</GID>
<name>IN_0</name></connection>
<intersection>-132 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-132,-3123,-132,-2989</points>
<intersection>-3123 6</intersection>
<intersection>-2998.5 5</intersection>
<intersection>-2989 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-132,-2998.5,25,-2998.5</points>
<connection>
<GID>7861</GID>
<name>IN_0</name></connection>
<intersection>-132 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3123,-132,-3123</points>
<connection>
<GID>7732</GID>
<name>OUT_14</name></connection>
<intersection>-132 4</intersection></hsegment></shape></wire>
<wire>
<ID>5384</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-131,-3008,13.5,-3008</points>
<connection>
<GID>7823</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-131,-3124,-131,-3008</points>
<intersection>-3124 6</intersection>
<intersection>-3017.5 4</intersection>
<intersection>-3008 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-131,-3017.5,25,-3017.5</points>
<connection>
<GID>7825</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3124,-131,-3124</points>
<connection>
<GID>7732</GID>
<name>OUT_13</name></connection>
<intersection>-131 3</intersection></hsegment></shape></wire>
<wire>
<ID>5385</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-130,-3026.5,13.5,-3026.5</points>
<connection>
<GID>7763</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-130,-3125,-130,-3026.5</points>
<intersection>-3125 5</intersection>
<intersection>-3036 4</intersection>
<intersection>-3026.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-130,-3036,25,-3036</points>
<connection>
<GID>7768</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3125,-130,-3125</points>
<connection>
<GID>7732</GID>
<name>OUT_12</name></connection>
<intersection>-130 3</intersection></hsegment></shape></wire>
<wire>
<ID>5386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-129,-3048.5,13.5,-3048.5</points>
<connection>
<GID>7677</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-129,-3126,-129,-3048.5</points>
<intersection>-3126 6</intersection>
<intersection>-3058 4</intersection>
<intersection>-3048.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-129,-3058,24.5,-3058</points>
<connection>
<GID>7678</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3126,-129,-3126</points>
<connection>
<GID>7732</GID>
<name>OUT_11</name></connection>
<intersection>-129 3</intersection></hsegment></shape></wire>
<wire>
<ID>5387</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-128,-3067,13.5,-3067</points>
<connection>
<GID>7641</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-3127,-128,-3067</points>
<intersection>-3127 5</intersection>
<intersection>-3076.5 4</intersection>
<intersection>-3067 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-3076.5,24.5,-3076.5</points>
<connection>
<GID>7643</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3127,-128,-3127</points>
<connection>
<GID>7732</GID>
<name>OUT_10</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>5388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127,-3086,13.5,-3086</points>
<connection>
<GID>7604</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-127,-3128,-127,-3086</points>
<intersection>-3128 5</intersection>
<intersection>-3095.5 4</intersection>
<intersection>-3086 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-127,-3095.5,24.5,-3095.5</points>
<connection>
<GID>7606</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3128,-127,-3128</points>
<connection>
<GID>7732</GID>
<name>OUT_9</name></connection>
<intersection>-127 3</intersection></hsegment></shape></wire>
<wire>
<ID>5389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,-3104.5,13.5,-3104.5</points>
<connection>
<GID>7931</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-3129,-126,-3104.5</points>
<intersection>-3129 5</intersection>
<intersection>-3114 4</intersection>
<intersection>-3104.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-3114,24.5,-3114</points>
<connection>
<GID>7933</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3129,-126,-3129</points>
<connection>
<GID>7732</GID>
<name>OUT_8</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>5390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-3128,12.5,-2963</points>
<connection>
<GID>7730</GID>
<name>N_in1</name></connection>
<connection>
<GID>7728</GID>
<name>N_in0</name></connection>
<intersection>-3106.5 10</intersection>
<intersection>-3088 9</intersection>
<intersection>-3069 8</intersection>
<intersection>-3050.5 7</intersection>
<intersection>-3028.5 6</intersection>
<intersection>-3010 5</intersection>
<intersection>-2991 4</intersection>
<intersection>-2972.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-2972.5,13.5,-2972.5</points>
<connection>
<GID>7895</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12.5,-2991,13.5,-2991</points>
<connection>
<GID>7859</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>12.5,-3010,13.5,-3010</points>
<connection>
<GID>7823</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>12.5,-3028.5,13.5,-3028.5</points>
<connection>
<GID>7763</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>12.5,-3050.5,13.5,-3050.5</points>
<connection>
<GID>7677</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>12.5,-3069,13.5,-3069</points>
<connection>
<GID>7641</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-3088,13.5,-3088</points>
<connection>
<GID>7604</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>12.5,-3106.5,13.5,-3106.5</points>
<connection>
<GID>7931</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-3128,22.5,-2963</points>
<connection>
<GID>7729</GID>
<name>N_in1</name></connection>
<connection>
<GID>7727</GID>
<name>N_in0</name></connection>
<intersection>-3116 3</intersection>
<intersection>-3097.5 5</intersection>
<intersection>-3078.5 7</intersection>
<intersection>-3060 9</intersection>
<intersection>-3038 11</intersection>
<intersection>-3019.5 13</intersection>
<intersection>-3000.5 15</intersection>
<intersection>-2982 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-3116,24.5,-3116</points>
<connection>
<GID>7933</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>22.5,-3097.5,24.5,-3097.5</points>
<connection>
<GID>7606</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22.5,-3078.5,24.5,-3078.5</points>
<connection>
<GID>7643</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22.5,-3060,24.5,-3060</points>
<connection>
<GID>7678</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>22.5,-3038,25,-3038</points>
<connection>
<GID>7768</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>22.5,-3019.5,25,-3019.5</points>
<connection>
<GID>7825</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>22.5,-3000.5,25,-3000.5</points>
<connection>
<GID>7861</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>22.5,-2982,25,-2982</points>
<connection>
<GID>7897</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3215.5,54,-3215.5</points>
<connection>
<GID>7828</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3215.5,48,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3200,48,-3200</points>
<connection>
<GID>7816</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5393</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3215.5,77,-3215.5</points>
<connection>
<GID>7854</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3215.5,71,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3200,71,-3200</points>
<connection>
<GID>7852</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3215.5,102,-3215.5</points>
<connection>
<GID>7862</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3215.5,96,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3200,96,-3200</points>
<connection>
<GID>7858</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5395</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3215.5,125,-3215.5</points>
<connection>
<GID>7870</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3215.5,119,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3200,119,-3200</points>
<connection>
<GID>7866</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3215.5,148,-3215.5</points>
<connection>
<GID>7876</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3215.5,142,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3200,142,-3200</points>
<connection>
<GID>7872</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3215.5,171,-3215.5</points>
<connection>
<GID>7880</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3215.5,165,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3200,165,-3200</points>
<connection>
<GID>7878</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5398</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3215.5,196,-3215.5</points>
<connection>
<GID>7884</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3215.5,190,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3200,190,-3200</points>
<connection>
<GID>7882</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3215.5,219,-3215.5</points>
<connection>
<GID>7888</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3215.5,213,-3200</points>
<intersection>-3215.5 1</intersection>
<intersection>-3200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3200,213,-3200</points>
<connection>
<GID>7886</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5400</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3203,206,-3203</points>
<connection>
<GID>7886</GID>
<name>clock</name></connection>
<connection>
<GID>7882</GID>
<name>clock</name></connection>
<connection>
<GID>7878</GID>
<name>clock</name></connection>
<connection>
<GID>7872</GID>
<name>clock</name></connection>
<connection>
<GID>7866</GID>
<name>clock</name></connection>
<connection>
<GID>7858</GID>
<name>clock</name></connection>
<connection>
<GID>7852</GID>
<name>clock</name></connection>
<connection>
<GID>7816</GID>
<name>clock</name></connection>
<connection>
<GID>7810</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3212.5,217,-3212.5</points>
<connection>
<GID>7888</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7884</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7880</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7876</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7870</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7862</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7854</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7828</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7812</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3197,54,-3197</points>
<connection>
<GID>7896</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3197,48,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3181.5,48,-3181.5</points>
<connection>
<GID>7894</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3197,77,-3197</points>
<connection>
<GID>7900</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3197,71,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3181.5,71,-3181.5</points>
<connection>
<GID>7898</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5404</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3197,102,-3197</points>
<connection>
<GID>7904</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3197,96,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3181.5,96,-3181.5</points>
<connection>
<GID>7902</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3197,125,-3197</points>
<connection>
<GID>7908</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3197,119,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3181.5,119,-3181.5</points>
<connection>
<GID>7906</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3197,148,-3197</points>
<connection>
<GID>7912</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3197,142,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3181.5,142,-3181.5</points>
<connection>
<GID>7910</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5407</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3197,171,-3197</points>
<connection>
<GID>7916</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3197,165,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3181.5,165,-3181.5</points>
<connection>
<GID>7914</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5408</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3197,196,-3197</points>
<connection>
<GID>7920</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3197,190,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3181.5,190,-3181.5</points>
<connection>
<GID>7918</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3197,219,-3197</points>
<connection>
<GID>7924</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3197,213,-3181.5</points>
<intersection>-3197 1</intersection>
<intersection>-3181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3181.5,213,-3181.5</points>
<connection>
<GID>7922</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5410</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3184.5,206,-3184.5</points>
<connection>
<GID>7922</GID>
<name>clock</name></connection>
<connection>
<GID>7918</GID>
<name>clock</name></connection>
<connection>
<GID>7914</GID>
<name>clock</name></connection>
<connection>
<GID>7910</GID>
<name>clock</name></connection>
<connection>
<GID>7906</GID>
<name>clock</name></connection>
<connection>
<GID>7902</GID>
<name>clock</name></connection>
<connection>
<GID>7898</GID>
<name>clock</name></connection>
<connection>
<GID>7894</GID>
<name>clock</name></connection>
<connection>
<GID>7890</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3194,217,-3194</points>
<connection>
<GID>7924</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7920</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7916</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7912</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7908</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7904</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7900</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7896</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7892</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3178,54,-3178</points>
<connection>
<GID>7932</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3178,48,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3162.5,48,-3162.5</points>
<connection>
<GID>7930</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3178,77,-3178</points>
<connection>
<GID>7936</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3178,71,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3162.5,71,-3162.5</points>
<connection>
<GID>7934</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3178,102,-3178</points>
<connection>
<GID>7940</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3178,96,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3162.5,96,-3162.5</points>
<connection>
<GID>7938</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3178,125,-3178</points>
<connection>
<GID>7944</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3178,119,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3162.5,119,-3162.5</points>
<connection>
<GID>7942</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3178,148,-3178</points>
<connection>
<GID>7585</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3178,142,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3162.5,142,-3162.5</points>
<connection>
<GID>7946</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3178,171,-3178</points>
<connection>
<GID>7589</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3178,165,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3162.5,165,-3162.5</points>
<connection>
<GID>7587</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5418</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3178,196,-3178</points>
<connection>
<GID>7593</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3178,190,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3162.5,190,-3162.5</points>
<connection>
<GID>7591</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3178,219,-3178</points>
<connection>
<GID>7597</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3178,213,-3162.5</points>
<intersection>-3178 1</intersection>
<intersection>-3162.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3162.5,213,-3162.5</points>
<connection>
<GID>7595</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3165.5,206,-3165.5</points>
<connection>
<GID>7946</GID>
<name>clock</name></connection>
<connection>
<GID>7942</GID>
<name>clock</name></connection>
<connection>
<GID>7938</GID>
<name>clock</name></connection>
<connection>
<GID>7934</GID>
<name>clock</name></connection>
<connection>
<GID>7930</GID>
<name>clock</name></connection>
<connection>
<GID>7926</GID>
<name>OUT</name></connection>
<connection>
<GID>7595</GID>
<name>clock</name></connection>
<connection>
<GID>7591</GID>
<name>clock</name></connection>
<connection>
<GID>7587</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3175,217,-3175</points>
<connection>
<GID>7944</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7940</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7936</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7932</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7928</GID>
<name>OUT</name></connection>
<connection>
<GID>7597</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7593</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7589</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7585</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3159.5,54,-3159.5</points>
<connection>
<GID>7605</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3159.5,48,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3144,48,-3144</points>
<connection>
<GID>7603</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3159.5,77,-3159.5</points>
<connection>
<GID>7609</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3159.5,71,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3144,71,-3144</points>
<connection>
<GID>7607</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3159.5,102,-3159.5</points>
<connection>
<GID>7613</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3159.5,96,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3144,96,-3144</points>
<connection>
<GID>7611</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3159.5,125,-3159.5</points>
<connection>
<GID>7617</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3159.5,119,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3144,119,-3144</points>
<connection>
<GID>7615</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3159.5,148,-3159.5</points>
<connection>
<GID>7621</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3159.5,142,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3144,142,-3144</points>
<connection>
<GID>7619</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3159.5,171,-3159.5</points>
<connection>
<GID>7625</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3159.5,165,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3144,165,-3144</points>
<connection>
<GID>7623</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3159.5,196,-3159.5</points>
<connection>
<GID>7629</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3159.5,190,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3144,190,-3144</points>
<connection>
<GID>7627</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5429</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3159.5,219,-3159.5</points>
<connection>
<GID>7633</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3159.5,213,-3144</points>
<intersection>-3159.5 1</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3144,213,-3144</points>
<connection>
<GID>7631</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3147,206,-3147</points>
<connection>
<GID>7631</GID>
<name>clock</name></connection>
<connection>
<GID>7627</GID>
<name>clock</name></connection>
<connection>
<GID>7623</GID>
<name>clock</name></connection>
<connection>
<GID>7619</GID>
<name>clock</name></connection>
<connection>
<GID>7615</GID>
<name>clock</name></connection>
<connection>
<GID>7611</GID>
<name>clock</name></connection>
<connection>
<GID>7607</GID>
<name>clock</name></connection>
<connection>
<GID>7603</GID>
<name>clock</name></connection>
<connection>
<GID>7599</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5431</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3156.5,217,-3156.5</points>
<connection>
<GID>7633</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7629</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7625</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7621</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7617</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7613</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7609</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7605</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7601</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5432</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3293.5,54,-3293.5</points>
<connection>
<GID>7642</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3293.5,48,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3278,48,-3278</points>
<connection>
<GID>7639</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5433</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3293.5,77,-3293.5</points>
<connection>
<GID>7647</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3293.5,71,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3278,71,-3278</points>
<connection>
<GID>7644</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3293.5,102,-3293.5</points>
<connection>
<GID>7652</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3293.5,96,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3278,96,-3278</points>
<connection>
<GID>7649</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3293.5,125,-3293.5</points>
<connection>
<GID>7657</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3293.5,119,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3278,119,-3278</points>
<connection>
<GID>7654</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3293.5,148,-3293.5</points>
<connection>
<GID>7662</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3293.5,142,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3278,142,-3278</points>
<connection>
<GID>7659</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5437</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3293.5,171,-3293.5</points>
<connection>
<GID>7667</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3293.5,165,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3278,165,-3278</points>
<connection>
<GID>7664</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3293.5,196,-3293.5</points>
<connection>
<GID>7734</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3293.5,190,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3278,190,-3278</points>
<connection>
<GID>7733</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5439</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3293.5,219,-3293.5</points>
<connection>
<GID>7736</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3293.5,213,-3278</points>
<intersection>-3293.5 1</intersection>
<intersection>-3278 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3278,213,-3278</points>
<connection>
<GID>7735</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5440</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3281,206,-3281</points>
<connection>
<GID>7735</GID>
<name>clock</name></connection>
<connection>
<GID>7733</GID>
<name>clock</name></connection>
<connection>
<GID>7664</GID>
<name>clock</name></connection>
<connection>
<GID>7659</GID>
<name>clock</name></connection>
<connection>
<GID>7654</GID>
<name>clock</name></connection>
<connection>
<GID>7649</GID>
<name>clock</name></connection>
<connection>
<GID>7644</GID>
<name>clock</name></connection>
<connection>
<GID>7639</GID>
<name>clock</name></connection>
<connection>
<GID>7635</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5441</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3290.5,217,-3290.5</points>
<connection>
<GID>7736</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7734</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7667</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7662</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7657</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7652</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7647</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7642</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7637</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5442</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3275,54,-3275</points>
<connection>
<GID>7740</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3275,48,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3259.5,48,-3259.5</points>
<connection>
<GID>7739</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3275,77,-3275</points>
<connection>
<GID>7742</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3275,71,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3259.5,71,-3259.5</points>
<connection>
<GID>7741</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5444</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3275,102,-3275</points>
<connection>
<GID>7744</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3275,96,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3259.5,96,-3259.5</points>
<connection>
<GID>7743</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5445</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3275,125,-3275</points>
<connection>
<GID>7746</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3275,119,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3259.5,119,-3259.5</points>
<connection>
<GID>7745</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3275,148,-3275</points>
<connection>
<GID>7748</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3275,142,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3259.5,142,-3259.5</points>
<connection>
<GID>7747</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5447</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3275,171,-3275</points>
<connection>
<GID>7750</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3275,165,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3259.5,165,-3259.5</points>
<connection>
<GID>7749</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5448</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3275,196,-3275</points>
<connection>
<GID>7752</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3275,190,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3259.5,190,-3259.5</points>
<connection>
<GID>7751</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3275,219,-3275</points>
<connection>
<GID>7754</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3275,213,-3259.5</points>
<intersection>-3275 1</intersection>
<intersection>-3259.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3259.5,213,-3259.5</points>
<connection>
<GID>7753</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3262.5,206,-3262.5</points>
<connection>
<GID>7753</GID>
<name>clock</name></connection>
<connection>
<GID>7751</GID>
<name>clock</name></connection>
<connection>
<GID>7749</GID>
<name>clock</name></connection>
<connection>
<GID>7747</GID>
<name>clock</name></connection>
<connection>
<GID>7745</GID>
<name>clock</name></connection>
<connection>
<GID>7743</GID>
<name>clock</name></connection>
<connection>
<GID>7741</GID>
<name>clock</name></connection>
<connection>
<GID>7739</GID>
<name>clock</name></connection>
<connection>
<GID>7737</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3272,217,-3272</points>
<connection>
<GID>7754</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7752</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7748</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7746</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7744</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7742</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7740</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7738</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3256,54,-3256</points>
<connection>
<GID>7650</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3256,48,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3240.5,48,-3240.5</points>
<connection>
<GID>7645</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5453</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3256,77,-3256</points>
<connection>
<GID>7660</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3256,71,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3240.5,71,-3240.5</points>
<connection>
<GID>7655</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3256,102,-3256</points>
<connection>
<GID>7669</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3256,96,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3240.5,96,-3240.5</points>
<connection>
<GID>7665</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3256,125,-3256</points>
<connection>
<GID>7756</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3256,119,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3240.5,119,-3240.5</points>
<connection>
<GID>7672</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3256,148,-3256</points>
<connection>
<GID>7758</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3256,142,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3240.5,142,-3240.5</points>
<connection>
<GID>7757</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5457</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3256,171,-3256</points>
<connection>
<GID>7760</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3256,165,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3240.5,165,-3240.5</points>
<connection>
<GID>7759</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3256,196,-3256</points>
<connection>
<GID>7762</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3256,190,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3240.5,190,-3240.5</points>
<connection>
<GID>7761</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3256,219,-3256</points>
<connection>
<GID>7765</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3256,213,-3240.5</points>
<intersection>-3256 1</intersection>
<intersection>-3240.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3240.5,213,-3240.5</points>
<connection>
<GID>7764</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3243.5,206,-3243.5</points>
<connection>
<GID>7764</GID>
<name>clock</name></connection>
<connection>
<GID>7761</GID>
<name>clock</name></connection>
<connection>
<GID>7759</GID>
<name>clock</name></connection>
<connection>
<GID>7757</GID>
<name>clock</name></connection>
<connection>
<GID>7755</GID>
<name>OUT</name></connection>
<connection>
<GID>7672</GID>
<name>clock</name></connection>
<connection>
<GID>7665</GID>
<name>clock</name></connection>
<connection>
<GID>7655</GID>
<name>clock</name></connection>
<connection>
<GID>7645</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3253,217,-3253</points>
<connection>
<GID>7765</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7762</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7760</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7758</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7756</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7669</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7660</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7650</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7640</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3237.5,54,-3237.5</points>
<connection>
<GID>7770</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3237.5,48,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3222,48,-3222</points>
<connection>
<GID>7769</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5463</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3237.5,77,-3237.5</points>
<connection>
<GID>7772</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3237.5,71,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3222,71,-3222</points>
<connection>
<GID>7771</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3237.5,102,-3237.5</points>
<connection>
<GID>7775</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3237.5,96,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3222,96,-3222</points>
<connection>
<GID>7774</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5465</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3237.5,125,-3237.5</points>
<connection>
<GID>7777</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3237.5,119,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3222,119,-3222</points>
<connection>
<GID>7776</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3237.5,148,-3237.5</points>
<connection>
<GID>7780</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3237.5,142,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3222,142,-3222</points>
<connection>
<GID>7778</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5467</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3237.5,171,-3237.5</points>
<connection>
<GID>7782</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3237.5,165,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3222,165,-3222</points>
<connection>
<GID>7781</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5468</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3237.5,196,-3237.5</points>
<connection>
<GID>7784</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3237.5,190,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3222,190,-3222</points>
<connection>
<GID>7783</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5469</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3237.5,219,-3237.5</points>
<connection>
<GID>7786</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3237.5,213,-3222</points>
<intersection>-3237.5 1</intersection>
<intersection>-3222 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3222,213,-3222</points>
<connection>
<GID>7785</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3225,206,-3225</points>
<connection>
<GID>7785</GID>
<name>clock</name></connection>
<connection>
<GID>7783</GID>
<name>clock</name></connection>
<connection>
<GID>7781</GID>
<name>clock</name></connection>
<connection>
<GID>7778</GID>
<name>clock</name></connection>
<connection>
<GID>7776</GID>
<name>clock</name></connection>
<connection>
<GID>7774</GID>
<name>clock</name></connection>
<connection>
<GID>7771</GID>
<name>clock</name></connection>
<connection>
<GID>7769</GID>
<name>clock</name></connection>
<connection>
<GID>7766</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5471</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3234.5,217,-3234.5</points>
<connection>
<GID>7786</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7784</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7782</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7780</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7777</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7775</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7772</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7770</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7767</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-3303.5,35.5,-3138.5</points>
<connection>
<GID>7814</GID>
<name>N_in1</name></connection>
<connection>
<GID>7787</GID>
<name>N_in0</name></connection>
<intersection>-3278 12</intersection>
<intersection>-3259.5 11</intersection>
<intersection>-3240.5 10</intersection>
<intersection>-3222 9</intersection>
<intersection>-3200 8</intersection>
<intersection>-3181.5 7</intersection>
<intersection>-3162.5 6</intersection>
<intersection>-3144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-3144,41,-3144</points>
<connection>
<GID>7603</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-3162.5,41,-3162.5</points>
<connection>
<GID>7930</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-3181.5,41,-3181.5</points>
<connection>
<GID>7894</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-3200,41,-3200</points>
<connection>
<GID>7816</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>35.5,-3222,41,-3222</points>
<connection>
<GID>7769</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>35.5,-3240.5,41,-3240.5</points>
<connection>
<GID>7645</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>35.5,-3259.5,41,-3259.5</points>
<connection>
<GID>7739</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>35.5,-3278,41,-3278</points>
<connection>
<GID>7639</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-3303,58.5,-3138</points>
<connection>
<GID>7818</GID>
<name>N_in1</name></connection>
<connection>
<GID>7788</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 4</intersection>
<intersection>-3267 5</intersection>
<intersection>-3248 6</intersection>
<intersection>-3229.5 7</intersection>
<intersection>-3207.5 8</intersection>
<intersection>-3189 9</intersection>
<intersection>-3170 10</intersection>
<intersection>-3151.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-3285.5,58.5,-3285.5</points>
<intersection>54 12</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54,-3267,58.5,-3267</points>
<intersection>54 14</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54,-3248,58.5,-3248</points>
<intersection>54 13</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54,-3229.5,58.5,-3229.5</points>
<intersection>54 15</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-3207.5,58.5,-3207.5</points>
<intersection>54 18</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>54,-3189,58.5,-3189</points>
<intersection>54 19</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>54,-3170,58.5,-3170</points>
<intersection>54 20</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>54,-3151.5,58.5,-3151.5</points>
<intersection>54 21</intersection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>54,-3288,54,-3285.5</points>
<connection>
<GID>7642</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>54,-3250.5,54,-3248</points>
<connection>
<GID>7650</GID>
<name>OUT_0</name></connection>
<intersection>-3248 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>54,-3269.5,54,-3267</points>
<connection>
<GID>7740</GID>
<name>OUT_0</name></connection>
<intersection>-3267 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>54,-3232,54,-3229.5</points>
<connection>
<GID>7770</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>54,-3210,54,-3207.5</points>
<connection>
<GID>7828</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>54,-3191.5,54,-3189</points>
<connection>
<GID>7896</GID>
<name>OUT_0</name></connection>
<intersection>-3189 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>54,-3172.5,54,-3170</points>
<connection>
<GID>7932</GID>
<name>OUT_0</name></connection>
<intersection>-3170 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>54,-3154,54,-3151.5</points>
<connection>
<GID>7605</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-3303,61.5,-3138.5</points>
<connection>
<GID>7820</GID>
<name>N_in1</name></connection>
<connection>
<GID>7789</GID>
<name>N_in0</name></connection>
<intersection>-3278 10</intersection>
<intersection>-3259.5 9</intersection>
<intersection>-3240.5 8</intersection>
<intersection>-3222 7</intersection>
<intersection>-3200 6</intersection>
<intersection>-3181.5 5</intersection>
<intersection>-3162.5 4</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-3144,64,-3144</points>
<connection>
<GID>7607</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-3162.5,64,-3162.5</points>
<connection>
<GID>7934</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61.5,-3181.5,64,-3181.5</points>
<connection>
<GID>7898</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61.5,-3200,64,-3200</points>
<connection>
<GID>7852</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61.5,-3222,64,-3222</points>
<connection>
<GID>7771</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61.5,-3240.5,64,-3240.5</points>
<connection>
<GID>7655</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61.5,-3259.5,64,-3259.5</points>
<connection>
<GID>7741</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61.5,-3278,64,-3278</points>
<connection>
<GID>7644</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-3303,81,-3138</points>
<connection>
<GID>7822</GID>
<name>N_in1</name></connection>
<connection>
<GID>7790</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 6</intersection>
<intersection>-3267 7</intersection>
<intersection>-3248 8</intersection>
<intersection>-3229.5 9</intersection>
<intersection>-3207.5 10</intersection>
<intersection>-3189 11</intersection>
<intersection>-3170 12</intersection>
<intersection>-3151.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-3285.5,81,-3285.5</points>
<intersection>77 14</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>77,-3267,81,-3267</points>
<intersection>77 16</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>77,-3248,81,-3248</points>
<intersection>77 15</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-3229.5,81,-3229.5</points>
<intersection>77 17</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>77,-3207.5,81,-3207.5</points>
<intersection>77 20</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>77,-3189,81,-3189</points>
<intersection>77 21</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>77,-3170,81,-3170</points>
<intersection>77 22</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>77,-3151.5,81,-3151.5</points>
<intersection>77 23</intersection>
<intersection>81 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>77,-3288,77,-3285.5</points>
<connection>
<GID>7647</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>77,-3250.5,77,-3248</points>
<connection>
<GID>7660</GID>
<name>OUT_0</name></connection>
<intersection>-3248 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>77,-3269.5,77,-3267</points>
<connection>
<GID>7742</GID>
<name>OUT_0</name></connection>
<intersection>-3267 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>77,-3232,77,-3229.5</points>
<connection>
<GID>7772</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>77,-3210,77,-3207.5</points>
<connection>
<GID>7854</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>77,-3191.5,77,-3189</points>
<connection>
<GID>7900</GID>
<name>OUT_0</name></connection>
<intersection>-3189 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>77,-3172.5,77,-3170</points>
<connection>
<GID>7936</GID>
<name>OUT_0</name></connection>
<intersection>-3170 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>77,-3154,77,-3151.5</points>
<connection>
<GID>7609</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-3303,84.5,-3138</points>
<connection>
<GID>7824</GID>
<name>N_in1</name></connection>
<connection>
<GID>7791</GID>
<name>N_in0</name></connection>
<intersection>-3278 13</intersection>
<intersection>-3259.5 12</intersection>
<intersection>-3240.5 11</intersection>
<intersection>-3222 10</intersection>
<intersection>-3200 9</intersection>
<intersection>-3181.5 8</intersection>
<intersection>-3162.5 7</intersection>
<intersection>-3144 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-3144,89,-3144</points>
<connection>
<GID>7611</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-3162.5,89,-3162.5</points>
<connection>
<GID>7938</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>84.5,-3181.5,89,-3181.5</points>
<connection>
<GID>7902</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84.5,-3200,89,-3200</points>
<connection>
<GID>7858</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84.5,-3222,89,-3222</points>
<connection>
<GID>7774</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84.5,-3240.5,89,-3240.5</points>
<connection>
<GID>7665</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>84.5,-3259.5,89,-3259.5</points>
<connection>
<GID>7743</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>84.5,-3278,89,-3278</points>
<connection>
<GID>7649</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3303,105.5,-3138.5</points>
<connection>
<GID>7826</GID>
<name>N_in1</name></connection>
<connection>
<GID>7792</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 6</intersection>
<intersection>-3267 7</intersection>
<intersection>-3248 8</intersection>
<intersection>-3229.5 9</intersection>
<intersection>-3207.5 10</intersection>
<intersection>-3189 11</intersection>
<intersection>-3170 12</intersection>
<intersection>-3151.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>102,-3285.5,105.5,-3285.5</points>
<intersection>102 14</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>102,-3267,105.5,-3267</points>
<intersection>102 16</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>102,-3248,105.5,-3248</points>
<intersection>102 15</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>102,-3229.5,105.5,-3229.5</points>
<intersection>102 17</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>102,-3207.5,105.5,-3207.5</points>
<intersection>102 20</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>102,-3189,105.5,-3189</points>
<intersection>102 21</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>102,-3170,105.5,-3170</points>
<intersection>102 22</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>102,-3151.5,105.5,-3151.5</points>
<intersection>102 23</intersection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>102,-3288,102,-3285.5</points>
<connection>
<GID>7652</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>102,-3250.5,102,-3248</points>
<connection>
<GID>7669</GID>
<name>OUT_0</name></connection>
<intersection>-3248 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>102,-3269.5,102,-3267</points>
<connection>
<GID>7744</GID>
<name>OUT_0</name></connection>
<intersection>-3267 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>102,-3232,102,-3229.5</points>
<connection>
<GID>7775</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>102,-3210,102,-3207.5</points>
<connection>
<GID>7862</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>102,-3191.5,102,-3189</points>
<connection>
<GID>7904</GID>
<name>OUT_0</name></connection>
<intersection>-3189 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>102,-3172.5,102,-3170</points>
<connection>
<GID>7940</GID>
<name>OUT_0</name></connection>
<intersection>-3170 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>102,-3154,102,-3151.5</points>
<connection>
<GID>7613</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3303,109.5,-3138</points>
<connection>
<GID>7830</GID>
<name>N_in1</name></connection>
<connection>
<GID>7793</GID>
<name>N_in0</name></connection>
<intersection>-3278 13</intersection>
<intersection>-3259.5 12</intersection>
<intersection>-3240.5 11</intersection>
<intersection>-3222 10</intersection>
<intersection>-3200 9</intersection>
<intersection>-3181.5 8</intersection>
<intersection>-3162.5 7</intersection>
<intersection>-3144 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109.5,-3144,112,-3144</points>
<connection>
<GID>7615</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>109.5,-3162.5,112,-3162.5</points>
<connection>
<GID>7942</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109.5,-3181.5,112,-3181.5</points>
<connection>
<GID>7906</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>109.5,-3200,112,-3200</points>
<connection>
<GID>7866</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>109.5,-3222,112,-3222</points>
<connection>
<GID>7776</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>109.5,-3240.5,112,-3240.5</points>
<connection>
<GID>7672</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109.5,-3259.5,112,-3259.5</points>
<connection>
<GID>7745</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>109.5,-3278,112,-3278</points>
<connection>
<GID>7654</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-3303,128,-3138</points>
<connection>
<GID>7832</GID>
<name>N_in1</name></connection>
<connection>
<GID>7794</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 6</intersection>
<intersection>-3267 7</intersection>
<intersection>-3248 8</intersection>
<intersection>-3229.5 9</intersection>
<intersection>-3207.5 10</intersection>
<intersection>-3189 11</intersection>
<intersection>-3170 12</intersection>
<intersection>-3151.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>125,-3285.5,128,-3285.5</points>
<intersection>125 14</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125,-3267,128,-3267</points>
<intersection>125 15</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>125,-3248,128,-3248</points>
<intersection>125 16</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>125,-3229.5,128,-3229.5</points>
<intersection>125 17</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125,-3207.5,128,-3207.5</points>
<intersection>125 20</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>125,-3189,128,-3189</points>
<intersection>125 21</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>125,-3170,128,-3170</points>
<intersection>125 22</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>125,-3151.5,128,-3151.5</points>
<intersection>125 23</intersection>
<intersection>128 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>125,-3288,125,-3285.5</points>
<connection>
<GID>7657</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>125,-3269.5,125,-3267</points>
<connection>
<GID>7746</GID>
<name>OUT_0</name></connection>
<intersection>-3267 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>125,-3250.5,125,-3248</points>
<connection>
<GID>7756</GID>
<name>OUT_0</name></connection>
<intersection>-3248 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>125,-3232,125,-3229.5</points>
<connection>
<GID>7777</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>125,-3210,125,-3207.5</points>
<connection>
<GID>7870</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>125,-3191.5,125,-3189</points>
<connection>
<GID>7908</GID>
<name>OUT_0</name></connection>
<intersection>-3189 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>125,-3172.5,125,-3170</points>
<connection>
<GID>7944</GID>
<name>OUT_0</name></connection>
<intersection>-3170 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>125,-3154,125,-3151.5</points>
<connection>
<GID>7617</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-3303,132,-3138</points>
<connection>
<GID>7834</GID>
<name>N_in1</name></connection>
<connection>
<GID>7796</GID>
<name>N_in0</name></connection>
<intersection>-3278 13</intersection>
<intersection>-3259.5 12</intersection>
<intersection>-3240.5 11</intersection>
<intersection>-3222 10</intersection>
<intersection>-3200 9</intersection>
<intersection>-3181.5 8</intersection>
<intersection>-3162.5 7</intersection>
<intersection>-3144 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>132,-3144,135,-3144</points>
<connection>
<GID>7619</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>132,-3162.5,135,-3162.5</points>
<connection>
<GID>7946</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>132,-3181.5,135,-3181.5</points>
<connection>
<GID>7910</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>132,-3200,135,-3200</points>
<connection>
<GID>7872</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132,-3222,135,-3222</points>
<connection>
<GID>7778</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132,-3240.5,135,-3240.5</points>
<connection>
<GID>7757</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>132,-3259.5,135,-3259.5</points>
<connection>
<GID>7747</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132,-3278,135,-3278</points>
<connection>
<GID>7659</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>5481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-3302.5,151,-3138</points>
<connection>
<GID>7836</GID>
<name>N_in1</name></connection>
<connection>
<GID>7798</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 6</intersection>
<intersection>-3267 7</intersection>
<intersection>-3248 8</intersection>
<intersection>-3229.5 9</intersection>
<intersection>-3207.5 10</intersection>
<intersection>-3189 11</intersection>
<intersection>-3170 12</intersection>
<intersection>-3151.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>148,-3285.5,151,-3285.5</points>
<intersection>148 15</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>148,-3267,151,-3267</points>
<intersection>148 16</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>148,-3248,151,-3248</points>
<intersection>148 17</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>148,-3229.5,151,-3229.5</points>
<intersection>148 18</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>148,-3207.5,151,-3207.5</points>
<intersection>148 21</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>148,-3189,151,-3189</points>
<intersection>148 22</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>148,-3170,151,-3170</points>
<intersection>148 23</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>148,-3151.5,151,-3151.5</points>
<intersection>148 14</intersection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>148,-3154,148,-3151.5</points>
<connection>
<GID>7621</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>148,-3288,148,-3285.5</points>
<connection>
<GID>7662</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>148,-3269.5,148,-3267</points>
<connection>
<GID>7748</GID>
<name>OUT_0</name></connection>
<intersection>-3267 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>148,-3250.5,148,-3248</points>
<connection>
<GID>7758</GID>
<name>OUT_0</name></connection>
<intersection>-3248 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>148,-3232,148,-3229.5</points>
<connection>
<GID>7780</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>148,-3210,148,-3207.5</points>
<connection>
<GID>7876</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>148,-3191.5,148,-3189</points>
<connection>
<GID>7912</GID>
<name>OUT_0</name></connection>
<intersection>-3189 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>148,-3172.5,148,-3170</points>
<connection>
<GID>7585</GID>
<name>OUT_0</name></connection>
<intersection>-3170 12</intersection></vsegment></shape></wire>
<wire>
<ID>5482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-3302.5,156,-3138</points>
<connection>
<GID>7838</GID>
<name>N_in1</name></connection>
<connection>
<GID>7800</GID>
<name>N_in0</name></connection>
<intersection>-3278 13</intersection>
<intersection>-3259.5 12</intersection>
<intersection>-3240.5 11</intersection>
<intersection>-3222 10</intersection>
<intersection>-3200 9</intersection>
<intersection>-3181.5 8</intersection>
<intersection>-3162.5 7</intersection>
<intersection>-3144 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>156,-3144,158,-3144</points>
<connection>
<GID>7623</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>156,-3162.5,158,-3162.5</points>
<connection>
<GID>7587</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>156,-3181.5,158,-3181.5</points>
<connection>
<GID>7914</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>156,-3200,158,-3200</points>
<connection>
<GID>7878</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156,-3222,158,-3222</points>
<connection>
<GID>7781</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>156,-3240.5,158,-3240.5</points>
<connection>
<GID>7759</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>156,-3259.5,158,-3259.5</points>
<connection>
<GID>7749</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>156,-3278,158,-3278</points>
<connection>
<GID>7664</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>5483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-3302,174,-3138</points>
<connection>
<GID>7840</GID>
<name>N_in1</name></connection>
<connection>
<GID>7804</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 16</intersection>
<intersection>-3267 15</intersection>
<intersection>-3248 14</intersection>
<intersection>-3229.5 13</intersection>
<intersection>-3207.5 12</intersection>
<intersection>-3189 11</intersection>
<intersection>-3170 10</intersection>
<intersection>-3151.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>171,-3151.5,174,-3151.5</points>
<intersection>171 17</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>171,-3170,174,-3170</points>
<intersection>171 26</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>171,-3189,174,-3189</points>
<intersection>171 25</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>171,-3207.5,174,-3207.5</points>
<intersection>171 24</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>171,-3229.5,174,-3229.5</points>
<intersection>171 21</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>171,-3248,174,-3248</points>
<intersection>171 20</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>171,-3267,174,-3267</points>
<intersection>171 19</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>171,-3285.5,174,-3285.5</points>
<intersection>171 18</intersection>
<intersection>174 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>171,-3154,171,-3151.5</points>
<connection>
<GID>7625</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>171,-3288,171,-3285.5</points>
<connection>
<GID>7667</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>171,-3269.5,171,-3267</points>
<connection>
<GID>7750</GID>
<name>OUT_0</name></connection>
<intersection>-3267 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>171,-3250.5,171,-3248</points>
<connection>
<GID>7760</GID>
<name>OUT_0</name></connection>
<intersection>-3248 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>171,-3232,171,-3229.5</points>
<connection>
<GID>7782</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>171,-3210,171,-3207.5</points>
<connection>
<GID>7880</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>171,-3191.5,171,-3189</points>
<connection>
<GID>7916</GID>
<name>OUT_0</name></connection>
<intersection>-3189 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>171,-3172.5,171,-3170</points>
<connection>
<GID>7589</GID>
<name>OUT_0</name></connection>
<intersection>-3170 10</intersection></vsegment></shape></wire>
<wire>
<ID>5484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-3302,178.5,-3138</points>
<connection>
<GID>7842</GID>
<name>N_in1</name></connection>
<connection>
<GID>7802</GID>
<name>N_in0</name></connection>
<intersection>-3278 13</intersection>
<intersection>-3259.5 12</intersection>
<intersection>-3240.5 11</intersection>
<intersection>-3222 10</intersection>
<intersection>-3200 9</intersection>
<intersection>-3181.5 8</intersection>
<intersection>-3162.5 7</intersection>
<intersection>-3144 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>178.5,-3144,183,-3144</points>
<connection>
<GID>7627</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>178.5,-3162.5,183,-3162.5</points>
<connection>
<GID>7591</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178.5,-3181.5,183,-3181.5</points>
<connection>
<GID>7918</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>178.5,-3200,183,-3200</points>
<connection>
<GID>7882</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>178.5,-3222,183,-3222</points>
<connection>
<GID>7783</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>178.5,-3240.5,183,-3240.5</points>
<connection>
<GID>7761</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>178.5,-3259.5,183,-3259.5</points>
<connection>
<GID>7751</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>178.5,-3278,183,-3278</points>
<connection>
<GID>7733</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-3301.5,199.5,-3138.5</points>
<connection>
<GID>7844</GID>
<name>N_in1</name></connection>
<connection>
<GID>7806</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 6</intersection>
<intersection>-3267 7</intersection>
<intersection>-3248 8</intersection>
<intersection>-3229.5 9</intersection>
<intersection>-3207.5 10</intersection>
<intersection>-3189 11</intersection>
<intersection>-3170 12</intersection>
<intersection>-3151.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196,-3285.5,199.5,-3285.5</points>
<intersection>196 15</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>196,-3267,199.5,-3267</points>
<intersection>196 16</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>196,-3248,199.5,-3248</points>
<intersection>196 17</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>196,-3229.5,199.5,-3229.5</points>
<intersection>196 18</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>196,-3207.5,199.5,-3207.5</points>
<intersection>196 21</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>196,-3189,199.5,-3189</points>
<intersection>196 22</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>196,-3170,199.5,-3170</points>
<intersection>196 23</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>196,-3151.5,199.5,-3151.5</points>
<intersection>196 14</intersection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>196,-3154,196,-3151.5</points>
<connection>
<GID>7629</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>196,-3288,196,-3285.5</points>
<connection>
<GID>7734</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>196,-3269.5,196,-3267</points>
<connection>
<GID>7752</GID>
<name>OUT_0</name></connection>
<intersection>-3267 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>196,-3250.5,196,-3248</points>
<connection>
<GID>7762</GID>
<name>OUT_0</name></connection>
<intersection>-3248 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>196,-3232,196,-3229.5</points>
<connection>
<GID>7784</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>196,-3210,196,-3207.5</points>
<connection>
<GID>7884</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>196,-3191.5,196,-3189</points>
<connection>
<GID>7920</GID>
<name>OUT_0</name></connection>
<intersection>-3189 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>196,-3172.5,196,-3170</points>
<connection>
<GID>7593</GID>
<name>OUT_0</name></connection>
<intersection>-3170 12</intersection></vsegment></shape></wire>
<wire>
<ID>5486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-3301.5,203,-3138.5</points>
<connection>
<GID>7846</GID>
<name>N_in1</name></connection>
<connection>
<GID>7848</GID>
<name>N_in0</name></connection>
<intersection>-3278 11</intersection>
<intersection>-3259.5 10</intersection>
<intersection>-3240.5 9</intersection>
<intersection>-3222 7</intersection>
<intersection>-3200 6</intersection>
<intersection>-3181.5 5</intersection>
<intersection>-3162.5 4</intersection>
<intersection>-3144 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-3144,206,-3144</points>
<connection>
<GID>7631</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>203,-3162.5,206,-3162.5</points>
<connection>
<GID>7595</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>203,-3181.5,206,-3181.5</points>
<connection>
<GID>7922</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>203,-3200,206,-3200</points>
<connection>
<GID>7886</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-3222,206,-3222</points>
<connection>
<GID>7785</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>203,-3240.5,206,-3240.5</points>
<connection>
<GID>7764</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>203,-3259.5,206,-3259.5</points>
<connection>
<GID>7753</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-3278,206,-3278</points>
<connection>
<GID>7735</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment></shape></wire>
<wire>
<ID>5487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-3301.5,224,-3139.5</points>
<connection>
<GID>7850</GID>
<name>N_in1</name></connection>
<connection>
<GID>7808</GID>
<name>N_in0</name></connection>
<intersection>-3285.5 11</intersection>
<intersection>-3267 10</intersection>
<intersection>-3248 9</intersection>
<intersection>-3229.5 8</intersection>
<intersection>-3207.5 7</intersection>
<intersection>-3189 6</intersection>
<intersection>-3170 5</intersection>
<intersection>-3151.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>219,-3151.5,224,-3151.5</points>
<intersection>219 12</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>219,-3170,224,-3170</points>
<intersection>219 21</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>219,-3189,224,-3189</points>
<intersection>219 20</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>219,-3207.5,224,-3207.5</points>
<intersection>219 19</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>219,-3229.5,224,-3229.5</points>
<intersection>219 16</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>219,-3248,224,-3248</points>
<intersection>219 15</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>219,-3267,224,-3267</points>
<intersection>219 14</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>219,-3285.5,224,-3285.5</points>
<intersection>219 13</intersection>
<intersection>224 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>219,-3154,219,-3151.5</points>
<connection>
<GID>7633</GID>
<name>OUT_0</name></connection>
<intersection>-3151.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>219,-3288,219,-3285.5</points>
<connection>
<GID>7736</GID>
<name>OUT_0</name></connection>
<intersection>-3285.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>219,-3269.5,219,-3267</points>
<connection>
<GID>7754</GID>
<name>OUT_0</name></connection>
<intersection>-3267 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>219,-3250.5,219,-3248</points>
<connection>
<GID>7765</GID>
<name>OUT_0</name></connection>
<intersection>-3248 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>219,-3232,219,-3229.5</points>
<connection>
<GID>7786</GID>
<name>OUT_0</name></connection>
<intersection>-3229.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>219,-3210,219,-3207.5</points>
<connection>
<GID>7888</GID>
<name>OUT_0</name></connection>
<intersection>-3207.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>219,-3191.5,219,-3189</points>
<connection>
<GID>7924</GID>
<name>OUT_0</name></connection>
<intersection>-3189 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>219,-3172.5,219,-3170</points>
<connection>
<GID>7597</GID>
<name>OUT_0</name></connection>
<intersection>-3170 5</intersection></vsegment></shape></wire>
<wire>
<ID>5488</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-126,-3146,13.5,-3146</points>
<connection>
<GID>7599</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-3155.5,-126,-3130</points>
<intersection>-3155.5 4</intersection>
<intersection>-3146 2</intersection>
<intersection>-3130 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-3155.5,25,-3155.5</points>
<connection>
<GID>7601</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3130,-126,-3130</points>
<connection>
<GID>7732</GID>
<name>OUT_7</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>5489</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-127,-3164.5,13.5,-3164.5</points>
<connection>
<GID>7926</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-127,-3174,-127,-3131</points>
<intersection>-3174 5</intersection>
<intersection>-3164.5 2</intersection>
<intersection>-3131 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-127,-3174,25,-3174</points>
<connection>
<GID>7928</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3131,-127,-3131</points>
<connection>
<GID>7732</GID>
<name>OUT_6</name></connection>
<intersection>-127 4</intersection></hsegment></shape></wire>
<wire>
<ID>5490</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-128,-3183.5,13.5,-3183.5</points>
<connection>
<GID>7890</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-3193,-128,-3132</points>
<intersection>-3193 4</intersection>
<intersection>-3183.5 2</intersection>
<intersection>-3132 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-3193,25,-3193</points>
<connection>
<GID>7892</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3132,-128,-3132</points>
<connection>
<GID>7732</GID>
<name>OUT_5</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>5491</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-129,-3202,13.5,-3202</points>
<connection>
<GID>7810</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-129,-3211.5,-129,-3133</points>
<intersection>-3211.5 4</intersection>
<intersection>-3202 2</intersection>
<intersection>-3133 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-129,-3211.5,25,-3211.5</points>
<connection>
<GID>7812</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3133,-129,-3133</points>
<connection>
<GID>7732</GID>
<name>OUT_4</name></connection>
<intersection>-129 3</intersection></hsegment></shape></wire>
<wire>
<ID>5492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-130,-3224,13.5,-3224</points>
<connection>
<GID>7766</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-130,-3233.5,-130,-3134</points>
<intersection>-3233.5 4</intersection>
<intersection>-3224 1</intersection>
<intersection>-3134 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-130,-3233.5,24.5,-3233.5</points>
<connection>
<GID>7767</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3134,-130,-3134</points>
<connection>
<GID>7732</GID>
<name>OUT_3</name></connection>
<intersection>-130 3</intersection></hsegment></shape></wire>
<wire>
<ID>5493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-131,-3242.5,13.5,-3242.5</points>
<connection>
<GID>7755</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-131,-3252,-131,-3135</points>
<intersection>-3252 4</intersection>
<intersection>-3242.5 1</intersection>
<intersection>-3135 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-131,-3252,24.5,-3252</points>
<connection>
<GID>7640</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3135,-131,-3135</points>
<connection>
<GID>7732</GID>
<name>OUT_2</name></connection>
<intersection>-131 3</intersection></hsegment></shape></wire>
<wire>
<ID>5494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-132,-3261.5,13.5,-3261.5</points>
<connection>
<GID>7737</GID>
<name>IN_0</name></connection>
<intersection>-132 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-132,-3271,-132,-3136</points>
<intersection>-3271 4</intersection>
<intersection>-3261.5 1</intersection>
<intersection>-3136 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-132,-3271,24.5,-3271</points>
<connection>
<GID>7738</GID>
<name>IN_0</name></connection>
<intersection>-132 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3136,-132,-3136</points>
<connection>
<GID>7732</GID>
<name>OUT_1</name></connection>
<intersection>-132 3</intersection></hsegment></shape></wire>
<wire>
<ID>5495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-133,-3280,13.5,-3280</points>
<connection>
<GID>7635</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-133,-3289.5,-133,-3137</points>
<connection>
<GID>7732</GID>
<name>OUT_0</name></connection>
<intersection>-3289.5 4</intersection>
<intersection>-3280 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-133,-3289.5,24.5,-3289.5</points>
<connection>
<GID>7637</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment></shape></wire>
<wire>
<ID>5496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-3303.5,12.5,-3138.5</points>
<connection>
<GID>7868</GID>
<name>N_in1</name></connection>
<connection>
<GID>7860</GID>
<name>N_in0</name></connection>
<intersection>-3282 10</intersection>
<intersection>-3263.5 9</intersection>
<intersection>-3244.5 8</intersection>
<intersection>-3226 7</intersection>
<intersection>-3204 6</intersection>
<intersection>-3185.5 5</intersection>
<intersection>-3166.5 4</intersection>
<intersection>-3148 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-3148,13.5,-3148</points>
<connection>
<GID>7599</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12.5,-3166.5,13.5,-3166.5</points>
<connection>
<GID>7926</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>12.5,-3185.5,13.5,-3185.5</points>
<connection>
<GID>7890</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>12.5,-3204,13.5,-3204</points>
<connection>
<GID>7810</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>12.5,-3226,13.5,-3226</points>
<connection>
<GID>7766</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>12.5,-3244.5,13.5,-3244.5</points>
<connection>
<GID>7755</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-3263.5,13.5,-3263.5</points>
<connection>
<GID>7737</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>12.5,-3282,13.5,-3282</points>
<connection>
<GID>7635</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-3303.5,22.5,-3138.5</points>
<connection>
<GID>7864</GID>
<name>N_in1</name></connection>
<connection>
<GID>7856</GID>
<name>N_in0</name></connection>
<intersection>-3291.5 3</intersection>
<intersection>-3273 5</intersection>
<intersection>-3254 7</intersection>
<intersection>-3235.5 9</intersection>
<intersection>-3213.5 11</intersection>
<intersection>-3195 13</intersection>
<intersection>-3176 15</intersection>
<intersection>-3157.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-3291.5,24.5,-3291.5</points>
<connection>
<GID>7637</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>22.5,-3273,24.5,-3273</points>
<connection>
<GID>7738</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22.5,-3254,24.5,-3254</points>
<connection>
<GID>7640</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22.5,-3235.5,24.5,-3235.5</points>
<connection>
<GID>7767</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>22.5,-3213.5,25,-3213.5</points>
<connection>
<GID>7812</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>22.5,-3195,25,-3195</points>
<connection>
<GID>7892</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>22.5,-3176,25,-3176</points>
<connection>
<GID>7928</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>22.5,-3157.5,25,-3157.5</points>
<connection>
<GID>7601</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-3136.5,12.5,-3130</points>
<connection>
<GID>7860</GID>
<name>N_in1</name></connection>
<connection>
<GID>7730</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-3136.5,22.5,-3130</points>
<connection>
<GID>7856</GID>
<name>N_in1</name></connection>
<connection>
<GID>7729</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-3136.5,35.5,-3130</points>
<connection>
<GID>7787</GID>
<name>N_in1</name></connection>
<connection>
<GID>7710</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-3136,58.5,-3129.5</points>
<connection>
<GID>7788</GID>
<name>N_in1</name></connection>
<connection>
<GID>7711</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-3136.5,61.5,-3129.5</points>
<connection>
<GID>7789</GID>
<name>N_in1</name></connection>
<connection>
<GID>7712</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-3136,81,-3129.5</points>
<connection>
<GID>7790</GID>
<name>N_in1</name></connection>
<connection>
<GID>7713</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-3136,84.5,-3129.5</points>
<connection>
<GID>7791</GID>
<name>N_in1</name></connection>
<connection>
<GID>7714</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3136.5,105.5,-3129.5</points>
<connection>
<GID>7792</GID>
<name>N_in1</name></connection>
<connection>
<GID>7715</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3136,109.5,-3129.5</points>
<connection>
<GID>7793</GID>
<name>N_in1</name></connection>
<connection>
<GID>7716</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-3136,128,-3129.5</points>
<connection>
<GID>7794</GID>
<name>N_in1</name></connection>
<connection>
<GID>7717</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-3136,132,-3129.5</points>
<connection>
<GID>7796</GID>
<name>N_in1</name></connection>
<connection>
<GID>7718</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-3136,151,-3129</points>
<connection>
<GID>7798</GID>
<name>N_in1</name></connection>
<connection>
<GID>7719</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-3136,156,-3129</points>
<connection>
<GID>7800</GID>
<name>N_in1</name></connection>
<connection>
<GID>7720</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-3136,174,-3128.5</points>
<connection>
<GID>7804</GID>
<name>N_in1</name></connection>
<connection>
<GID>7721</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-3136,178.5,-3128.5</points>
<connection>
<GID>7802</GID>
<name>N_in1</name></connection>
<connection>
<GID>7722</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-3136.5,199.5,-3128</points>
<connection>
<GID>7806</GID>
<name>N_in1</name></connection>
<connection>
<GID>7723</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-3136.5,203,-3128</points>
<connection>
<GID>7848</GID>
<name>N_in1</name></connection>
<connection>
<GID>7724</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-3137.5,224,-3128</points>
<connection>
<GID>7808</GID>
<name>N_in1</name></connection>
<connection>
<GID>7726</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3392,54,-3392</points>
<connection>
<GID>8144</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3392,48,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3376.5,48,-3376.5</points>
<connection>
<GID>8138</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3392,77,-3392</points>
<connection>
<GID>8162</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3392,71,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3376.5,71,-3376.5</points>
<connection>
<GID>8160</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3392,102,-3392</points>
<connection>
<GID>8166</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3392,96,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3376.5,96,-3376.5</points>
<connection>
<GID>8164</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5519</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3392,125,-3392</points>
<connection>
<GID>8170</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3392,119,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3376.5,119,-3376.5</points>
<connection>
<GID>8168</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3392,148,-3392</points>
<connection>
<GID>8174</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3392,142,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3376.5,142,-3376.5</points>
<connection>
<GID>8172</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3392,171,-3392</points>
<connection>
<GID>8178</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3392,165,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3376.5,165,-3376.5</points>
<connection>
<GID>8176</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3392,196,-3392</points>
<connection>
<GID>8182</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3392,190,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3376.5,190,-3376.5</points>
<connection>
<GID>8180</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3392,219,-3392</points>
<connection>
<GID>8186</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3392,213,-3376.5</points>
<intersection>-3392 1</intersection>
<intersection>-3376.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3376.5,213,-3376.5</points>
<connection>
<GID>8184</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3379.5,206,-3379.5</points>
<connection>
<GID>8128</GID>
<name>OUT</name></connection>
<connection>
<GID>8138</GID>
<name>clock</name></connection>
<connection>
<GID>8160</GID>
<name>clock</name></connection>
<connection>
<GID>8164</GID>
<name>clock</name></connection>
<connection>
<GID>8168</GID>
<name>clock</name></connection>
<connection>
<GID>8172</GID>
<name>clock</name></connection>
<connection>
<GID>8176</GID>
<name>clock</name></connection>
<connection>
<GID>8180</GID>
<name>clock</name></connection>
<connection>
<GID>8184</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3389,217,-3389</points>
<connection>
<GID>8133</GID>
<name>OUT</name></connection>
<connection>
<GID>8144</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8162</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8166</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8170</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8174</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8178</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8182</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8186</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3373.5,54,-3373.5</points>
<connection>
<GID>8194</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3373.5,48,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3358,48,-3358</points>
<connection>
<GID>8192</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3373.5,77,-3373.5</points>
<connection>
<GID>8198</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3373.5,71,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3358,71,-3358</points>
<connection>
<GID>8196</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3373.5,102,-3373.5</points>
<connection>
<GID>8202</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3373.5,96,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3358,96,-3358</points>
<connection>
<GID>8200</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3373.5,125,-3373.5</points>
<connection>
<GID>8206</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3373.5,119,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3358,119,-3358</points>
<connection>
<GID>8204</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3373.5,148,-3373.5</points>
<connection>
<GID>8210</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3373.5,142,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3358,142,-3358</points>
<connection>
<GID>8208</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3373.5,171,-3373.5</points>
<connection>
<GID>8214</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3373.5,165,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3358,165,-3358</points>
<connection>
<GID>8212</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3373.5,196,-3373.5</points>
<connection>
<GID>8218</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3373.5,190,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3358,190,-3358</points>
<connection>
<GID>8216</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3373.5,219,-3373.5</points>
<connection>
<GID>8222</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3373.5,213,-3358</points>
<intersection>-3373.5 1</intersection>
<intersection>-3358 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3358,213,-3358</points>
<connection>
<GID>8220</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3361,206,-3361</points>
<connection>
<GID>8188</GID>
<name>OUT</name></connection>
<connection>
<GID>8192</GID>
<name>clock</name></connection>
<connection>
<GID>8196</GID>
<name>clock</name></connection>
<connection>
<GID>8200</GID>
<name>clock</name></connection>
<connection>
<GID>8204</GID>
<name>clock</name></connection>
<connection>
<GID>8208</GID>
<name>clock</name></connection>
<connection>
<GID>8212</GID>
<name>clock</name></connection>
<connection>
<GID>8216</GID>
<name>clock</name></connection>
<connection>
<GID>8220</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3370.5,217,-3370.5</points>
<connection>
<GID>8190</GID>
<name>OUT</name></connection>
<connection>
<GID>8194</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8198</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8202</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8206</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8210</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8214</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8218</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8222</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3354.5,54,-3354.5</points>
<connection>
<GID>8230</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3354.5,48,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3339,48,-3339</points>
<connection>
<GID>8228</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3354.5,77,-3354.5</points>
<connection>
<GID>8234</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3354.5,71,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3339,71,-3339</points>
<connection>
<GID>8232</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5538</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3354.5,102,-3354.5</points>
<connection>
<GID>8238</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3354.5,96,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3339,96,-3339</points>
<connection>
<GID>8236</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3354.5,125,-3354.5</points>
<connection>
<GID>8242</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3354.5,119,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3339,119,-3339</points>
<connection>
<GID>8240</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5540</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3354.5,148,-3354.5</points>
<connection>
<GID>8246</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3354.5,142,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3339,142,-3339</points>
<connection>
<GID>8244</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5541</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3354.5,171,-3354.5</points>
<connection>
<GID>8250</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3354.5,165,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3339,165,-3339</points>
<connection>
<GID>8248</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5542</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3354.5,196,-3354.5</points>
<connection>
<GID>8254</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3354.5,190,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3339,190,-3339</points>
<connection>
<GID>8252</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5543</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3354.5,219,-3354.5</points>
<connection>
<GID>8258</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3354.5,213,-3339</points>
<intersection>-3354.5 1</intersection>
<intersection>-3339 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3339,213,-3339</points>
<connection>
<GID>8256</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5544</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3342,206,-3342</points>
<connection>
<GID>8224</GID>
<name>OUT</name></connection>
<connection>
<GID>8228</GID>
<name>clock</name></connection>
<connection>
<GID>8232</GID>
<name>clock</name></connection>
<connection>
<GID>8236</GID>
<name>clock</name></connection>
<connection>
<GID>8240</GID>
<name>clock</name></connection>
<connection>
<GID>8244</GID>
<name>clock</name></connection>
<connection>
<GID>8248</GID>
<name>clock</name></connection>
<connection>
<GID>8252</GID>
<name>clock</name></connection>
<connection>
<GID>8256</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5545</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3351.5,217,-3351.5</points>
<connection>
<GID>8226</GID>
<name>OUT</name></connection>
<connection>
<GID>8230</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8234</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8238</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8242</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8246</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8250</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8254</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8258</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3336,54,-3336</points>
<connection>
<GID>8266</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3336,48,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3320.5,48,-3320.5</points>
<connection>
<GID>8264</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5547</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3336,77,-3336</points>
<connection>
<GID>8270</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3336,71,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3320.5,71,-3320.5</points>
<connection>
<GID>8268</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3336,102,-3336</points>
<connection>
<GID>8274</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3336,96,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3320.5,96,-3320.5</points>
<connection>
<GID>8272</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3336,125,-3336</points>
<connection>
<GID>8278</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3336,119,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3320.5,119,-3320.5</points>
<connection>
<GID>8276</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3336,148,-3336</points>
<connection>
<GID>8282</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3336,142,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3320.5,142,-3320.5</points>
<connection>
<GID>8280</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5551</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3336,171,-3336</points>
<connection>
<GID>8286</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3336,165,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3320.5,165,-3320.5</points>
<connection>
<GID>8284</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5552</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3336,196,-3336</points>
<connection>
<GID>8290</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3336,190,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3320.5,190,-3320.5</points>
<connection>
<GID>8288</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5553</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3336,219,-3336</points>
<connection>
<GID>8294</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3336,213,-3320.5</points>
<intersection>-3336 1</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3320.5,213,-3320.5</points>
<connection>
<GID>8292</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5554</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3323.5,206,-3323.5</points>
<connection>
<GID>8260</GID>
<name>OUT</name></connection>
<connection>
<GID>8264</GID>
<name>clock</name></connection>
<connection>
<GID>8268</GID>
<name>clock</name></connection>
<connection>
<GID>8272</GID>
<name>clock</name></connection>
<connection>
<GID>8276</GID>
<name>clock</name></connection>
<connection>
<GID>8280</GID>
<name>clock</name></connection>
<connection>
<GID>8284</GID>
<name>clock</name></connection>
<connection>
<GID>8288</GID>
<name>clock</name></connection>
<connection>
<GID>8292</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3333,217,-3333</points>
<connection>
<GID>8262</GID>
<name>OUT</name></connection>
<connection>
<GID>8266</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8270</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8274</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8278</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8282</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8286</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8290</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8294</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3470,54,-3470</points>
<connection>
<GID>8302</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3470,48,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3454.5,48,-3454.5</points>
<connection>
<GID>8300</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3470,77,-3470</points>
<connection>
<GID>8306</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3470,71,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3454.5,71,-3454.5</points>
<connection>
<GID>8304</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5558</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3470,102,-3470</points>
<connection>
<GID>8310</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3470,96,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3454.5,96,-3454.5</points>
<connection>
<GID>8308</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5559</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3470,125,-3470</points>
<connection>
<GID>7951</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3470,119,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3454.5,119,-3454.5</points>
<connection>
<GID>7949</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5560</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3470,148,-3470</points>
<connection>
<GID>7955</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3470,142,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3454.5,142,-3454.5</points>
<connection>
<GID>7953</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3470,171,-3470</points>
<connection>
<GID>7959</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3470,165,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3454.5,165,-3454.5</points>
<connection>
<GID>7957</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5562</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3470,196,-3470</points>
<connection>
<GID>7963</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3470,190,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3454.5,190,-3454.5</points>
<connection>
<GID>7961</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5563</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3470,219,-3470</points>
<connection>
<GID>7967</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3470,213,-3454.5</points>
<intersection>-3470 1</intersection>
<intersection>-3454.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3454.5,213,-3454.5</points>
<connection>
<GID>7965</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3457.5,206,-3457.5</points>
<connection>
<GID>8308</GID>
<name>clock</name></connection>
<connection>
<GID>8304</GID>
<name>clock</name></connection>
<connection>
<GID>8300</GID>
<name>clock</name></connection>
<connection>
<GID>8296</GID>
<name>OUT</name></connection>
<connection>
<GID>7965</GID>
<name>clock</name></connection>
<connection>
<GID>7961</GID>
<name>clock</name></connection>
<connection>
<GID>7957</GID>
<name>clock</name></connection>
<connection>
<GID>7953</GID>
<name>clock</name></connection>
<connection>
<GID>7949</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3467,217,-3467</points>
<connection>
<GID>8310</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8306</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8302</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8298</GID>
<name>OUT</name></connection>
<connection>
<GID>7967</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7963</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7959</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7955</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7951</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5566</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3451.5,54,-3451.5</points>
<connection>
<GID>7975</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3451.5,48,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3436,48,-3436</points>
<connection>
<GID>7973</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5567</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3451.5,77,-3451.5</points>
<connection>
<GID>7979</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3451.5,71,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3436,71,-3436</points>
<connection>
<GID>7977</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5568</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3451.5,102,-3451.5</points>
<connection>
<GID>7983</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3451.5,96,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3436,96,-3436</points>
<connection>
<GID>7981</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5569</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3451.5,125,-3451.5</points>
<connection>
<GID>7987</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3451.5,119,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3436,119,-3436</points>
<connection>
<GID>7985</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5570</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3451.5,148,-3451.5</points>
<connection>
<GID>7991</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3451.5,142,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3436,142,-3436</points>
<connection>
<GID>7989</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5571</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3451.5,171,-3451.5</points>
<connection>
<GID>7995</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3451.5,165,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3436,165,-3436</points>
<connection>
<GID>7993</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5572</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3451.5,196,-3451.5</points>
<connection>
<GID>7999</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3451.5,190,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3436,190,-3436</points>
<connection>
<GID>7997</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3451.5,219,-3451.5</points>
<connection>
<GID>8003</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3451.5,213,-3436</points>
<intersection>-3451.5 1</intersection>
<intersection>-3436 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3436,213,-3436</points>
<connection>
<GID>8001</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3439,206,-3439</points>
<connection>
<GID>7969</GID>
<name>OUT</name></connection>
<connection>
<GID>7973</GID>
<name>clock</name></connection>
<connection>
<GID>7977</GID>
<name>clock</name></connection>
<connection>
<GID>7981</GID>
<name>clock</name></connection>
<connection>
<GID>7985</GID>
<name>clock</name></connection>
<connection>
<GID>7989</GID>
<name>clock</name></connection>
<connection>
<GID>7993</GID>
<name>clock</name></connection>
<connection>
<GID>7997</GID>
<name>clock</name></connection>
<connection>
<GID>8001</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5575</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3448.5,217,-3448.5</points>
<connection>
<GID>7971</GID>
<name>OUT</name></connection>
<connection>
<GID>7975</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7979</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7983</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7987</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7991</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7995</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7999</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8003</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5576</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3432.5,54,-3432.5</points>
<connection>
<GID>8013</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3432.5,48,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3417,48,-3417</points>
<connection>
<GID>8011</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3432.5,77,-3432.5</points>
<connection>
<GID>8018</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3432.5,71,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3417,71,-3417</points>
<connection>
<GID>8016</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3432.5,102,-3432.5</points>
<connection>
<GID>8023</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3432.5,96,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3417,96,-3417</points>
<connection>
<GID>8021</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3432.5,125,-3432.5</points>
<connection>
<GID>8028</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3432.5,119,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3417,119,-3417</points>
<connection>
<GID>8026</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3432.5,148,-3432.5</points>
<connection>
<GID>8033</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3432.5,142,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3417,142,-3417</points>
<connection>
<GID>8031</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3432.5,171,-3432.5</points>
<connection>
<GID>8036</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3432.5,165,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3417,165,-3417</points>
<connection>
<GID>8035</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3432.5,196,-3432.5</points>
<connection>
<GID>8039</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3432.5,190,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3417,190,-3417</points>
<connection>
<GID>8038</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3432.5,219,-3432.5</points>
<connection>
<GID>8041</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3432.5,213,-3417</points>
<intersection>-3432.5 1</intersection>
<intersection>-3417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3417,213,-3417</points>
<connection>
<GID>8040</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3420,206,-3420</points>
<connection>
<GID>8006</GID>
<name>OUT</name></connection>
<connection>
<GID>8011</GID>
<name>clock</name></connection>
<connection>
<GID>8016</GID>
<name>clock</name></connection>
<connection>
<GID>8021</GID>
<name>clock</name></connection>
<connection>
<GID>8026</GID>
<name>clock</name></connection>
<connection>
<GID>8031</GID>
<name>clock</name></connection>
<connection>
<GID>8035</GID>
<name>clock</name></connection>
<connection>
<GID>8038</GID>
<name>clock</name></connection>
<connection>
<GID>8040</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3429.5,217,-3429.5</points>
<connection>
<GID>8008</GID>
<name>OUT</name></connection>
<connection>
<GID>8013</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8018</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8023</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8028</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8033</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8036</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8039</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8041</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3414,54,-3414</points>
<connection>
<GID>8045</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3414,48,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3398.5,48,-3398.5</points>
<connection>
<GID>8044</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3414,77,-3414</points>
<connection>
<GID>8047</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3414,71,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3398.5,71,-3398.5</points>
<connection>
<GID>8046</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5588</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3414,102,-3414</points>
<connection>
<GID>8049</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3414,96,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3398.5,96,-3398.5</points>
<connection>
<GID>8048</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5589</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3414,125,-3414</points>
<connection>
<GID>8051</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3414,119,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3398.5,119,-3398.5</points>
<connection>
<GID>8050</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5590</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3414,148,-3414</points>
<connection>
<GID>8053</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3414,142,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3398.5,142,-3398.5</points>
<connection>
<GID>8052</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5591</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3414,171,-3414</points>
<connection>
<GID>8055</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3414,165,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3398.5,165,-3398.5</points>
<connection>
<GID>8054</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5592</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3414,196,-3414</points>
<connection>
<GID>8057</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3414,190,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3398.5,190,-3398.5</points>
<connection>
<GID>8056</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3414,219,-3414</points>
<connection>
<GID>8059</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3414,213,-3398.5</points>
<intersection>-3414 1</intersection>
<intersection>-3398.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3398.5,213,-3398.5</points>
<connection>
<GID>8058</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3401.5,206,-3401.5</points>
<connection>
<GID>8042</GID>
<name>OUT</name></connection>
<connection>
<GID>8044</GID>
<name>clock</name></connection>
<connection>
<GID>8046</GID>
<name>clock</name></connection>
<connection>
<GID>8048</GID>
<name>clock</name></connection>
<connection>
<GID>8050</GID>
<name>clock</name></connection>
<connection>
<GID>8052</GID>
<name>clock</name></connection>
<connection>
<GID>8054</GID>
<name>clock</name></connection>
<connection>
<GID>8056</GID>
<name>clock</name></connection>
<connection>
<GID>8058</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3411,217,-3411</points>
<connection>
<GID>8043</GID>
<name>OUT</name></connection>
<connection>
<GID>8045</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8047</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8049</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8051</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8053</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8055</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8057</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8059</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-3480,35.5,-3315</points>
<connection>
<GID>8075</GID>
<name>N_in1</name></connection>
<connection>
<GID>8060</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 12</intersection>
<intersection>-3436 11</intersection>
<intersection>-3417 10</intersection>
<intersection>-3398.5 9</intersection>
<intersection>-3376.5 8</intersection>
<intersection>-3358 7</intersection>
<intersection>-3339 6</intersection>
<intersection>-3320.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-3320.5,41,-3320.5</points>
<connection>
<GID>8264</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-3339,41,-3339</points>
<connection>
<GID>8228</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-3358,41,-3358</points>
<connection>
<GID>8192</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-3376.5,41,-3376.5</points>
<connection>
<GID>8138</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>35.5,-3398.5,41,-3398.5</points>
<connection>
<GID>8044</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>35.5,-3417,41,-3417</points>
<connection>
<GID>8011</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>35.5,-3436,41,-3436</points>
<connection>
<GID>7973</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>35.5,-3454.5,41,-3454.5</points>
<connection>
<GID>8300</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-3479.5,58.5,-3314.5</points>
<connection>
<GID>8076</GID>
<name>N_in1</name></connection>
<connection>
<GID>8061</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 4</intersection>
<intersection>-3445 5</intersection>
<intersection>-3426 6</intersection>
<intersection>-3407.5 7</intersection>
<intersection>-3385.5 8</intersection>
<intersection>-3367 9</intersection>
<intersection>-3348 10</intersection>
<intersection>-3329.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-3463.5,58.5,-3463.5</points>
<intersection>54 12</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54,-3445,58.5,-3445</points>
<intersection>54 13</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54,-3426,58.5,-3426</points>
<intersection>54 14</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54,-3407.5,58.5,-3407.5</points>
<intersection>54 15</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-3385.5,58.5,-3385.5</points>
<intersection>54 18</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>54,-3367,58.5,-3367</points>
<intersection>54 19</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>54,-3348,58.5,-3348</points>
<intersection>54 20</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>54,-3329.5,58.5,-3329.5</points>
<intersection>54 21</intersection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>54,-3464.5,54,-3463.5</points>
<connection>
<GID>8302</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>54,-3446,54,-3445</points>
<connection>
<GID>7975</GID>
<name>OUT_0</name></connection>
<intersection>-3445 5</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>54,-3427,54,-3426</points>
<connection>
<GID>8013</GID>
<name>OUT_0</name></connection>
<intersection>-3426 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>54,-3408.5,54,-3407.5</points>
<connection>
<GID>8045</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>54,-3386.5,54,-3385.5</points>
<connection>
<GID>8144</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>54,-3368,54,-3367</points>
<connection>
<GID>8194</GID>
<name>OUT_0</name></connection>
<intersection>-3367 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>54,-3349,54,-3348</points>
<connection>
<GID>8230</GID>
<name>OUT_0</name></connection>
<intersection>-3348 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>54,-3330.5,54,-3329.5</points>
<connection>
<GID>8266</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-3479.5,61.5,-3315</points>
<connection>
<GID>8077</GID>
<name>N_in1</name></connection>
<connection>
<GID>8062</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 10</intersection>
<intersection>-3436 9</intersection>
<intersection>-3417 8</intersection>
<intersection>-3398.5 7</intersection>
<intersection>-3376.5 6</intersection>
<intersection>-3358 5</intersection>
<intersection>-3339 4</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-3320.5,64,-3320.5</points>
<connection>
<GID>8268</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-3339,64,-3339</points>
<connection>
<GID>8232</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61.5,-3358,64,-3358</points>
<connection>
<GID>8196</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61.5,-3376.5,64,-3376.5</points>
<connection>
<GID>8160</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61.5,-3398.5,64,-3398.5</points>
<connection>
<GID>8046</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61.5,-3417,64,-3417</points>
<connection>
<GID>8016</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61.5,-3436,64,-3436</points>
<connection>
<GID>7977</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61.5,-3454.5,64,-3454.5</points>
<connection>
<GID>8304</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-3479.5,81,-3314.5</points>
<connection>
<GID>8078</GID>
<name>N_in1</name></connection>
<connection>
<GID>8063</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 6</intersection>
<intersection>-3445 7</intersection>
<intersection>-3426 8</intersection>
<intersection>-3407.5 9</intersection>
<intersection>-3385.5 10</intersection>
<intersection>-3367 11</intersection>
<intersection>-3348 12</intersection>
<intersection>-3329.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-3463.5,81,-3463.5</points>
<intersection>77 14</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>77,-3445,81,-3445</points>
<intersection>77 15</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>77,-3426,81,-3426</points>
<intersection>77 16</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-3407.5,81,-3407.5</points>
<intersection>77 17</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>77,-3385.5,81,-3385.5</points>
<intersection>77 20</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>77,-3367,81,-3367</points>
<intersection>77 21</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>77,-3348,81,-3348</points>
<intersection>77 22</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>77,-3329.5,81,-3329.5</points>
<intersection>77 23</intersection>
<intersection>81 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>77,-3464.5,77,-3463.5</points>
<connection>
<GID>8306</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>77,-3446,77,-3445</points>
<connection>
<GID>7979</GID>
<name>OUT_0</name></connection>
<intersection>-3445 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>77,-3427,77,-3426</points>
<connection>
<GID>8018</GID>
<name>OUT_0</name></connection>
<intersection>-3426 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>77,-3408.5,77,-3407.5</points>
<connection>
<GID>8047</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>77,-3386.5,77,-3385.5</points>
<connection>
<GID>8162</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>77,-3368,77,-3367</points>
<connection>
<GID>8198</GID>
<name>OUT_0</name></connection>
<intersection>-3367 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>77,-3349,77,-3348</points>
<connection>
<GID>8234</GID>
<name>OUT_0</name></connection>
<intersection>-3348 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>77,-3330.5,77,-3329.5</points>
<connection>
<GID>8270</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-3479.5,84.5,-3314.5</points>
<connection>
<GID>8079</GID>
<name>N_in1</name></connection>
<connection>
<GID>8064</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 13</intersection>
<intersection>-3436 12</intersection>
<intersection>-3417 11</intersection>
<intersection>-3398.5 10</intersection>
<intersection>-3376.5 9</intersection>
<intersection>-3358 8</intersection>
<intersection>-3339 7</intersection>
<intersection>-3320.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-3320.5,89,-3320.5</points>
<connection>
<GID>8272</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-3339,89,-3339</points>
<connection>
<GID>8236</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>84.5,-3358,89,-3358</points>
<connection>
<GID>8200</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84.5,-3376.5,89,-3376.5</points>
<connection>
<GID>8164</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84.5,-3398.5,89,-3398.5</points>
<connection>
<GID>8048</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84.5,-3417,89,-3417</points>
<connection>
<GID>8021</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>84.5,-3436,89,-3436</points>
<connection>
<GID>7981</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>84.5,-3454.5,89,-3454.5</points>
<connection>
<GID>8308</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3479.5,105.5,-3315</points>
<connection>
<GID>8080</GID>
<name>N_in1</name></connection>
<connection>
<GID>8065</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 6</intersection>
<intersection>-3445 7</intersection>
<intersection>-3426 8</intersection>
<intersection>-3407.5 9</intersection>
<intersection>-3385.5 10</intersection>
<intersection>-3367 11</intersection>
<intersection>-3348 12</intersection>
<intersection>-3329.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>102,-3463.5,105.5,-3463.5</points>
<intersection>102 14</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>102,-3445,105.5,-3445</points>
<intersection>102 15</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>102,-3426,105.5,-3426</points>
<intersection>102 16</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>102,-3407.5,105.5,-3407.5</points>
<intersection>102 17</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>102,-3385.5,105.5,-3385.5</points>
<intersection>102 20</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>102,-3367,105.5,-3367</points>
<intersection>102 21</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>102,-3348,105.5,-3348</points>
<intersection>102 22</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>102,-3329.5,105.5,-3329.5</points>
<intersection>102 23</intersection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>102,-3464.5,102,-3463.5</points>
<connection>
<GID>8310</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>102,-3446,102,-3445</points>
<connection>
<GID>7983</GID>
<name>OUT_0</name></connection>
<intersection>-3445 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>102,-3427,102,-3426</points>
<connection>
<GID>8023</GID>
<name>OUT_0</name></connection>
<intersection>-3426 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>102,-3408.5,102,-3407.5</points>
<connection>
<GID>8049</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>102,-3386.5,102,-3385.5</points>
<connection>
<GID>8166</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>102,-3368,102,-3367</points>
<connection>
<GID>8202</GID>
<name>OUT_0</name></connection>
<intersection>-3367 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>102,-3349,102,-3348</points>
<connection>
<GID>8238</GID>
<name>OUT_0</name></connection>
<intersection>-3348 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>102,-3330.5,102,-3329.5</points>
<connection>
<GID>8274</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3479.5,109.5,-3314.5</points>
<connection>
<GID>8081</GID>
<name>N_in1</name></connection>
<connection>
<GID>8066</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 13</intersection>
<intersection>-3436 12</intersection>
<intersection>-3417 11</intersection>
<intersection>-3398.5 10</intersection>
<intersection>-3376.5 9</intersection>
<intersection>-3358 8</intersection>
<intersection>-3339 7</intersection>
<intersection>-3320.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109.5,-3320.5,112,-3320.5</points>
<connection>
<GID>8276</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>109.5,-3339,112,-3339</points>
<connection>
<GID>8240</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109.5,-3358,112,-3358</points>
<connection>
<GID>8204</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>109.5,-3376.5,112,-3376.5</points>
<connection>
<GID>8168</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>109.5,-3398.5,112,-3398.5</points>
<connection>
<GID>8050</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>109.5,-3417,112,-3417</points>
<connection>
<GID>8026</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109.5,-3436,112,-3436</points>
<connection>
<GID>7985</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>109.5,-3454.5,112,-3454.5</points>
<connection>
<GID>7949</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-3479.5,128,-3314.5</points>
<connection>
<GID>8082</GID>
<name>N_in1</name></connection>
<connection>
<GID>8067</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 6</intersection>
<intersection>-3445 7</intersection>
<intersection>-3426 8</intersection>
<intersection>-3407.5 9</intersection>
<intersection>-3385.5 10</intersection>
<intersection>-3367 11</intersection>
<intersection>-3348 12</intersection>
<intersection>-3329.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>125,-3463.5,128,-3463.5</points>
<intersection>125 14</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125,-3445,128,-3445</points>
<intersection>125 15</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>125,-3426,128,-3426</points>
<intersection>125 16</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>125,-3407.5,128,-3407.5</points>
<intersection>125 17</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125,-3385.5,128,-3385.5</points>
<intersection>125 20</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>125,-3367,128,-3367</points>
<intersection>125 21</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>125,-3348,128,-3348</points>
<intersection>125 22</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>125,-3329.5,128,-3329.5</points>
<intersection>125 23</intersection>
<intersection>128 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>125,-3464.5,125,-3463.5</points>
<connection>
<GID>7951</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>125,-3446,125,-3445</points>
<connection>
<GID>7987</GID>
<name>OUT_0</name></connection>
<intersection>-3445 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>125,-3427,125,-3426</points>
<connection>
<GID>8028</GID>
<name>OUT_0</name></connection>
<intersection>-3426 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>125,-3408.5,125,-3407.5</points>
<connection>
<GID>8051</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>125,-3386.5,125,-3385.5</points>
<connection>
<GID>8170</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>125,-3368,125,-3367</points>
<connection>
<GID>8206</GID>
<name>OUT_0</name></connection>
<intersection>-3367 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>125,-3349,125,-3348</points>
<connection>
<GID>8242</GID>
<name>OUT_0</name></connection>
<intersection>-3348 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>125,-3330.5,125,-3329.5</points>
<connection>
<GID>8278</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-3479.5,132,-3314.5</points>
<connection>
<GID>8083</GID>
<name>N_in1</name></connection>
<connection>
<GID>8068</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 13</intersection>
<intersection>-3436 12</intersection>
<intersection>-3417 11</intersection>
<intersection>-3398.5 10</intersection>
<intersection>-3376.5 9</intersection>
<intersection>-3358 8</intersection>
<intersection>-3339 7</intersection>
<intersection>-3320.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>132,-3320.5,135,-3320.5</points>
<connection>
<GID>8280</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>132,-3339,135,-3339</points>
<connection>
<GID>8244</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>132,-3358,135,-3358</points>
<connection>
<GID>8208</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>132,-3376.5,135,-3376.5</points>
<connection>
<GID>8172</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132,-3398.5,135,-3398.5</points>
<connection>
<GID>8052</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132,-3417,135,-3417</points>
<connection>
<GID>8031</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>132,-3436,135,-3436</points>
<connection>
<GID>7989</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132,-3454.5,135,-3454.5</points>
<connection>
<GID>7953</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>5605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-3479,151,-3314.5</points>
<connection>
<GID>8084</GID>
<name>N_in1</name></connection>
<connection>
<GID>8069</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 6</intersection>
<intersection>-3445 7</intersection>
<intersection>-3426 8</intersection>
<intersection>-3407.5 9</intersection>
<intersection>-3385.5 10</intersection>
<intersection>-3367 11</intersection>
<intersection>-3348 12</intersection>
<intersection>-3329.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>148,-3463.5,151,-3463.5</points>
<intersection>148 14</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>148,-3445,151,-3445</points>
<intersection>148 15</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>148,-3426,151,-3426</points>
<intersection>148 16</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>148,-3407.5,151,-3407.5</points>
<intersection>148 17</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>148,-3385.5,151,-3385.5</points>
<intersection>148 20</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>148,-3367,151,-3367</points>
<intersection>148 21</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>148,-3348,151,-3348</points>
<intersection>148 22</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>148,-3329.5,151,-3329.5</points>
<intersection>148 23</intersection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>148,-3464.5,148,-3463.5</points>
<connection>
<GID>7955</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>148,-3446,148,-3445</points>
<connection>
<GID>7991</GID>
<name>OUT_0</name></connection>
<intersection>-3445 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>148,-3427,148,-3426</points>
<connection>
<GID>8033</GID>
<name>OUT_0</name></connection>
<intersection>-3426 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>148,-3408.5,148,-3407.5</points>
<connection>
<GID>8053</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>148,-3386.5,148,-3385.5</points>
<connection>
<GID>8174</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>148,-3368,148,-3367</points>
<connection>
<GID>8210</GID>
<name>OUT_0</name></connection>
<intersection>-3367 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>148,-3349,148,-3348</points>
<connection>
<GID>8246</GID>
<name>OUT_0</name></connection>
<intersection>-3348 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>148,-3330.5,148,-3329.5</points>
<connection>
<GID>8282</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-3479,156,-3314.5</points>
<connection>
<GID>8085</GID>
<name>N_in1</name></connection>
<connection>
<GID>8070</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 13</intersection>
<intersection>-3436 12</intersection>
<intersection>-3417 11</intersection>
<intersection>-3398.5 10</intersection>
<intersection>-3376.5 9</intersection>
<intersection>-3358 8</intersection>
<intersection>-3339 7</intersection>
<intersection>-3320.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>156,-3320.5,158,-3320.5</points>
<connection>
<GID>8284</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>156,-3339,158,-3339</points>
<connection>
<GID>8248</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>156,-3358,158,-3358</points>
<connection>
<GID>8212</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>156,-3376.5,158,-3376.5</points>
<connection>
<GID>8176</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156,-3398.5,158,-3398.5</points>
<connection>
<GID>8054</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>156,-3417,158,-3417</points>
<connection>
<GID>8035</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>156,-3436,158,-3436</points>
<connection>
<GID>7993</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>156,-3454.5,158,-3454.5</points>
<connection>
<GID>7957</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>5607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-3478.5,174,-3314.5</points>
<connection>
<GID>8086</GID>
<name>N_in1</name></connection>
<connection>
<GID>8072</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 16</intersection>
<intersection>-3445 15</intersection>
<intersection>-3426 14</intersection>
<intersection>-3407.5 13</intersection>
<intersection>-3385.5 12</intersection>
<intersection>-3367 11</intersection>
<intersection>-3348 10</intersection>
<intersection>-3329.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>171,-3329.5,174,-3329.5</points>
<intersection>171 26</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>171,-3348,174,-3348</points>
<intersection>171 25</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>171,-3367,174,-3367</points>
<intersection>171 24</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>171,-3385.5,174,-3385.5</points>
<intersection>171 23</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>171,-3407.5,174,-3407.5</points>
<intersection>171 20</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>171,-3426,174,-3426</points>
<intersection>171 19</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>171,-3445,174,-3445</points>
<intersection>171 18</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>171,-3463.5,174,-3463.5</points>
<intersection>171 17</intersection>
<intersection>174 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>171,-3464.5,171,-3463.5</points>
<connection>
<GID>7959</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>171,-3446,171,-3445</points>
<connection>
<GID>7995</GID>
<name>OUT_0</name></connection>
<intersection>-3445 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>171,-3427,171,-3426</points>
<connection>
<GID>8036</GID>
<name>OUT_0</name></connection>
<intersection>-3426 14</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>171,-3408.5,171,-3407.5</points>
<connection>
<GID>8055</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 13</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>171,-3386.5,171,-3385.5</points>
<connection>
<GID>8178</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 12</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>171,-3368,171,-3367</points>
<connection>
<GID>8214</GID>
<name>OUT_0</name></connection>
<intersection>-3367 11</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>171,-3349,171,-3348</points>
<connection>
<GID>8250</GID>
<name>OUT_0</name></connection>
<intersection>-3348 10</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>171,-3330.5,171,-3329.5</points>
<connection>
<GID>8286</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>5608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-3478.5,178.5,-3314.5</points>
<connection>
<GID>8087</GID>
<name>N_in1</name></connection>
<connection>
<GID>8071</GID>
<name>N_in0</name></connection>
<intersection>-3454.5 13</intersection>
<intersection>-3436 12</intersection>
<intersection>-3417 11</intersection>
<intersection>-3398.5 10</intersection>
<intersection>-3376.5 9</intersection>
<intersection>-3358 8</intersection>
<intersection>-3339 7</intersection>
<intersection>-3320.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>178.5,-3320.5,183,-3320.5</points>
<connection>
<GID>8288</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>178.5,-3339,183,-3339</points>
<connection>
<GID>8252</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178.5,-3358,183,-3358</points>
<connection>
<GID>8216</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>178.5,-3376.5,183,-3376.5</points>
<connection>
<GID>8180</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>178.5,-3398.5,183,-3398.5</points>
<connection>
<GID>8056</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>178.5,-3417,183,-3417</points>
<connection>
<GID>8038</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>178.5,-3436,183,-3436</points>
<connection>
<GID>7997</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>178.5,-3454.5,183,-3454.5</points>
<connection>
<GID>7961</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-3478,199.5,-3315</points>
<connection>
<GID>8088</GID>
<name>N_in1</name></connection>
<connection>
<GID>8073</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 6</intersection>
<intersection>-3445 7</intersection>
<intersection>-3426 8</intersection>
<intersection>-3407.5 9</intersection>
<intersection>-3385.5 10</intersection>
<intersection>-3367 11</intersection>
<intersection>-3348 12</intersection>
<intersection>-3329.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196,-3463.5,199.5,-3463.5</points>
<intersection>196 14</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>196,-3445,199.5,-3445</points>
<intersection>196 15</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>196,-3426,199.5,-3426</points>
<intersection>196 16</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>196,-3407.5,199.5,-3407.5</points>
<intersection>196 17</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>196,-3385.5,199.5,-3385.5</points>
<intersection>196 20</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>196,-3367,199.5,-3367</points>
<intersection>196 21</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>196,-3348,199.5,-3348</points>
<intersection>196 22</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>196,-3329.5,199.5,-3329.5</points>
<intersection>196 23</intersection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>196,-3464.5,196,-3463.5</points>
<connection>
<GID>7963</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>196,-3446,196,-3445</points>
<connection>
<GID>7999</GID>
<name>OUT_0</name></connection>
<intersection>-3445 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>196,-3427,196,-3426</points>
<connection>
<GID>8039</GID>
<name>OUT_0</name></connection>
<intersection>-3426 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>196,-3408.5,196,-3407.5</points>
<connection>
<GID>8057</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>196,-3386.5,196,-3385.5</points>
<connection>
<GID>8182</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>196,-3368,196,-3367</points>
<connection>
<GID>8218</GID>
<name>OUT_0</name></connection>
<intersection>-3367 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>196,-3349,196,-3348</points>
<connection>
<GID>8254</GID>
<name>OUT_0</name></connection>
<intersection>-3348 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>196,-3330.5,196,-3329.5</points>
<connection>
<GID>8290</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-3478,203,-3315</points>
<connection>
<GID>8090</GID>
<name>N_in0</name></connection>
<connection>
<GID>8089</GID>
<name>N_in1</name></connection>
<intersection>-3454.5 11</intersection>
<intersection>-3436 10</intersection>
<intersection>-3417 9</intersection>
<intersection>-3398.5 7</intersection>
<intersection>-3376.5 6</intersection>
<intersection>-3358 5</intersection>
<intersection>-3339 4</intersection>
<intersection>-3320.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-3320.5,206,-3320.5</points>
<connection>
<GID>8292</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>203,-3339,206,-3339</points>
<connection>
<GID>8256</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>203,-3358,206,-3358</points>
<connection>
<GID>8220</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>203,-3376.5,206,-3376.5</points>
<connection>
<GID>8184</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-3398.5,206,-3398.5</points>
<connection>
<GID>8058</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>203,-3417,206,-3417</points>
<connection>
<GID>8040</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>203,-3436,206,-3436</points>
<connection>
<GID>8001</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-3454.5,206,-3454.5</points>
<connection>
<GID>7965</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment></shape></wire>
<wire>
<ID>5611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-3478,224,-3316</points>
<connection>
<GID>8091</GID>
<name>N_in1</name></connection>
<connection>
<GID>8074</GID>
<name>N_in0</name></connection>
<intersection>-3463.5 11</intersection>
<intersection>-3445 10</intersection>
<intersection>-3426 9</intersection>
<intersection>-3407.5 8</intersection>
<intersection>-3385.5 7</intersection>
<intersection>-3367 6</intersection>
<intersection>-3348 5</intersection>
<intersection>-3329.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>219,-3329.5,224,-3329.5</points>
<intersection>219 21</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>219,-3348,224,-3348</points>
<intersection>219 20</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>219,-3367,224,-3367</points>
<intersection>219 19</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>219,-3385.5,224,-3385.5</points>
<intersection>219 18</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>219,-3407.5,224,-3407.5</points>
<intersection>219 15</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>219,-3426,224,-3426</points>
<intersection>219 14</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>219,-3445,224,-3445</points>
<intersection>219 13</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>219,-3463.5,224,-3463.5</points>
<intersection>219 12</intersection>
<intersection>224 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>219,-3464.5,219,-3463.5</points>
<connection>
<GID>7967</GID>
<name>OUT_0</name></connection>
<intersection>-3463.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>219,-3446,219,-3445</points>
<connection>
<GID>8003</GID>
<name>OUT_0</name></connection>
<intersection>-3445 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>219,-3427,219,-3426</points>
<connection>
<GID>8041</GID>
<name>OUT_0</name></connection>
<intersection>-3426 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>219,-3408.5,219,-3407.5</points>
<connection>
<GID>8059</GID>
<name>OUT_0</name></connection>
<intersection>-3407.5 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>219,-3386.5,219,-3385.5</points>
<connection>
<GID>8186</GID>
<name>OUT_0</name></connection>
<intersection>-3385.5 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>219,-3368,219,-3367</points>
<connection>
<GID>8222</GID>
<name>OUT_0</name></connection>
<intersection>-3367 6</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>219,-3349,219,-3348</points>
<connection>
<GID>8258</GID>
<name>OUT_0</name></connection>
<intersection>-3348 5</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>219,-3330.5,219,-3329.5</points>
<connection>
<GID>8294</GID>
<name>OUT_0</name></connection>
<intersection>-3329.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>5612</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-133,-3322.5,13.5,-3322.5</points>
<connection>
<GID>8260</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-133,-3474,-133,-3322.5</points>
<connection>
<GID>8097</GID>
<name>OUT_15</name></connection>
<intersection>-3332 4</intersection>
<intersection>-3322.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-133,-3332,25,-3332</points>
<connection>
<GID>8262</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment></shape></wire>
<wire>
<ID>5613</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-132,-3341,13.5,-3341</points>
<connection>
<GID>8224</GID>
<name>IN_0</name></connection>
<intersection>-132 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-132,-3475,-132,-3341</points>
<intersection>-3475 6</intersection>
<intersection>-3350.5 5</intersection>
<intersection>-3341 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-132,-3350.5,25,-3350.5</points>
<connection>
<GID>8226</GID>
<name>IN_0</name></connection>
<intersection>-132 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3475,-132,-3475</points>
<connection>
<GID>8097</GID>
<name>OUT_14</name></connection>
<intersection>-132 4</intersection></hsegment></shape></wire>
<wire>
<ID>5614</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-131,-3360,13.5,-3360</points>
<connection>
<GID>8188</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-131,-3476,-131,-3360</points>
<intersection>-3476 6</intersection>
<intersection>-3369.5 4</intersection>
<intersection>-3360 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-131,-3369.5,25,-3369.5</points>
<connection>
<GID>8190</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3476,-131,-3476</points>
<connection>
<GID>8097</GID>
<name>OUT_13</name></connection>
<intersection>-131 3</intersection></hsegment></shape></wire>
<wire>
<ID>5615</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-130,-3378.5,13.5,-3378.5</points>
<connection>
<GID>8128</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-130,-3477,-130,-3378.5</points>
<intersection>-3477 5</intersection>
<intersection>-3388 4</intersection>
<intersection>-3378.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-130,-3388,25,-3388</points>
<connection>
<GID>8133</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3477,-130,-3477</points>
<connection>
<GID>8097</GID>
<name>OUT_12</name></connection>
<intersection>-130 3</intersection></hsegment></shape></wire>
<wire>
<ID>5616</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-129,-3400.5,13.5,-3400.5</points>
<connection>
<GID>8042</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-129,-3478,-129,-3400.5</points>
<intersection>-3478 6</intersection>
<intersection>-3410 4</intersection>
<intersection>-3400.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-129,-3410,24.5,-3410</points>
<connection>
<GID>8043</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3478,-129,-3478</points>
<connection>
<GID>8097</GID>
<name>OUT_11</name></connection>
<intersection>-129 3</intersection></hsegment></shape></wire>
<wire>
<ID>5617</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-128,-3419,13.5,-3419</points>
<connection>
<GID>8006</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-3479,-128,-3419</points>
<intersection>-3479 5</intersection>
<intersection>-3428.5 4</intersection>
<intersection>-3419 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-3428.5,24.5,-3428.5</points>
<connection>
<GID>8008</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3479,-128,-3479</points>
<connection>
<GID>8097</GID>
<name>OUT_10</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>5618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127,-3438,13.5,-3438</points>
<connection>
<GID>7969</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-127,-3480,-127,-3438</points>
<intersection>-3480 5</intersection>
<intersection>-3447.5 4</intersection>
<intersection>-3438 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-127,-3447.5,24.5,-3447.5</points>
<connection>
<GID>7971</GID>
<name>IN_0</name></connection>
<intersection>-127 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3480,-127,-3480</points>
<connection>
<GID>8097</GID>
<name>OUT_9</name></connection>
<intersection>-127 3</intersection></hsegment></shape></wire>
<wire>
<ID>5619</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,-3456.5,13.5,-3456.5</points>
<connection>
<GID>8296</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-3481,-126,-3456.5</points>
<intersection>-3481 5</intersection>
<intersection>-3466 4</intersection>
<intersection>-3456.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-3466,24.5,-3466</points>
<connection>
<GID>8298</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3481,-126,-3481</points>
<connection>
<GID>8097</GID>
<name>OUT_8</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>5620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-3480,12.5,-3315</points>
<connection>
<GID>8095</GID>
<name>N_in1</name></connection>
<connection>
<GID>8093</GID>
<name>N_in0</name></connection>
<intersection>-3458.5 10</intersection>
<intersection>-3440 9</intersection>
<intersection>-3421 8</intersection>
<intersection>-3402.5 7</intersection>
<intersection>-3380.5 6</intersection>
<intersection>-3362 5</intersection>
<intersection>-3343 4</intersection>
<intersection>-3324.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-3324.5,13.5,-3324.5</points>
<connection>
<GID>8260</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12.5,-3343,13.5,-3343</points>
<connection>
<GID>8224</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>12.5,-3362,13.5,-3362</points>
<connection>
<GID>8188</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>12.5,-3380.5,13.5,-3380.5</points>
<connection>
<GID>8128</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>12.5,-3402.5,13.5,-3402.5</points>
<connection>
<GID>8042</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>12.5,-3421,13.5,-3421</points>
<connection>
<GID>8006</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-3440,13.5,-3440</points>
<connection>
<GID>7969</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>12.5,-3458.5,13.5,-3458.5</points>
<connection>
<GID>8296</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-3480,22.5,-3315</points>
<connection>
<GID>8094</GID>
<name>N_in1</name></connection>
<connection>
<GID>8092</GID>
<name>N_in0</name></connection>
<intersection>-3468 3</intersection>
<intersection>-3449.5 5</intersection>
<intersection>-3430.5 7</intersection>
<intersection>-3412 9</intersection>
<intersection>-3390 11</intersection>
<intersection>-3371.5 13</intersection>
<intersection>-3352.5 15</intersection>
<intersection>-3334 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-3468,24.5,-3468</points>
<connection>
<GID>8298</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>22.5,-3449.5,24.5,-3449.5</points>
<connection>
<GID>7971</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22.5,-3430.5,24.5,-3430.5</points>
<connection>
<GID>8008</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22.5,-3412,24.5,-3412</points>
<connection>
<GID>8043</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>22.5,-3390,25,-3390</points>
<connection>
<GID>8133</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>22.5,-3371.5,25,-3371.5</points>
<connection>
<GID>8190</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>22.5,-3352.5,25,-3352.5</points>
<connection>
<GID>8226</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>22.5,-3334,25,-3334</points>
<connection>
<GID>8262</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3567.5,54,-3567.5</points>
<connection>
<GID>8193</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3567.5,48,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3552,48,-3552</points>
<connection>
<GID>8181</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5623</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3567.5,77,-3567.5</points>
<connection>
<GID>8219</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3567.5,71,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3552,71,-3552</points>
<connection>
<GID>8217</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5624</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3567.5,102,-3567.5</points>
<connection>
<GID>8227</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3567.5,96,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3552,96,-3552</points>
<connection>
<GID>8223</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3567.5,125,-3567.5</points>
<connection>
<GID>8235</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3567.5,119,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3552,119,-3552</points>
<connection>
<GID>8231</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3567.5,148,-3567.5</points>
<connection>
<GID>8241</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3567.5,142,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3552,142,-3552</points>
<connection>
<GID>8237</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3567.5,171,-3567.5</points>
<connection>
<GID>8245</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3567.5,165,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3552,165,-3552</points>
<connection>
<GID>8243</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5628</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3567.5,196,-3567.5</points>
<connection>
<GID>8249</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3567.5,190,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3552,190,-3552</points>
<connection>
<GID>8247</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3567.5,219,-3567.5</points>
<connection>
<GID>8253</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3567.5,213,-3552</points>
<intersection>-3567.5 1</intersection>
<intersection>-3552 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3552,213,-3552</points>
<connection>
<GID>8251</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5630</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3555,206,-3555</points>
<connection>
<GID>8175</GID>
<name>OUT</name></connection>
<connection>
<GID>8181</GID>
<name>clock</name></connection>
<connection>
<GID>8217</GID>
<name>clock</name></connection>
<connection>
<GID>8223</GID>
<name>clock</name></connection>
<connection>
<GID>8231</GID>
<name>clock</name></connection>
<connection>
<GID>8237</GID>
<name>clock</name></connection>
<connection>
<GID>8243</GID>
<name>clock</name></connection>
<connection>
<GID>8247</GID>
<name>clock</name></connection>
<connection>
<GID>8251</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3564.5,217,-3564.5</points>
<connection>
<GID>8177</GID>
<name>OUT</name></connection>
<connection>
<GID>8193</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8219</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8227</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8235</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8241</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8245</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8249</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8253</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5632</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3549,54,-3549</points>
<connection>
<GID>8261</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3549,48,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3533.5,48,-3533.5</points>
<connection>
<GID>8259</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5633</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3549,77,-3549</points>
<connection>
<GID>8265</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3549,71,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3533.5,71,-3533.5</points>
<connection>
<GID>8263</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5634</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3549,102,-3549</points>
<connection>
<GID>8269</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3549,96,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3533.5,96,-3533.5</points>
<connection>
<GID>8267</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3549,125,-3549</points>
<connection>
<GID>8273</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3549,119,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3533.5,119,-3533.5</points>
<connection>
<GID>8271</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5636</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3549,148,-3549</points>
<connection>
<GID>8277</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3549,142,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3533.5,142,-3533.5</points>
<connection>
<GID>8275</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3549,171,-3549</points>
<connection>
<GID>8281</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3549,165,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3533.5,165,-3533.5</points>
<connection>
<GID>8279</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3549,196,-3549</points>
<connection>
<GID>8285</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3549,190,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3533.5,190,-3533.5</points>
<connection>
<GID>8283</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3549,219,-3549</points>
<connection>
<GID>8289</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3549,213,-3533.5</points>
<intersection>-3549 1</intersection>
<intersection>-3533.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3533.5,213,-3533.5</points>
<connection>
<GID>8287</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5640</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3536.5,206,-3536.5</points>
<connection>
<GID>8255</GID>
<name>OUT</name></connection>
<connection>
<GID>8259</GID>
<name>clock</name></connection>
<connection>
<GID>8263</GID>
<name>clock</name></connection>
<connection>
<GID>8267</GID>
<name>clock</name></connection>
<connection>
<GID>8271</GID>
<name>clock</name></connection>
<connection>
<GID>8275</GID>
<name>clock</name></connection>
<connection>
<GID>8279</GID>
<name>clock</name></connection>
<connection>
<GID>8283</GID>
<name>clock</name></connection>
<connection>
<GID>8287</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5641</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3546,217,-3546</points>
<connection>
<GID>8257</GID>
<name>OUT</name></connection>
<connection>
<GID>8261</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8265</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8269</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8273</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8277</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8281</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8285</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8289</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5642</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3530,54,-3530</points>
<connection>
<GID>8297</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3530,48,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3514.5,48,-3514.5</points>
<connection>
<GID>8295</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5643</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3530,77,-3530</points>
<connection>
<GID>8301</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3530,71,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3514.5,71,-3514.5</points>
<connection>
<GID>8299</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5644</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3530,102,-3530</points>
<connection>
<GID>8305</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3530,96,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3514.5,96,-3514.5</points>
<connection>
<GID>8303</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3530,125,-3530</points>
<connection>
<GID>8309</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3530,119,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3514.5,119,-3514.5</points>
<connection>
<GID>8307</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3530,148,-3530</points>
<connection>
<GID>7950</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3530,142,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3514.5,142,-3514.5</points>
<connection>
<GID>8311</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3530,171,-3530</points>
<connection>
<GID>7954</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3530,165,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3514.5,165,-3514.5</points>
<connection>
<GID>7952</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3530,196,-3530</points>
<connection>
<GID>7958</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3530,190,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3514.5,190,-3514.5</points>
<connection>
<GID>7956</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5649</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3530,219,-3530</points>
<connection>
<GID>7962</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3530,213,-3514.5</points>
<intersection>-3530 1</intersection>
<intersection>-3514.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3514.5,213,-3514.5</points>
<connection>
<GID>7960</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3517.5,206,-3517.5</points>
<connection>
<GID>8311</GID>
<name>clock</name></connection>
<connection>
<GID>8307</GID>
<name>clock</name></connection>
<connection>
<GID>8303</GID>
<name>clock</name></connection>
<connection>
<GID>8299</GID>
<name>clock</name></connection>
<connection>
<GID>8295</GID>
<name>clock</name></connection>
<connection>
<GID>8291</GID>
<name>OUT</name></connection>
<connection>
<GID>7960</GID>
<name>clock</name></connection>
<connection>
<GID>7956</GID>
<name>clock</name></connection>
<connection>
<GID>7952</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3527,217,-3527</points>
<connection>
<GID>8309</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8305</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8301</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8297</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8293</GID>
<name>OUT</name></connection>
<connection>
<GID>7962</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7958</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7954</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7950</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5652</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3511.5,54,-3511.5</points>
<connection>
<GID>7970</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3511.5,48,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3496,48,-3496</points>
<connection>
<GID>7968</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3511.5,77,-3511.5</points>
<connection>
<GID>7974</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3511.5,71,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3496,71,-3496</points>
<connection>
<GID>7972</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5654</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3511.5,102,-3511.5</points>
<connection>
<GID>7978</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3511.5,96,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3496,96,-3496</points>
<connection>
<GID>7976</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5655</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3511.5,125,-3511.5</points>
<connection>
<GID>7982</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3511.5,119,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3496,119,-3496</points>
<connection>
<GID>7980</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5656</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3511.5,148,-3511.5</points>
<connection>
<GID>7986</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3511.5,142,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3496,142,-3496</points>
<connection>
<GID>7984</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5657</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3511.5,171,-3511.5</points>
<connection>
<GID>7990</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3511.5,165,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3496,165,-3496</points>
<connection>
<GID>7988</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3511.5,196,-3511.5</points>
<connection>
<GID>7994</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3511.5,190,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3496,190,-3496</points>
<connection>
<GID>7992</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5659</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3511.5,219,-3511.5</points>
<connection>
<GID>7998</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3511.5,213,-3496</points>
<intersection>-3511.5 1</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3496,213,-3496</points>
<connection>
<GID>7996</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5660</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3499,206,-3499</points>
<connection>
<GID>7964</GID>
<name>OUT</name></connection>
<connection>
<GID>7968</GID>
<name>clock</name></connection>
<connection>
<GID>7972</GID>
<name>clock</name></connection>
<connection>
<GID>7976</GID>
<name>clock</name></connection>
<connection>
<GID>7980</GID>
<name>clock</name></connection>
<connection>
<GID>7984</GID>
<name>clock</name></connection>
<connection>
<GID>7988</GID>
<name>clock</name></connection>
<connection>
<GID>7992</GID>
<name>clock</name></connection>
<connection>
<GID>7996</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5661</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-3508.5,217,-3508.5</points>
<connection>
<GID>7966</GID>
<name>OUT</name></connection>
<connection>
<GID>7970</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7974</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7978</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7982</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7986</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7990</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7994</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>7998</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5662</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3645.5,54,-3645.5</points>
<connection>
<GID>8007</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3645.5,48,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3630,48,-3630</points>
<connection>
<GID>8004</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5663</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3645.5,77,-3645.5</points>
<connection>
<GID>8012</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3645.5,71,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3630,71,-3630</points>
<connection>
<GID>8009</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5664</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3645.5,102,-3645.5</points>
<connection>
<GID>8017</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3645.5,96,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3630,96,-3630</points>
<connection>
<GID>8014</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5665</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3645.5,125,-3645.5</points>
<connection>
<GID>8022</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3645.5,119,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3630,119,-3630</points>
<connection>
<GID>8019</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5666</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3645.5,148,-3645.5</points>
<connection>
<GID>8027</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3645.5,142,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3630,142,-3630</points>
<connection>
<GID>8024</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5667</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3645.5,171,-3645.5</points>
<connection>
<GID>8032</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3645.5,165,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3630,165,-3630</points>
<connection>
<GID>8029</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3645.5,196,-3645.5</points>
<connection>
<GID>8099</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3645.5,190,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3630,190,-3630</points>
<connection>
<GID>8098</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3645.5,219,-3645.5</points>
<connection>
<GID>8101</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3645.5,213,-3630</points>
<intersection>-3645.5 1</intersection>
<intersection>-3630 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3630,213,-3630</points>
<connection>
<GID>8100</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5670</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3633,206,-3633</points>
<connection>
<GID>8000</GID>
<name>OUT</name></connection>
<connection>
<GID>8004</GID>
<name>clock</name></connection>
<connection>
<GID>8009</GID>
<name>clock</name></connection>
<connection>
<GID>8014</GID>
<name>clock</name></connection>
<connection>
<GID>8019</GID>
<name>clock</name></connection>
<connection>
<GID>8024</GID>
<name>clock</name></connection>
<connection>
<GID>8029</GID>
<name>clock</name></connection>
<connection>
<GID>8098</GID>
<name>clock</name></connection>
<connection>
<GID>8100</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5671</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3642.5,217,-3642.5</points>
<connection>
<GID>8002</GID>
<name>OUT</name></connection>
<connection>
<GID>8007</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8012</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8017</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8022</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8027</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8032</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8099</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8101</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5672</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3627,54,-3627</points>
<connection>
<GID>8105</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3627,48,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3611.5,48,-3611.5</points>
<connection>
<GID>8104</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5673</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3627,77,-3627</points>
<connection>
<GID>8107</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3627,71,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3611.5,71,-3611.5</points>
<connection>
<GID>8106</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5674</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3627,102,-3627</points>
<connection>
<GID>8109</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3627,96,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3611.5,96,-3611.5</points>
<connection>
<GID>8108</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5675</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3627,125,-3627</points>
<connection>
<GID>8111</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3627,119,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3611.5,119,-3611.5</points>
<connection>
<GID>8110</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5676</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3627,148,-3627</points>
<connection>
<GID>8113</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3627,142,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3611.5,142,-3611.5</points>
<connection>
<GID>8112</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5677</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3627,171,-3627</points>
<connection>
<GID>8115</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3627,165,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3611.5,165,-3611.5</points>
<connection>
<GID>8114</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5678</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3627,196,-3627</points>
<connection>
<GID>8117</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3627,190,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3611.5,190,-3611.5</points>
<connection>
<GID>8116</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5679</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3627,219,-3627</points>
<connection>
<GID>8119</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3627,213,-3611.5</points>
<intersection>-3627 1</intersection>
<intersection>-3611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3611.5,213,-3611.5</points>
<connection>
<GID>8118</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5680</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3614.5,206,-3614.5</points>
<connection>
<GID>8102</GID>
<name>OUT</name></connection>
<connection>
<GID>8104</GID>
<name>clock</name></connection>
<connection>
<GID>8106</GID>
<name>clock</name></connection>
<connection>
<GID>8108</GID>
<name>clock</name></connection>
<connection>
<GID>8110</GID>
<name>clock</name></connection>
<connection>
<GID>8112</GID>
<name>clock</name></connection>
<connection>
<GID>8114</GID>
<name>clock</name></connection>
<connection>
<GID>8116</GID>
<name>clock</name></connection>
<connection>
<GID>8118</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5681</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3624,217,-3624</points>
<connection>
<GID>8103</GID>
<name>OUT</name></connection>
<connection>
<GID>8105</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8107</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8109</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8111</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8113</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8115</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8117</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8119</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5682</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3608,54,-3608</points>
<connection>
<GID>8015</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3608,48,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3592.5,48,-3592.5</points>
<connection>
<GID>8010</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5683</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3608,77,-3608</points>
<connection>
<GID>8025</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3608,71,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3592.5,71,-3592.5</points>
<connection>
<GID>8020</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5684</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3608,102,-3608</points>
<connection>
<GID>8034</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3608,96,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3592.5,96,-3592.5</points>
<connection>
<GID>8030</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5685</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3608,125,-3608</points>
<connection>
<GID>8121</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3608,119,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3592.5,119,-3592.5</points>
<connection>
<GID>8037</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5686</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3608,148,-3608</points>
<connection>
<GID>8123</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3608,142,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3592.5,142,-3592.5</points>
<connection>
<GID>8122</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5687</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3608,171,-3608</points>
<connection>
<GID>8125</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3608,165,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3592.5,165,-3592.5</points>
<connection>
<GID>8124</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5688</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3608,196,-3608</points>
<connection>
<GID>8127</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3608,190,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3592.5,190,-3592.5</points>
<connection>
<GID>8126</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5689</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3608,219,-3608</points>
<connection>
<GID>8130</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3608,213,-3592.5</points>
<intersection>-3608 1</intersection>
<intersection>-3592.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3592.5,213,-3592.5</points>
<connection>
<GID>8129</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5690</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3595.5,206,-3595.5</points>
<connection>
<GID>8129</GID>
<name>clock</name></connection>
<connection>
<GID>8126</GID>
<name>clock</name></connection>
<connection>
<GID>8124</GID>
<name>clock</name></connection>
<connection>
<GID>8122</GID>
<name>clock</name></connection>
<connection>
<GID>8120</GID>
<name>OUT</name></connection>
<connection>
<GID>8037</GID>
<name>clock</name></connection>
<connection>
<GID>8030</GID>
<name>clock</name></connection>
<connection>
<GID>8020</GID>
<name>clock</name></connection>
<connection>
<GID>8010</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5691</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3605,217,-3605</points>
<connection>
<GID>8005</GID>
<name>OUT</name></connection>
<connection>
<GID>8015</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8025</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8034</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8121</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8123</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8125</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8127</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8130</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5692</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-3589.5,54,-3589.5</points>
<connection>
<GID>8135</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-3589.5,48,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47,-3574,48,-3574</points>
<connection>
<GID>8134</GID>
<name>OUT_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>5693</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-3589.5,77,-3589.5</points>
<connection>
<GID>8137</GID>
<name>IN_0</name></connection>
<intersection>71 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,-3589.5,71,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-3574,71,-3574</points>
<connection>
<GID>8136</GID>
<name>OUT_0</name></connection>
<intersection>71 2</intersection></hsegment></shape></wire>
<wire>
<ID>5694</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-3589.5,102,-3589.5</points>
<connection>
<GID>8140</GID>
<name>IN_0</name></connection>
<intersection>96 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-3589.5,96,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-3574,96,-3574</points>
<connection>
<GID>8139</GID>
<name>OUT_0</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>5695</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>119,-3589.5,125,-3589.5</points>
<connection>
<GID>8142</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,-3589.5,119,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-3574,119,-3574</points>
<connection>
<GID>8141</GID>
<name>OUT_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>5696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-3589.5,148,-3589.5</points>
<connection>
<GID>8145</GID>
<name>IN_0</name></connection>
<intersection>142 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142,-3589.5,142,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-3574,142,-3574</points>
<connection>
<GID>8143</GID>
<name>OUT_0</name></connection>
<intersection>142 2</intersection></hsegment></shape></wire>
<wire>
<ID>5697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-3589.5,171,-3589.5</points>
<connection>
<GID>8147</GID>
<name>IN_0</name></connection>
<intersection>165 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>165,-3589.5,165,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164,-3574,165,-3574</points>
<connection>
<GID>8146</GID>
<name>OUT_0</name></connection>
<intersection>165 2</intersection></hsegment></shape></wire>
<wire>
<ID>5698</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-3589.5,196,-3589.5</points>
<connection>
<GID>8149</GID>
<name>IN_0</name></connection>
<intersection>190 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>190,-3589.5,190,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189,-3574,190,-3574</points>
<connection>
<GID>8148</GID>
<name>OUT_0</name></connection>
<intersection>190 2</intersection></hsegment></shape></wire>
<wire>
<ID>5699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213,-3589.5,219,-3589.5</points>
<connection>
<GID>8151</GID>
<name>IN_0</name></connection>
<intersection>213 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>213,-3589.5,213,-3574</points>
<intersection>-3589.5 1</intersection>
<intersection>-3574 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>212,-3574,213,-3574</points>
<connection>
<GID>8150</GID>
<name>OUT_0</name></connection>
<intersection>213 2</intersection></hsegment></shape></wire>
<wire>
<ID>5700</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-3577,206,-3577</points>
<connection>
<GID>8131</GID>
<name>OUT</name></connection>
<connection>
<GID>8134</GID>
<name>clock</name></connection>
<connection>
<GID>8136</GID>
<name>clock</name></connection>
<connection>
<GID>8139</GID>
<name>clock</name></connection>
<connection>
<GID>8141</GID>
<name>clock</name></connection>
<connection>
<GID>8143</GID>
<name>clock</name></connection>
<connection>
<GID>8146</GID>
<name>clock</name></connection>
<connection>
<GID>8148</GID>
<name>clock</name></connection>
<connection>
<GID>8150</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>5701</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-3586.5,217,-3586.5</points>
<connection>
<GID>8132</GID>
<name>OUT</name></connection>
<connection>
<GID>8135</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8137</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8140</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8142</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8145</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8147</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8149</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>8151</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-3655.5,35.5,-3490.5</points>
<connection>
<GID>8179</GID>
<name>N_in1</name></connection>
<connection>
<GID>8152</GID>
<name>N_in0</name></connection>
<intersection>-3630 12</intersection>
<intersection>-3611.5 11</intersection>
<intersection>-3592.5 10</intersection>
<intersection>-3574 9</intersection>
<intersection>-3552 8</intersection>
<intersection>-3533.5 7</intersection>
<intersection>-3514.5 6</intersection>
<intersection>-3496 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-3496,41,-3496</points>
<connection>
<GID>7968</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-3514.5,41,-3514.5</points>
<connection>
<GID>8295</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-3533.5,41,-3533.5</points>
<connection>
<GID>8259</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-3552,41,-3552</points>
<connection>
<GID>8181</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>35.5,-3574,41,-3574</points>
<connection>
<GID>8134</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>35.5,-3592.5,41,-3592.5</points>
<connection>
<GID>8010</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>35.5,-3611.5,41,-3611.5</points>
<connection>
<GID>8104</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>35.5,-3630,41,-3630</points>
<connection>
<GID>8004</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-3655,58.5,-3490</points>
<connection>
<GID>8183</GID>
<name>N_in1</name></connection>
<connection>
<GID>8153</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 4</intersection>
<intersection>-3620 5</intersection>
<intersection>-3601 6</intersection>
<intersection>-3582.5 7</intersection>
<intersection>-3560.5 8</intersection>
<intersection>-3542 9</intersection>
<intersection>-3523 10</intersection>
<intersection>-3504.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-3638.5,58.5,-3638.5</points>
<intersection>54 12</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54,-3620,58.5,-3620</points>
<intersection>54 14</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54,-3601,58.5,-3601</points>
<intersection>54 13</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54,-3582.5,58.5,-3582.5</points>
<intersection>54 15</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-3560.5,58.5,-3560.5</points>
<intersection>54 18</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>54,-3542,58.5,-3542</points>
<intersection>54 19</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>54,-3523,58.5,-3523</points>
<intersection>54 20</intersection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>54,-3504.5,58.5,-3504.5</points>
<intersection>54 21</intersection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>54,-3640,54,-3638.5</points>
<connection>
<GID>8007</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>54,-3602.5,54,-3601</points>
<connection>
<GID>8015</GID>
<name>OUT_0</name></connection>
<intersection>-3601 6</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>54,-3621.5,54,-3620</points>
<connection>
<GID>8105</GID>
<name>OUT_0</name></connection>
<intersection>-3620 5</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>54,-3584,54,-3582.5</points>
<connection>
<GID>8135</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 7</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>54,-3562,54,-3560.5</points>
<connection>
<GID>8193</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>54,-3543.5,54,-3542</points>
<connection>
<GID>8261</GID>
<name>OUT_0</name></connection>
<intersection>-3542 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>54,-3524.5,54,-3523</points>
<connection>
<GID>8297</GID>
<name>OUT_0</name></connection>
<intersection>-3523 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>54,-3506,54,-3504.5</points>
<connection>
<GID>7970</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>5704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-3655,61.5,-3490.5</points>
<connection>
<GID>8185</GID>
<name>N_in1</name></connection>
<connection>
<GID>8154</GID>
<name>N_in0</name></connection>
<intersection>-3630 10</intersection>
<intersection>-3611.5 9</intersection>
<intersection>-3592.5 8</intersection>
<intersection>-3574 7</intersection>
<intersection>-3552 6</intersection>
<intersection>-3533.5 5</intersection>
<intersection>-3514.5 4</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-3496,64,-3496</points>
<connection>
<GID>7972</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-3514.5,64,-3514.5</points>
<connection>
<GID>8299</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61.5,-3533.5,64,-3533.5</points>
<connection>
<GID>8263</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61.5,-3552,64,-3552</points>
<connection>
<GID>8217</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61.5,-3574,64,-3574</points>
<connection>
<GID>8136</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61.5,-3592.5,64,-3592.5</points>
<connection>
<GID>8020</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61.5,-3611.5,64,-3611.5</points>
<connection>
<GID>8106</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61.5,-3630,64,-3630</points>
<connection>
<GID>8009</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-3655,81,-3490</points>
<connection>
<GID>8187</GID>
<name>N_in1</name></connection>
<connection>
<GID>8155</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 6</intersection>
<intersection>-3620 7</intersection>
<intersection>-3601 8</intersection>
<intersection>-3582.5 9</intersection>
<intersection>-3560.5 10</intersection>
<intersection>-3542 11</intersection>
<intersection>-3523 12</intersection>
<intersection>-3504.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-3638.5,81,-3638.5</points>
<intersection>77 14</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>77,-3620,81,-3620</points>
<intersection>77 16</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>77,-3601,81,-3601</points>
<intersection>77 15</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-3582.5,81,-3582.5</points>
<intersection>77 17</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>77,-3560.5,81,-3560.5</points>
<intersection>77 20</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>77,-3542,81,-3542</points>
<intersection>77 21</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>77,-3523,81,-3523</points>
<intersection>77 22</intersection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>77,-3504.5,81,-3504.5</points>
<intersection>77 23</intersection>
<intersection>81 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>77,-3640,77,-3638.5</points>
<connection>
<GID>8012</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>77,-3602.5,77,-3601</points>
<connection>
<GID>8025</GID>
<name>OUT_0</name></connection>
<intersection>-3601 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>77,-3621.5,77,-3620</points>
<connection>
<GID>8107</GID>
<name>OUT_0</name></connection>
<intersection>-3620 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>77,-3584,77,-3582.5</points>
<connection>
<GID>8137</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>77,-3562,77,-3560.5</points>
<connection>
<GID>8219</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>77,-3543.5,77,-3542</points>
<connection>
<GID>8265</GID>
<name>OUT_0</name></connection>
<intersection>-3542 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>77,-3524.5,77,-3523</points>
<connection>
<GID>8301</GID>
<name>OUT_0</name></connection>
<intersection>-3523 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>77,-3506,77,-3504.5</points>
<connection>
<GID>7974</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5706</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-3655,84.5,-3490</points>
<connection>
<GID>8189</GID>
<name>N_in1</name></connection>
<connection>
<GID>8156</GID>
<name>N_in0</name></connection>
<intersection>-3630 13</intersection>
<intersection>-3611.5 12</intersection>
<intersection>-3592.5 11</intersection>
<intersection>-3574 10</intersection>
<intersection>-3552 9</intersection>
<intersection>-3533.5 8</intersection>
<intersection>-3514.5 7</intersection>
<intersection>-3496 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-3496,89,-3496</points>
<connection>
<GID>7976</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-3514.5,89,-3514.5</points>
<connection>
<GID>8303</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>84.5,-3533.5,89,-3533.5</points>
<connection>
<GID>8267</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84.5,-3552,89,-3552</points>
<connection>
<GID>8223</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84.5,-3574,89,-3574</points>
<connection>
<GID>8139</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84.5,-3592.5,89,-3592.5</points>
<connection>
<GID>8030</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>84.5,-3611.5,89,-3611.5</points>
<connection>
<GID>8108</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>84.5,-3630,89,-3630</points>
<connection>
<GID>8014</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3655,105.5,-3490.5</points>
<connection>
<GID>8191</GID>
<name>N_in1</name></connection>
<connection>
<GID>8157</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 6</intersection>
<intersection>-3620 7</intersection>
<intersection>-3601 8</intersection>
<intersection>-3582.5 9</intersection>
<intersection>-3560.5 10</intersection>
<intersection>-3542 11</intersection>
<intersection>-3523 12</intersection>
<intersection>-3504.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>102,-3638.5,105.5,-3638.5</points>
<intersection>102 14</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>102,-3620,105.5,-3620</points>
<intersection>102 16</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>102,-3601,105.5,-3601</points>
<intersection>102 15</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>102,-3582.5,105.5,-3582.5</points>
<intersection>102 17</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>102,-3560.5,105.5,-3560.5</points>
<intersection>102 20</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>102,-3542,105.5,-3542</points>
<intersection>102 21</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>102,-3523,105.5,-3523</points>
<intersection>102 22</intersection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>102,-3504.5,105.5,-3504.5</points>
<intersection>102 23</intersection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>102,-3640,102,-3638.5</points>
<connection>
<GID>8017</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>102,-3602.5,102,-3601</points>
<connection>
<GID>8034</GID>
<name>OUT_0</name></connection>
<intersection>-3601 8</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>102,-3621.5,102,-3620</points>
<connection>
<GID>8109</GID>
<name>OUT_0</name></connection>
<intersection>-3620 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>102,-3584,102,-3582.5</points>
<connection>
<GID>8140</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>102,-3562,102,-3560.5</points>
<connection>
<GID>8227</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>102,-3543.5,102,-3542</points>
<connection>
<GID>8269</GID>
<name>OUT_0</name></connection>
<intersection>-3542 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>102,-3524.5,102,-3523</points>
<connection>
<GID>8305</GID>
<name>OUT_0</name></connection>
<intersection>-3523 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>102,-3506,102,-3504.5</points>
<connection>
<GID>7978</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3655,109.5,-3490</points>
<connection>
<GID>8195</GID>
<name>N_in1</name></connection>
<connection>
<GID>8158</GID>
<name>N_in0</name></connection>
<intersection>-3630 13</intersection>
<intersection>-3611.5 12</intersection>
<intersection>-3592.5 11</intersection>
<intersection>-3574 10</intersection>
<intersection>-3552 9</intersection>
<intersection>-3533.5 8</intersection>
<intersection>-3514.5 7</intersection>
<intersection>-3496 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109.5,-3496,112,-3496</points>
<connection>
<GID>7980</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>109.5,-3514.5,112,-3514.5</points>
<connection>
<GID>8307</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109.5,-3533.5,112,-3533.5</points>
<connection>
<GID>8271</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>109.5,-3552,112,-3552</points>
<connection>
<GID>8231</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>109.5,-3574,112,-3574</points>
<connection>
<GID>8141</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>109.5,-3592.5,112,-3592.5</points>
<connection>
<GID>8037</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109.5,-3611.5,112,-3611.5</points>
<connection>
<GID>8110</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>109.5,-3630,112,-3630</points>
<connection>
<GID>8019</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-3655,128,-3490</points>
<connection>
<GID>8197</GID>
<name>N_in1</name></connection>
<connection>
<GID>8159</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 6</intersection>
<intersection>-3620 7</intersection>
<intersection>-3601 8</intersection>
<intersection>-3582.5 9</intersection>
<intersection>-3560.5 10</intersection>
<intersection>-3542 11</intersection>
<intersection>-3523 12</intersection>
<intersection>-3504.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>125,-3638.5,128,-3638.5</points>
<intersection>125 14</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125,-3620,128,-3620</points>
<intersection>125 15</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>125,-3601,128,-3601</points>
<intersection>125 16</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>125,-3582.5,128,-3582.5</points>
<intersection>125 17</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125,-3560.5,128,-3560.5</points>
<intersection>125 20</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>125,-3542,128,-3542</points>
<intersection>125 21</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>125,-3523,128,-3523</points>
<intersection>125 22</intersection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>125,-3504.5,128,-3504.5</points>
<intersection>125 23</intersection>
<intersection>128 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>125,-3640,125,-3638.5</points>
<connection>
<GID>8022</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 6</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>125,-3621.5,125,-3620</points>
<connection>
<GID>8111</GID>
<name>OUT_0</name></connection>
<intersection>-3620 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>125,-3602.5,125,-3601</points>
<connection>
<GID>8121</GID>
<name>OUT_0</name></connection>
<intersection>-3601 8</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>125,-3584,125,-3582.5</points>
<connection>
<GID>8142</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 9</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>125,-3562,125,-3560.5</points>
<connection>
<GID>8235</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>125,-3543.5,125,-3542</points>
<connection>
<GID>8273</GID>
<name>OUT_0</name></connection>
<intersection>-3542 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>125,-3524.5,125,-3523</points>
<connection>
<GID>8309</GID>
<name>OUT_0</name></connection>
<intersection>-3523 12</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>125,-3506,125,-3504.5</points>
<connection>
<GID>7982</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>5710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-3655,132,-3490</points>
<connection>
<GID>8199</GID>
<name>N_in1</name></connection>
<connection>
<GID>8161</GID>
<name>N_in0</name></connection>
<intersection>-3630 13</intersection>
<intersection>-3611.5 12</intersection>
<intersection>-3592.5 11</intersection>
<intersection>-3574 10</intersection>
<intersection>-3552 9</intersection>
<intersection>-3533.5 8</intersection>
<intersection>-3514.5 7</intersection>
<intersection>-3496 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>132,-3496,135,-3496</points>
<connection>
<GID>7984</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>132,-3514.5,135,-3514.5</points>
<connection>
<GID>8311</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>132,-3533.5,135,-3533.5</points>
<connection>
<GID>8275</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>132,-3552,135,-3552</points>
<connection>
<GID>8237</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132,-3574,135,-3574</points>
<connection>
<GID>8143</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132,-3592.5,135,-3592.5</points>
<connection>
<GID>8122</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>132,-3611.5,135,-3611.5</points>
<connection>
<GID>8112</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132,-3630,135,-3630</points>
<connection>
<GID>8024</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>5711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-3654.5,151,-3490</points>
<connection>
<GID>8201</GID>
<name>N_in1</name></connection>
<connection>
<GID>8163</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 6</intersection>
<intersection>-3620 7</intersection>
<intersection>-3601 8</intersection>
<intersection>-3582.5 9</intersection>
<intersection>-3560.5 10</intersection>
<intersection>-3542 11</intersection>
<intersection>-3523 12</intersection>
<intersection>-3504.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>148,-3638.5,151,-3638.5</points>
<intersection>148 15</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>148,-3620,151,-3620</points>
<intersection>148 16</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>148,-3601,151,-3601</points>
<intersection>148 17</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>148,-3582.5,151,-3582.5</points>
<intersection>148 18</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>148,-3560.5,151,-3560.5</points>
<intersection>148 21</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>148,-3542,151,-3542</points>
<intersection>148 22</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>148,-3523,151,-3523</points>
<intersection>148 23</intersection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>148,-3504.5,151,-3504.5</points>
<intersection>148 14</intersection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>148,-3506,148,-3504.5</points>
<connection>
<GID>7986</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>148,-3640,148,-3638.5</points>
<connection>
<GID>8027</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>148,-3621.5,148,-3620</points>
<connection>
<GID>8113</GID>
<name>OUT_0</name></connection>
<intersection>-3620 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>148,-3602.5,148,-3601</points>
<connection>
<GID>8123</GID>
<name>OUT_0</name></connection>
<intersection>-3601 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>148,-3584,148,-3582.5</points>
<connection>
<GID>8145</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>148,-3562,148,-3560.5</points>
<connection>
<GID>8241</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>148,-3543.5,148,-3542</points>
<connection>
<GID>8277</GID>
<name>OUT_0</name></connection>
<intersection>-3542 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>148,-3524.5,148,-3523</points>
<connection>
<GID>7950</GID>
<name>OUT_0</name></connection>
<intersection>-3523 12</intersection></vsegment></shape></wire>
<wire>
<ID>5712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-3654.5,156,-3490</points>
<connection>
<GID>8203</GID>
<name>N_in1</name></connection>
<connection>
<GID>8165</GID>
<name>N_in0</name></connection>
<intersection>-3630 13</intersection>
<intersection>-3611.5 12</intersection>
<intersection>-3592.5 11</intersection>
<intersection>-3574 10</intersection>
<intersection>-3552 9</intersection>
<intersection>-3533.5 8</intersection>
<intersection>-3514.5 7</intersection>
<intersection>-3496 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>156,-3496,158,-3496</points>
<connection>
<GID>7988</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>156,-3514.5,158,-3514.5</points>
<connection>
<GID>7952</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>156,-3533.5,158,-3533.5</points>
<connection>
<GID>8279</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>156,-3552,158,-3552</points>
<connection>
<GID>8243</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156,-3574,158,-3574</points>
<connection>
<GID>8146</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>156,-3592.5,158,-3592.5</points>
<connection>
<GID>8124</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>156,-3611.5,158,-3611.5</points>
<connection>
<GID>8114</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>156,-3630,158,-3630</points>
<connection>
<GID>8029</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>5713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-3654,174,-3490</points>
<connection>
<GID>8205</GID>
<name>N_in1</name></connection>
<connection>
<GID>8169</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 16</intersection>
<intersection>-3620 15</intersection>
<intersection>-3601 14</intersection>
<intersection>-3582.5 13</intersection>
<intersection>-3560.5 12</intersection>
<intersection>-3542 11</intersection>
<intersection>-3523 10</intersection>
<intersection>-3504.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>171,-3504.5,174,-3504.5</points>
<intersection>171 17</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>171,-3523,174,-3523</points>
<intersection>171 26</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>171,-3542,174,-3542</points>
<intersection>171 25</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>171,-3560.5,174,-3560.5</points>
<intersection>171 24</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>171,-3582.5,174,-3582.5</points>
<intersection>171 21</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>171,-3601,174,-3601</points>
<intersection>171 20</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>171,-3620,174,-3620</points>
<intersection>171 19</intersection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>171,-3638.5,174,-3638.5</points>
<intersection>171 18</intersection>
<intersection>174 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>171,-3506,171,-3504.5</points>
<connection>
<GID>7990</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 9</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>171,-3640,171,-3638.5</points>
<connection>
<GID>8032</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 16</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>171,-3621.5,171,-3620</points>
<connection>
<GID>8115</GID>
<name>OUT_0</name></connection>
<intersection>-3620 15</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>171,-3602.5,171,-3601</points>
<connection>
<GID>8125</GID>
<name>OUT_0</name></connection>
<intersection>-3601 14</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>171,-3584,171,-3582.5</points>
<connection>
<GID>8147</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 13</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>171,-3562,171,-3560.5</points>
<connection>
<GID>8245</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 12</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>171,-3543.5,171,-3542</points>
<connection>
<GID>8281</GID>
<name>OUT_0</name></connection>
<intersection>-3542 11</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>171,-3524.5,171,-3523</points>
<connection>
<GID>7954</GID>
<name>OUT_0</name></connection>
<intersection>-3523 10</intersection></vsegment></shape></wire>
<wire>
<ID>5714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-3654,178.5,-3490</points>
<connection>
<GID>8207</GID>
<name>N_in1</name></connection>
<connection>
<GID>8167</GID>
<name>N_in0</name></connection>
<intersection>-3630 13</intersection>
<intersection>-3611.5 12</intersection>
<intersection>-3592.5 11</intersection>
<intersection>-3574 10</intersection>
<intersection>-3552 9</intersection>
<intersection>-3533.5 8</intersection>
<intersection>-3514.5 7</intersection>
<intersection>-3496 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>178.5,-3496,183,-3496</points>
<connection>
<GID>7992</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>178.5,-3514.5,183,-3514.5</points>
<connection>
<GID>7956</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178.5,-3533.5,183,-3533.5</points>
<connection>
<GID>8283</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>178.5,-3552,183,-3552</points>
<connection>
<GID>8247</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>178.5,-3574,183,-3574</points>
<connection>
<GID>8148</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>178.5,-3592.5,183,-3592.5</points>
<connection>
<GID>8126</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>178.5,-3611.5,183,-3611.5</points>
<connection>
<GID>8116</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>178.5,-3630,183,-3630</points>
<connection>
<GID>8098</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-3653.5,199.5,-3490.5</points>
<connection>
<GID>8209</GID>
<name>N_in1</name></connection>
<connection>
<GID>8171</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 6</intersection>
<intersection>-3620 7</intersection>
<intersection>-3601 8</intersection>
<intersection>-3582.5 9</intersection>
<intersection>-3560.5 10</intersection>
<intersection>-3542 11</intersection>
<intersection>-3523 12</intersection>
<intersection>-3504.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>196,-3638.5,199.5,-3638.5</points>
<intersection>196 15</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>196,-3620,199.5,-3620</points>
<intersection>196 16</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>196,-3601,199.5,-3601</points>
<intersection>196 17</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>196,-3582.5,199.5,-3582.5</points>
<intersection>196 18</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>196,-3560.5,199.5,-3560.5</points>
<intersection>196 21</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>196,-3542,199.5,-3542</points>
<intersection>196 22</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>196,-3523,199.5,-3523</points>
<intersection>196 23</intersection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>196,-3504.5,199.5,-3504.5</points>
<intersection>196 14</intersection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>196,-3506,196,-3504.5</points>
<connection>
<GID>7994</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>196,-3640,196,-3638.5</points>
<connection>
<GID>8099</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 6</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>196,-3621.5,196,-3620</points>
<connection>
<GID>8117</GID>
<name>OUT_0</name></connection>
<intersection>-3620 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>196,-3602.5,196,-3601</points>
<connection>
<GID>8127</GID>
<name>OUT_0</name></connection>
<intersection>-3601 8</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>196,-3584,196,-3582.5</points>
<connection>
<GID>8149</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>196,-3562,196,-3560.5</points>
<connection>
<GID>8249</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 10</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>196,-3543.5,196,-3542</points>
<connection>
<GID>8285</GID>
<name>OUT_0</name></connection>
<intersection>-3542 11</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>196,-3524.5,196,-3523</points>
<connection>
<GID>7958</GID>
<name>OUT_0</name></connection>
<intersection>-3523 12</intersection></vsegment></shape></wire>
<wire>
<ID>5716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-3653.5,203,-3490.5</points>
<connection>
<GID>8213</GID>
<name>N_in0</name></connection>
<connection>
<GID>8211</GID>
<name>N_in1</name></connection>
<intersection>-3630 11</intersection>
<intersection>-3611.5 10</intersection>
<intersection>-3592.5 9</intersection>
<intersection>-3574 7</intersection>
<intersection>-3552 6</intersection>
<intersection>-3533.5 5</intersection>
<intersection>-3514.5 4</intersection>
<intersection>-3496 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203,-3496,206,-3496</points>
<connection>
<GID>7996</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>203,-3514.5,206,-3514.5</points>
<connection>
<GID>7960</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>203,-3533.5,206,-3533.5</points>
<connection>
<GID>8287</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>203,-3552,206,-3552</points>
<connection>
<GID>8251</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-3574,206,-3574</points>
<connection>
<GID>8150</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>203,-3592.5,206,-3592.5</points>
<connection>
<GID>8129</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>203,-3611.5,206,-3611.5</points>
<connection>
<GID>8118</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-3630,206,-3630</points>
<connection>
<GID>8100</GID>
<name>IN_0</name></connection>
<intersection>203 0</intersection></hsegment></shape></wire>
<wire>
<ID>5717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-3653.5,224,-3491.5</points>
<connection>
<GID>8215</GID>
<name>N_in1</name></connection>
<connection>
<GID>8173</GID>
<name>N_in0</name></connection>
<intersection>-3638.5 11</intersection>
<intersection>-3620 10</intersection>
<intersection>-3601 9</intersection>
<intersection>-3582.5 8</intersection>
<intersection>-3560.5 7</intersection>
<intersection>-3542 6</intersection>
<intersection>-3523 5</intersection>
<intersection>-3504.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>219,-3504.5,224,-3504.5</points>
<intersection>219 12</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>219,-3523,224,-3523</points>
<intersection>219 21</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>219,-3542,224,-3542</points>
<intersection>219 20</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>219,-3560.5,224,-3560.5</points>
<intersection>219 19</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>219,-3582.5,224,-3582.5</points>
<intersection>219 16</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>219,-3601,224,-3601</points>
<intersection>219 15</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>219,-3620,224,-3620</points>
<intersection>219 14</intersection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>219,-3638.5,224,-3638.5</points>
<intersection>219 13</intersection>
<intersection>224 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>219,-3506,219,-3504.5</points>
<connection>
<GID>7998</GID>
<name>OUT_0</name></connection>
<intersection>-3504.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>219,-3640,219,-3638.5</points>
<connection>
<GID>8101</GID>
<name>OUT_0</name></connection>
<intersection>-3638.5 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>219,-3621.5,219,-3620</points>
<connection>
<GID>8119</GID>
<name>OUT_0</name></connection>
<intersection>-3620 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>219,-3602.5,219,-3601</points>
<connection>
<GID>8130</GID>
<name>OUT_0</name></connection>
<intersection>-3601 9</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>219,-3584,219,-3582.5</points>
<connection>
<GID>8151</GID>
<name>OUT_0</name></connection>
<intersection>-3582.5 8</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>219,-3562,219,-3560.5</points>
<connection>
<GID>8253</GID>
<name>OUT_0</name></connection>
<intersection>-3560.5 7</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>219,-3543.5,219,-3542</points>
<connection>
<GID>8289</GID>
<name>OUT_0</name></connection>
<intersection>-3542 6</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>219,-3524.5,219,-3523</points>
<connection>
<GID>7962</GID>
<name>OUT_0</name></connection>
<intersection>-3523 5</intersection></vsegment></shape></wire>
<wire>
<ID>5718</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-126,-3498,13.5,-3498</points>
<connection>
<GID>7964</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-126,-3507.5,-126,-3482</points>
<intersection>-3507.5 4</intersection>
<intersection>-3498 2</intersection>
<intersection>-3482 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-126,-3507.5,25,-3507.5</points>
<connection>
<GID>7966</GID>
<name>IN_0</name></connection>
<intersection>-126 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3482,-126,-3482</points>
<connection>
<GID>8097</GID>
<name>OUT_7</name></connection>
<intersection>-126 3</intersection></hsegment></shape></wire>
<wire>
<ID>5719</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-127,-3516.5,13.5,-3516.5</points>
<connection>
<GID>8291</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-127,-3526,-127,-3483</points>
<intersection>-3526 5</intersection>
<intersection>-3516.5 2</intersection>
<intersection>-3483 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-127,-3526,25,-3526</points>
<connection>
<GID>8293</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3483,-127,-3483</points>
<connection>
<GID>8097</GID>
<name>OUT_6</name></connection>
<intersection>-127 4</intersection></hsegment></shape></wire>
<wire>
<ID>5720</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-128,-3535.5,13.5,-3535.5</points>
<connection>
<GID>8255</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-128,-3545,-128,-3484</points>
<intersection>-3545 4</intersection>
<intersection>-3535.5 2</intersection>
<intersection>-3484 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-128,-3545,25,-3545</points>
<connection>
<GID>8257</GID>
<name>IN_0</name></connection>
<intersection>-128 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-133,-3484,-128,-3484</points>
<connection>
<GID>8097</GID>
<name>OUT_5</name></connection>
<intersection>-128 3</intersection></hsegment></shape></wire>
<wire>
<ID>5721</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-129,-3554,13.5,-3554</points>
<connection>
<GID>8175</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-129,-3563.5,-129,-3485</points>
<intersection>-3563.5 4</intersection>
<intersection>-3554 2</intersection>
<intersection>-3485 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-129,-3563.5,25,-3563.5</points>
<connection>
<GID>8177</GID>
<name>IN_0</name></connection>
<intersection>-129 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3485,-129,-3485</points>
<connection>
<GID>8097</GID>
<name>OUT_4</name></connection>
<intersection>-129 3</intersection></hsegment></shape></wire>
<wire>
<ID>5722</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-130,-3576,13.5,-3576</points>
<connection>
<GID>8131</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-130,-3585.5,-130,-3486</points>
<intersection>-3585.5 4</intersection>
<intersection>-3576 1</intersection>
<intersection>-3486 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-130,-3585.5,24.5,-3585.5</points>
<connection>
<GID>8132</GID>
<name>IN_0</name></connection>
<intersection>-130 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3486,-130,-3486</points>
<connection>
<GID>8097</GID>
<name>OUT_3</name></connection>
<intersection>-130 3</intersection></hsegment></shape></wire>
<wire>
<ID>5723</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-131,-3594.5,13.5,-3594.5</points>
<connection>
<GID>8120</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-131,-3604,-131,-3487</points>
<intersection>-3604 4</intersection>
<intersection>-3594.5 1</intersection>
<intersection>-3487 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-131,-3604,24.5,-3604</points>
<connection>
<GID>8005</GID>
<name>IN_0</name></connection>
<intersection>-131 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3487,-131,-3487</points>
<connection>
<GID>8097</GID>
<name>OUT_2</name></connection>
<intersection>-131 3</intersection></hsegment></shape></wire>
<wire>
<ID>5724</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-132,-3613.5,13.5,-3613.5</points>
<connection>
<GID>8102</GID>
<name>IN_0</name></connection>
<intersection>-132 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-132,-3623,-132,-3488</points>
<intersection>-3623 4</intersection>
<intersection>-3613.5 1</intersection>
<intersection>-3488 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-132,-3623,24.5,-3623</points>
<connection>
<GID>8103</GID>
<name>IN_0</name></connection>
<intersection>-132 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-133,-3488,-132,-3488</points>
<connection>
<GID>8097</GID>
<name>OUT_1</name></connection>
<intersection>-132 3</intersection></hsegment></shape></wire>
<wire>
<ID>5725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-133,-3632,13.5,-3632</points>
<connection>
<GID>8000</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-133,-3641.5,-133,-3489</points>
<connection>
<GID>8097</GID>
<name>OUT_0</name></connection>
<intersection>-3641.5 4</intersection>
<intersection>-3632 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-133,-3641.5,24.5,-3641.5</points>
<connection>
<GID>8002</GID>
<name>IN_0</name></connection>
<intersection>-133 3</intersection></hsegment></shape></wire>
<wire>
<ID>5726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-3655.5,12.5,-3490.5</points>
<connection>
<GID>8233</GID>
<name>N_in1</name></connection>
<connection>
<GID>8225</GID>
<name>N_in0</name></connection>
<intersection>-3634 10</intersection>
<intersection>-3615.5 9</intersection>
<intersection>-3596.5 8</intersection>
<intersection>-3578 7</intersection>
<intersection>-3556 6</intersection>
<intersection>-3537.5 5</intersection>
<intersection>-3518.5 4</intersection>
<intersection>-3500 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-3500,13.5,-3500</points>
<connection>
<GID>7964</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12.5,-3518.5,13.5,-3518.5</points>
<connection>
<GID>8291</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>12.5,-3537.5,13.5,-3537.5</points>
<connection>
<GID>8255</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>12.5,-3556,13.5,-3556</points>
<connection>
<GID>8175</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>12.5,-3578,13.5,-3578</points>
<connection>
<GID>8131</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>12.5,-3596.5,13.5,-3596.5</points>
<connection>
<GID>8120</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-3615.5,13.5,-3615.5</points>
<connection>
<GID>8102</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>12.5,-3634,13.5,-3634</points>
<connection>
<GID>8000</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-3655.5,22.5,-3490.5</points>
<connection>
<GID>8229</GID>
<name>N_in1</name></connection>
<connection>
<GID>8221</GID>
<name>N_in0</name></connection>
<intersection>-3643.5 3</intersection>
<intersection>-3625 5</intersection>
<intersection>-3606 7</intersection>
<intersection>-3587.5 9</intersection>
<intersection>-3565.5 11</intersection>
<intersection>-3547 13</intersection>
<intersection>-3528 15</intersection>
<intersection>-3509.5 17</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-3643.5,24.5,-3643.5</points>
<connection>
<GID>8002</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>22.5,-3625,24.5,-3625</points>
<connection>
<GID>8103</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22.5,-3606,24.5,-3606</points>
<connection>
<GID>8005</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22.5,-3587.5,24.5,-3587.5</points>
<connection>
<GID>8132</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>22.5,-3565.5,25,-3565.5</points>
<connection>
<GID>8177</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>22.5,-3547,25,-3547</points>
<connection>
<GID>8257</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>22.5,-3528,25,-3528</points>
<connection>
<GID>8293</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>22.5,-3509.5,25,-3509.5</points>
<connection>
<GID>7966</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-3488.5,12.5,-3482</points>
<connection>
<GID>8225</GID>
<name>N_in1</name></connection>
<connection>
<GID>8095</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-3488.5,22.5,-3482</points>
<connection>
<GID>8221</GID>
<name>N_in1</name></connection>
<connection>
<GID>8094</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5730</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-3488.5,35.5,-3482</points>
<connection>
<GID>8152</GID>
<name>N_in1</name></connection>
<connection>
<GID>8075</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-3488,58.5,-3481.5</points>
<connection>
<GID>8153</GID>
<name>N_in1</name></connection>
<connection>
<GID>8076</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-3488.5,61.5,-3481.5</points>
<connection>
<GID>8154</GID>
<name>N_in1</name></connection>
<connection>
<GID>8077</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-3488,81,-3481.5</points>
<connection>
<GID>8155</GID>
<name>N_in1</name></connection>
<connection>
<GID>8078</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-3488,84.5,-3481.5</points>
<connection>
<GID>8156</GID>
<name>N_in1</name></connection>
<connection>
<GID>8079</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3488.5,105.5,-3481.5</points>
<connection>
<GID>8157</GID>
<name>N_in1</name></connection>
<connection>
<GID>8080</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3488,109.5,-3481.5</points>
<connection>
<GID>8158</GID>
<name>N_in1</name></connection>
<connection>
<GID>8081</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-3488,128,-3481.5</points>
<connection>
<GID>8159</GID>
<name>N_in1</name></connection>
<connection>
<GID>8082</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-3488,132,-3481.5</points>
<connection>
<GID>8161</GID>
<name>N_in1</name></connection>
<connection>
<GID>8083</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-3488,151,-3481</points>
<connection>
<GID>8163</GID>
<name>N_in1</name></connection>
<connection>
<GID>8084</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-3488,156,-3481</points>
<connection>
<GID>8165</GID>
<name>N_in1</name></connection>
<connection>
<GID>8085</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-3488,174,-3480.5</points>
<connection>
<GID>8169</GID>
<name>N_in1</name></connection>
<connection>
<GID>8086</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-3488,178.5,-3480.5</points>
<connection>
<GID>8167</GID>
<name>N_in1</name></connection>
<connection>
<GID>8087</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-3488.5,199.5,-3480</points>
<connection>
<GID>8171</GID>
<name>N_in1</name></connection>
<connection>
<GID>8088</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-3488.5,203,-3480</points>
<connection>
<GID>8213</GID>
<name>N_in1</name></connection>
<connection>
<GID>8089</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>5745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-3489.5,224,-3480</points>
<connection>
<GID>8173</GID>
<name>N_in1</name></connection>
<connection>
<GID>8091</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,7.07075e-007,122.4,-60.5</PageViewport></page 9></circuit>