<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-38.7038,787.47,348.141,596.26</PageViewport></page 0>
<page 1>
<PageViewport>-285.586,111.285,230.208,-143.662</PageViewport></page 1>
<page 2>
<PageViewport>-195.034,41.0687,320.759,-213.878</PageViewport>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>56,-13</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_TRI_STATE</type>
<position>76,-21</position>
<input>
<ID>ENABLE_0</ID>4 </input>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>68,-21</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_DFF_LOW</type>
<position>21,-13</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_TRI_STATE</type>
<position>41,-21</position>
<input>
<ID>ENABLE_0</ID>6 </input>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>33,-21</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>124,-13</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>11</ID>
<type>BA_TRI_STATE</type>
<position>144,-21</position>
<input>
<ID>ENABLE_0</ID>8 </input>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>136,-21</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_DFF_LOW</type>
<position>89,-13</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_TRI_STATE</type>
<position>109,-21</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>101,-21</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_DFF_LOW</type>
<position>193.5,-13</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>11 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>17</ID>
<type>BA_TRI_STATE</type>
<position>213.5,-21</position>
<input>
<ID>ENABLE_0</ID>12 </input>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>205.5,-21</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_DFF_LOW</type>
<position>158.5,-13</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>BA_TRI_STATE</type>
<position>178.5,-21</position>
<input>
<ID>ENABLE_0</ID>14 </input>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>170.5,-21</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_DFF_LOW</type>
<position>261.5,-13</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>BA_TRI_STATE</type>
<position>281.5,-21</position>
<input>
<ID>ENABLE_0</ID>16 </input>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>273.5,-21</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>226.5,-13</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_TRI_STATE</type>
<position>246.5,-21</position>
<input>
<ID>ENABLE_0</ID>18 </input>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND2</type>
<position>238.5,-21</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>2,-14</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>BA_TRI_STATE</type>
<position>5,-22</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>59</ID>
<type>HA_JUNC_2</type>
<position>14.5,-5</position>
<input>
<ID>N_in0</ID>514 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>61</ID>
<type>HA_JUNC_2</type>
<position>45,0</position>
<input>
<ID>N_in0</ID>515 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>62</ID>
<type>HA_JUNC_2</type>
<position>50,-5</position>
<input>
<ID>N_in0</ID>516 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>63</ID>
<type>HA_JUNC_2</type>
<position>80,0</position>
<input>
<ID>N_in0</ID>517 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>64</ID>
<type>HA_JUNC_2</type>
<position>84,-5</position>
<input>
<ID>N_in0</ID>518 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>65</ID>
<type>HA_JUNC_2</type>
<position>115,0</position>
<input>
<ID>N_in0</ID>519 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>66</ID>
<type>HA_JUNC_2</type>
<position>118,-5</position>
<input>
<ID>N_in0</ID>520 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>67</ID>
<type>HA_JUNC_2</type>
<position>150,0</position>
<input>
<ID>N_in0</ID>521 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>68</ID>
<type>HA_JUNC_2</type>
<position>153,-5</position>
<input>
<ID>N_in0</ID>522 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>69</ID>
<type>HA_JUNC_2</type>
<position>184,0</position>
<input>
<ID>N_in0</ID>523 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>70</ID>
<type>HA_JUNC_2</type>
<position>187,-5</position>
<input>
<ID>N_in0</ID>524 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>71</ID>
<type>HA_JUNC_2</type>
<position>219,0</position>
<input>
<ID>N_in0</ID>525 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>72</ID>
<type>HA_JUNC_2</type>
<position>222,-5</position>
<input>
<ID>N_in0</ID>526 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>73</ID>
<type>HA_JUNC_2</type>
<position>251,0</position>
<input>
<ID>N_in0</ID>527 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>74</ID>
<type>HA_JUNC_2</type>
<position>256,-5</position>
<input>
<ID>N_in0</ID>528 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>75</ID>
<type>HA_JUNC_2</type>
<position>288,0</position>
<input>
<ID>N_in0</ID>529 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>547</ID>
<type>AE_DFF_LOW</type>
<position>57,-32</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>381 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>548</ID>
<type>BA_TRI_STATE</type>
<position>77,-40</position>
<input>
<ID>ENABLE_0</ID>382 </input>
<input>
<ID>IN_0</ID>381 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>549</ID>
<type>AA_AND2</type>
<position>69,-40</position>
<input>
<ID>IN_0</ID>381 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>550</ID>
<type>AE_DFF_LOW</type>
<position>22,-32</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>383 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>551</ID>
<type>BA_TRI_STATE</type>
<position>42,-40</position>
<input>
<ID>ENABLE_0</ID>384 </input>
<input>
<ID>IN_0</ID>383 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>552</ID>
<type>AA_AND2</type>
<position>34,-40</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>384 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>553</ID>
<type>AE_DFF_LOW</type>
<position>125,-32</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>385 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>554</ID>
<type>BA_TRI_STATE</type>
<position>145,-40</position>
<input>
<ID>ENABLE_0</ID>386 </input>
<input>
<ID>IN_0</ID>385 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>555</ID>
<type>AA_AND2</type>
<position>137,-40</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>AE_DFF_LOW</type>
<position>90,-32</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>387 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>557</ID>
<type>BA_TRI_STATE</type>
<position>110,-40</position>
<input>
<ID>ENABLE_0</ID>388 </input>
<input>
<ID>IN_0</ID>387 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND2</type>
<position>102,-40</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>388 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>559</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-32</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>389 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>560</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-40</position>
<input>
<ID>ENABLE_0</ID>390 </input>
<input>
<ID>IN_0</ID>389 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_AND2</type>
<position>206.5,-40</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>390 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>562</ID>
<type>AE_DFF_LOW</type>
<position>159.5,-32</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>391 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>563</ID>
<type>BA_TRI_STATE</type>
<position>179.5,-40</position>
<input>
<ID>ENABLE_0</ID>392 </input>
<input>
<ID>IN_0</ID>391 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>564</ID>
<type>AA_AND2</type>
<position>171.5,-40</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>565</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-32</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>393 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>566</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-40</position>
<input>
<ID>ENABLE_0</ID>394 </input>
<input>
<ID>IN_0</ID>393 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>567</ID>
<type>AA_AND2</type>
<position>274.5,-40</position>
<input>
<ID>IN_0</ID>393 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>568</ID>
<type>AE_DFF_LOW</type>
<position>227.5,-32</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>395 </output>
<input>
<ID>clock</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>569</ID>
<type>BA_TRI_STATE</type>
<position>247.5,-40</position>
<input>
<ID>ENABLE_0</ID>396 </input>
<input>
<ID>IN_0</ID>395 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>570</ID>
<type>AA_AND2</type>
<position>239.5,-40</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>571</ID>
<type>AA_AND2</type>
<position>3,-33</position>
<input>
<ID>IN_0</ID>399 </input>
<output>
<ID>OUT</ID>398 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>BA_TRI_STATE</type>
<position>6,-41</position>
<input>
<ID>ENABLE_0</ID>399 </input>
<output>
<ID>OUT_0</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>573</ID>
<type>AE_DFF_LOW</type>
<position>57.5,-52.5</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>400 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>574</ID>
<type>BA_TRI_STATE</type>
<position>77.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>401 </input>
<input>
<ID>IN_0</ID>400 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>575</ID>
<type>AA_AND2</type>
<position>69.5,-60.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>576</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-52.5</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>402 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>577</ID>
<type>BA_TRI_STATE</type>
<position>42.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>403 </input>
<input>
<ID>IN_0</ID>402 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>578</ID>
<type>AA_AND2</type>
<position>34.5,-60.5</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>403 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>579</ID>
<type>AE_DFF_LOW</type>
<position>125.5,-52.5</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>404 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>580</ID>
<type>BA_TRI_STATE</type>
<position>145.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>405 </input>
<input>
<ID>IN_0</ID>404 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>581</ID>
<type>AA_AND2</type>
<position>137.5,-60.5</position>
<input>
<ID>IN_0</ID>404 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>405 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>583</ID>
<type>BA_TRI_STATE</type>
<position>110.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>407 </input>
<input>
<ID>IN_0</ID>406 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>584</ID>
<type>AA_AND2</type>
<position>102.5,-60.5</position>
<input>
<ID>IN_0</ID>406 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>407 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>585</ID>
<type>AE_DFF_LOW</type>
<position>195,-52.5</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>408 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>586</ID>
<type>BA_TRI_STATE</type>
<position>215,-60.5</position>
<input>
<ID>ENABLE_0</ID>409 </input>
<input>
<ID>IN_0</ID>408 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>587</ID>
<type>AA_AND2</type>
<position>207,-60.5</position>
<input>
<ID>IN_0</ID>408 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>588</ID>
<type>AE_DFF_LOW</type>
<position>160,-52.5</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>410 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>589</ID>
<type>BA_TRI_STATE</type>
<position>180,-60.5</position>
<input>
<ID>ENABLE_0</ID>411 </input>
<input>
<ID>IN_0</ID>410 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>590</ID>
<type>AA_AND2</type>
<position>172,-60.5</position>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>591</ID>
<type>AE_DFF_LOW</type>
<position>263,-52.5</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>412 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>592</ID>
<type>BA_TRI_STATE</type>
<position>283,-60.5</position>
<input>
<ID>ENABLE_0</ID>413 </input>
<input>
<ID>IN_0</ID>412 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>593</ID>
<type>AA_AND2</type>
<position>275,-60.5</position>
<input>
<ID>IN_0</ID>412 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>594</ID>
<type>AE_DFF_LOW</type>
<position>228,-52.5</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>414 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>595</ID>
<type>BA_TRI_STATE</type>
<position>248,-60.5</position>
<input>
<ID>ENABLE_0</ID>415 </input>
<input>
<ID>IN_0</ID>414 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_AND2</type>
<position>240,-60.5</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>597</ID>
<type>AA_AND2</type>
<position>3.5,-53.5</position>
<input>
<ID>IN_0</ID>418 </input>
<output>
<ID>OUT</ID>417 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>BA_TRI_STATE</type>
<position>6.5,-61.5</position>
<input>
<ID>ENABLE_0</ID>418 </input>
<output>
<ID>OUT_0</ID>416 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>599</ID>
<type>AE_DFF_LOW</type>
<position>57,-76</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>419 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>600</ID>
<type>BA_TRI_STATE</type>
<position>77,-84</position>
<input>
<ID>ENABLE_0</ID>420 </input>
<input>
<ID>IN_0</ID>419 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>601</ID>
<type>AA_AND2</type>
<position>69,-84</position>
<input>
<ID>IN_0</ID>419 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>602</ID>
<type>AE_DFF_LOW</type>
<position>22,-76</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>421 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>603</ID>
<type>BA_TRI_STATE</type>
<position>42,-84</position>
<input>
<ID>ENABLE_0</ID>422 </input>
<input>
<ID>IN_0</ID>421 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>604</ID>
<type>AA_AND2</type>
<position>34,-84</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>605</ID>
<type>AE_DFF_LOW</type>
<position>125,-76</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>423 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>606</ID>
<type>BA_TRI_STATE</type>
<position>145,-84</position>
<input>
<ID>ENABLE_0</ID>424 </input>
<input>
<ID>IN_0</ID>423 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_AND2</type>
<position>137,-84</position>
<input>
<ID>IN_0</ID>423 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>608</ID>
<type>AE_DFF_LOW</type>
<position>90,-76</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>425 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>609</ID>
<type>BA_TRI_STATE</type>
<position>110,-84</position>
<input>
<ID>ENABLE_0</ID>426 </input>
<input>
<ID>IN_0</ID>425 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_AND2</type>
<position>102,-84</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>426 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>611</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-76</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>427 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>612</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-84</position>
<input>
<ID>ENABLE_0</ID>428 </input>
<input>
<ID>IN_0</ID>427 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>613</ID>
<type>AA_AND2</type>
<position>206.5,-84</position>
<input>
<ID>IN_0</ID>427 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>614</ID>
<type>AE_DFF_LOW</type>
<position>159.5,-76</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>429 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>615</ID>
<type>BA_TRI_STATE</type>
<position>179.5,-84</position>
<input>
<ID>ENABLE_0</ID>430 </input>
<input>
<ID>IN_0</ID>429 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_AND2</type>
<position>171.5,-84</position>
<input>
<ID>IN_0</ID>429 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>617</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-76</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>431 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>618</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-84</position>
<input>
<ID>ENABLE_0</ID>432 </input>
<input>
<ID>IN_0</ID>431 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>619</ID>
<type>AA_AND2</type>
<position>274.5,-84</position>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>620</ID>
<type>AE_DFF_LOW</type>
<position>227.5,-76</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>433 </output>
<input>
<ID>clock</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>621</ID>
<type>BA_TRI_STATE</type>
<position>247.5,-84</position>
<input>
<ID>ENABLE_0</ID>434 </input>
<input>
<ID>IN_0</ID>433 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>622</ID>
<type>AA_AND2</type>
<position>239.5,-84</position>
<input>
<ID>IN_0</ID>433 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>623</ID>
<type>AA_AND2</type>
<position>3,-77</position>
<input>
<ID>IN_0</ID>437 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>624</ID>
<type>BA_TRI_STATE</type>
<position>6,-85</position>
<input>
<ID>ENABLE_0</ID>437 </input>
<output>
<ID>OUT_0</ID>435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>625</ID>
<type>AE_DFF_LOW</type>
<position>57,-100.5</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>438 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>626</ID>
<type>BA_TRI_STATE</type>
<position>77,-108.5</position>
<input>
<ID>ENABLE_0</ID>439 </input>
<input>
<ID>IN_0</ID>438 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>627</ID>
<type>AA_AND2</type>
<position>69,-108.5</position>
<input>
<ID>IN_0</ID>438 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>628</ID>
<type>AE_DFF_LOW</type>
<position>22,-100.5</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>440 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>629</ID>
<type>BA_TRI_STATE</type>
<position>42,-108.5</position>
<input>
<ID>ENABLE_0</ID>441 </input>
<input>
<ID>IN_0</ID>440 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>630</ID>
<type>AA_AND2</type>
<position>34,-108.5</position>
<input>
<ID>IN_0</ID>440 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>441 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>631</ID>
<type>AE_DFF_LOW</type>
<position>125,-100.5</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>442 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>632</ID>
<type>BA_TRI_STATE</type>
<position>145.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>443 </input>
<input>
<ID>IN_0</ID>442 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>633</ID>
<type>AA_AND2</type>
<position>137,-108.5</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>443 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>634</ID>
<type>AE_DFF_LOW</type>
<position>90,-100.5</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>444 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>635</ID>
<type>BA_TRI_STATE</type>
<position>110,-108.5</position>
<input>
<ID>ENABLE_0</ID>445 </input>
<input>
<ID>IN_0</ID>444 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>636</ID>
<type>AA_AND2</type>
<position>102,-108.5</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>637</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-100.5</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>446 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>638</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>447 </input>
<input>
<ID>IN_0</ID>446 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>639</ID>
<type>AA_AND2</type>
<position>206.5,-108.5</position>
<input>
<ID>IN_0</ID>446 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>447 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>640</ID>
<type>AE_DFF_LOW</type>
<position>159.5,-100.5</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>448 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>641</ID>
<type>BA_TRI_STATE</type>
<position>179.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>449 </input>
<input>
<ID>IN_0</ID>448 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>642</ID>
<type>AA_AND2</type>
<position>171.5,-108.5</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>643</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-100.5</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>450 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>644</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>451 </input>
<input>
<ID>IN_0</ID>450 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>645</ID>
<type>AA_AND2</type>
<position>274.5,-108.5</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_DFF_LOW</type>
<position>227.5,-100.5</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>452 </output>
<input>
<ID>clock</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>647</ID>
<type>BA_TRI_STATE</type>
<position>247.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>453 </input>
<input>
<ID>IN_0</ID>452 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>648</ID>
<type>AA_AND2</type>
<position>239.5,-108.5</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>649</ID>
<type>AA_AND2</type>
<position>3,-101.5</position>
<input>
<ID>IN_0</ID>456 </input>
<output>
<ID>OUT</ID>455 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>650</ID>
<type>BA_TRI_STATE</type>
<position>6,-109.5</position>
<input>
<ID>ENABLE_0</ID>456 </input>
<output>
<ID>OUT_0</ID>454 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>651</ID>
<type>AE_DFF_LOW</type>
<position>57,-125</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>457 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>652</ID>
<type>BA_TRI_STATE</type>
<position>77,-133</position>
<input>
<ID>ENABLE_0</ID>458 </input>
<input>
<ID>IN_0</ID>457 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>653</ID>
<type>AA_AND2</type>
<position>69,-133</position>
<input>
<ID>IN_0</ID>457 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>458 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>654</ID>
<type>AE_DFF_LOW</type>
<position>22,-125</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>459 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>655</ID>
<type>BA_TRI_STATE</type>
<position>42,-133</position>
<input>
<ID>ENABLE_0</ID>460 </input>
<input>
<ID>IN_0</ID>459 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>656</ID>
<type>AA_AND2</type>
<position>34,-133</position>
<input>
<ID>IN_0</ID>459 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>657</ID>
<type>AE_DFF_LOW</type>
<position>125,-125</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>461 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>658</ID>
<type>BA_TRI_STATE</type>
<position>145,-133.5</position>
<input>
<ID>ENABLE_0</ID>462 </input>
<input>
<ID>IN_0</ID>461 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_AND2</type>
<position>137,-133</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>660</ID>
<type>AE_DFF_LOW</type>
<position>90,-125</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>463 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>661</ID>
<type>BA_TRI_STATE</type>
<position>110,-133</position>
<input>
<ID>ENABLE_0</ID>464 </input>
<input>
<ID>IN_0</ID>463 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>662</ID>
<type>AA_AND2</type>
<position>102,-133</position>
<input>
<ID>IN_0</ID>463 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>464 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>663</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-125</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>465 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>664</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-133</position>
<input>
<ID>ENABLE_0</ID>466 </input>
<input>
<ID>IN_0</ID>465 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>665</ID>
<type>AA_AND2</type>
<position>206.5,-133</position>
<input>
<ID>IN_0</ID>465 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>666</ID>
<type>AE_DFF_LOW</type>
<position>159.5,-125</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>467 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>667</ID>
<type>BA_TRI_STATE</type>
<position>179.5,-133</position>
<input>
<ID>ENABLE_0</ID>468 </input>
<input>
<ID>IN_0</ID>467 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>668</ID>
<type>AA_AND2</type>
<position>171.5,-133</position>
<input>
<ID>IN_0</ID>467 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>669</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-125</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>469 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>670</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-133</position>
<input>
<ID>ENABLE_0</ID>470 </input>
<input>
<ID>IN_0</ID>469 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>671</ID>
<type>AA_AND2</type>
<position>274.5,-133</position>
<input>
<ID>IN_0</ID>469 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>470 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>672</ID>
<type>AE_DFF_LOW</type>
<position>227.5,-125</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>471 </output>
<input>
<ID>clock</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>673</ID>
<type>BA_TRI_STATE</type>
<position>247.5,-133</position>
<input>
<ID>ENABLE_0</ID>472 </input>
<input>
<ID>IN_0</ID>471 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>674</ID>
<type>AA_AND2</type>
<position>239.5,-133</position>
<input>
<ID>IN_0</ID>471 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_AND2</type>
<position>3,-126</position>
<input>
<ID>IN_0</ID>475 </input>
<output>
<ID>OUT</ID>474 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>676</ID>
<type>BA_TRI_STATE</type>
<position>6,-134</position>
<input>
<ID>ENABLE_0</ID>475 </input>
<output>
<ID>OUT_0</ID>473 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>677</ID>
<type>AE_DFF_LOW</type>
<position>57.5,-148.5</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>476 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>678</ID>
<type>BA_TRI_STATE</type>
<position>77.5,-156.5</position>
<input>
<ID>ENABLE_0</ID>477 </input>
<input>
<ID>IN_0</ID>476 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>679</ID>
<type>AA_AND2</type>
<position>69.5,-156.5</position>
<input>
<ID>IN_0</ID>476 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>477 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>680</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-148.5</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>478 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>681</ID>
<type>BA_TRI_STATE</type>
<position>42.5,-156.5</position>
<input>
<ID>ENABLE_0</ID>479 </input>
<input>
<ID>IN_0</ID>478 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>682</ID>
<type>AA_AND2</type>
<position>34.5,-156.5</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>683</ID>
<type>AE_DFF_LOW</type>
<position>125.5,-148.5</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>480 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>684</ID>
<type>BA_TRI_STATE</type>
<position>145.5,-156.5</position>
<input>
<ID>ENABLE_0</ID>481 </input>
<input>
<ID>IN_0</ID>480 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>685</ID>
<type>AA_AND2</type>
<position>137.5,-156.5</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>686</ID>
<type>AE_DFF_LOW</type>
<position>90.5,-148.5</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>482 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>687</ID>
<type>BA_TRI_STATE</type>
<position>110.5,-156.5</position>
<input>
<ID>ENABLE_0</ID>483 </input>
<input>
<ID>IN_0</ID>482 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>688</ID>
<type>AA_AND2</type>
<position>102.5,-156.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>689</ID>
<type>AE_DFF_LOW</type>
<position>195,-148.5</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>484 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>690</ID>
<type>BA_TRI_STATE</type>
<position>215,-156.5</position>
<input>
<ID>ENABLE_0</ID>485 </input>
<input>
<ID>IN_0</ID>484 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>691</ID>
<type>AA_AND2</type>
<position>207,-156.5</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_DFF_LOW</type>
<position>160,-148.5</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>486 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>693</ID>
<type>BA_TRI_STATE</type>
<position>180,-156.5</position>
<input>
<ID>ENABLE_0</ID>487 </input>
<input>
<ID>IN_0</ID>486 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>694</ID>
<type>AA_AND2</type>
<position>172,-156.5</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>695</ID>
<type>AE_DFF_LOW</type>
<position>263,-148.5</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>488 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>696</ID>
<type>BA_TRI_STATE</type>
<position>283,-156.5</position>
<input>
<ID>ENABLE_0</ID>489 </input>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>697</ID>
<type>AA_AND2</type>
<position>275,-156.5</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>489 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>698</ID>
<type>AE_DFF_LOW</type>
<position>228,-148.5</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>490 </output>
<input>
<ID>clock</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>699</ID>
<type>BA_TRI_STATE</type>
<position>248,-156.5</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>490 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>700</ID>
<type>AA_AND2</type>
<position>240,-156.5</position>
<input>
<ID>IN_0</ID>490 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>491 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_AND2</type>
<position>3.5,-149.5</position>
<input>
<ID>IN_0</ID>494 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>702</ID>
<type>BA_TRI_STATE</type>
<position>6.5,-157.5</position>
<input>
<ID>ENABLE_0</ID>494 </input>
<output>
<ID>OUT_0</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>703</ID>
<type>AE_DFF_LOW</type>
<position>57,-171</position>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>495 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>704</ID>
<type>BA_TRI_STATE</type>
<position>77,-179</position>
<input>
<ID>ENABLE_0</ID>496 </input>
<input>
<ID>IN_0</ID>495 </input>
<output>
<ID>OUT_0</ID>517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>705</ID>
<type>AA_AND2</type>
<position>69,-179</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>706</ID>
<type>AE_DFF_LOW</type>
<position>22,-171</position>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>497 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>707</ID>
<type>BA_TRI_STATE</type>
<position>42,-179</position>
<input>
<ID>ENABLE_0</ID>498 </input>
<input>
<ID>IN_0</ID>497 </input>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>708</ID>
<type>AA_AND2</type>
<position>34,-179</position>
<input>
<ID>IN_0</ID>497 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>498 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>709</ID>
<type>AE_DFF_LOW</type>
<position>125,-171</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>499 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>710</ID>
<type>BA_TRI_STATE</type>
<position>145,-179.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>499 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>711</ID>
<type>AA_AND2</type>
<position>137,-179</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>500 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>712</ID>
<type>AE_DFF_LOW</type>
<position>90,-171</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>501 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>713</ID>
<type>BA_TRI_STATE</type>
<position>110,-179</position>
<input>
<ID>ENABLE_0</ID>502 </input>
<input>
<ID>IN_0</ID>501 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>714</ID>
<type>AA_AND2</type>
<position>102,-179</position>
<input>
<ID>IN_0</ID>501 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>502 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>715</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-171</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>503 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>716</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-179</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>503 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>717</ID>
<type>AA_AND2</type>
<position>206.5,-179</position>
<input>
<ID>IN_0</ID>503 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>718</ID>
<type>AE_DFF_LOW</type>
<position>159.5,-171</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>505 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>719</ID>
<type>BA_TRI_STATE</type>
<position>179.5,-179</position>
<input>
<ID>ENABLE_0</ID>506 </input>
<input>
<ID>IN_0</ID>505 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>720</ID>
<type>AA_AND2</type>
<position>171.5,-179</position>
<input>
<ID>IN_0</ID>505 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>721</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-171</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>507 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>722</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-179</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>507 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>723</ID>
<type>AA_AND2</type>
<position>274.5,-179</position>
<input>
<ID>IN_0</ID>507 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>724</ID>
<type>AE_DFF_LOW</type>
<position>227.5,-171</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>509 </output>
<input>
<ID>clock</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>725</ID>
<type>BA_TRI_STATE</type>
<position>247.5,-179</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>509 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>726</ID>
<type>AA_AND2</type>
<position>239.5,-179</position>
<input>
<ID>IN_0</ID>509 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>727</ID>
<type>AA_AND2</type>
<position>3,-172</position>
<input>
<ID>IN_0</ID>513 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>728</ID>
<type>BA_TRI_STATE</type>
<position>6,-180</position>
<input>
<ID>ENABLE_0</ID>513 </input>
<output>
<ID>OUT_0</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>729</ID>
<type>HA_JUNC_2</type>
<position>14.5,-198.5</position>
<input>
<ID>N_in1</ID>514 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>730</ID>
<type>HA_JUNC_2</type>
<position>45,-193.5</position>
<input>
<ID>N_in1</ID>515 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>731</ID>
<type>HA_JUNC_2</type>
<position>50,-198.5</position>
<input>
<ID>N_in1</ID>516 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>732</ID>
<type>HA_JUNC_2</type>
<position>80,-194</position>
<input>
<ID>N_in1</ID>517 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>733</ID>
<type>HA_JUNC_2</type>
<position>84,-198.5</position>
<input>
<ID>N_in1</ID>518 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>734</ID>
<type>HA_JUNC_2</type>
<position>115,-193.5</position>
<input>
<ID>N_in1</ID>519 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>735</ID>
<type>HA_JUNC_2</type>
<position>118,-198.5</position>
<input>
<ID>N_in1</ID>520 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>736</ID>
<type>HA_JUNC_2</type>
<position>150,-193.5</position>
<input>
<ID>N_in1</ID>521 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>737</ID>
<type>HA_JUNC_2</type>
<position>153,-198.5</position>
<input>
<ID>N_in1</ID>522 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>738</ID>
<type>HA_JUNC_2</type>
<position>184,-193</position>
<input>
<ID>N_in1</ID>523 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>739</ID>
<type>HA_JUNC_2</type>
<position>187,-198.5</position>
<input>
<ID>N_in1</ID>524 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>740</ID>
<type>HA_JUNC_2</type>
<position>219,-193.5</position>
<input>
<ID>N_in1</ID>525 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>741</ID>
<type>HA_JUNC_2</type>
<position>222,-198.5</position>
<input>
<ID>N_in1</ID>526 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>742</ID>
<type>HA_JUNC_2</type>
<position>251,-193</position>
<input>
<ID>N_in1</ID>527 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>743</ID>
<type>HA_JUNC_2</type>
<position>256,-198.5</position>
<input>
<ID>N_in1</ID>528 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>744</ID>
<type>HA_JUNC_2</type>
<position>288,-193</position>
<input>
<ID>N_in1</ID>529 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>746</ID>
<type>AE_DFF_LOW</type>
<position>90.5,-52.5</position>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>406 </output>
<input>
<ID>clock</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>748</ID>
<type>BE_DECODER_3x8</type>
<position>-87,-90</position>
<output>
<ID>OUT_0</ID>513 </output>
<output>
<ID>OUT_1</ID>494 </output>
<output>
<ID>OUT_2</ID>475 </output>
<output>
<ID>OUT_3</ID>456 </output>
<output>
<ID>OUT_4</ID>437 </output>
<output>
<ID>OUT_5</ID>418 </output>
<output>
<ID>OUT_6</ID>399 </output>
<output>
<ID>OUT_7</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,-40,143,-40</points>
<connection>
<GID>554</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>555</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-43,95,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-39,99,-39</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-30,95,-30</points>
<connection>
<GID>556</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-43,110,-43</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-40,108,-40</points>
<connection>
<GID>558</GID>
<name>OUT</name></connection>
<connection>
<GID>557</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-43,199.5,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-39,203.5,-39</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197.5,-30,199.5,-30</points>
<connection>
<GID>559</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199.5,-43,214.5,-43</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-24,61,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-20,65,-20</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-11,61,-11</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61,-24,76,-24</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-40,212.5,-40</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<connection>
<GID>560</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-21,74,-21</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>5</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-43,164.5,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-39,168.5,-39</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-30,164.5,-30</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-43,179.5,-43</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-24,26,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-20,30,-20</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-11,26,-11</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26,-24,41,-24</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-40,177.5,-40</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<connection>
<GID>563</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-21,39,-21</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-43,267.5,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-39,271.5,-39</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-30,267.5,-30</points>
<connection>
<GID>565</GID>
<name>OUT_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>267.5,-43,282.5,-43</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-24,129,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-20,133,-20</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,-11,129,-11</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>129,-24,144,-24</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-40,280.5,-40</points>
<connection>
<GID>567</GID>
<name>OUT</name></connection>
<connection>
<GID>566</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139,-21,142,-21</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>11</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-43,232.5,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,-39,236.5,-39</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230.5,-30,232.5,-30</points>
<connection>
<GID>568</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>232.5,-43,247.5,-43</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-24,94,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-20,98,-20</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,-11,94,-11</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>94,-24,109,-24</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,-40,245.5,-40</points>
<connection>
<GID>570</GID>
<name>OUT</name></connection>
<connection>
<GID>569</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-21,107,-21</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-41,271.5,-41</points>
<connection>
<GID>567</GID>
<name>IN_1</name></connection>
<connection>
<GID>570</GID>
<name>IN_1</name></connection>
<connection>
<GID>561</GID>
<name>IN_1</name></connection>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<connection>
<GID>555</GID>
<name>IN_1</name></connection>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<connection>
<GID>549</GID>
<name>IN_1</name></connection>
<connection>
<GID>572</GID>
<name>OUT_0</name></connection>
<connection>
<GID>552</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-24,198.5,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198.5,-20,202.5,-20</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>196.5,-11,198.5,-11</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,-24,213.5,-24</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-33,259.5,-33</points>
<connection>
<GID>565</GID>
<name>clock</name></connection>
<connection>
<GID>568</GID>
<name>clock</name></connection>
<connection>
<GID>559</GID>
<name>clock</name></connection>
<connection>
<GID>562</GID>
<name>clock</name></connection>
<connection>
<GID>550</GID>
<name>clock</name></connection>
<connection>
<GID>571</GID>
<name>OUT</name></connection>
<connection>
<GID>547</GID>
<name>clock</name></connection>
<connection>
<GID>556</GID>
<name>clock</name></connection>
<connection>
<GID>553</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>208.5,-21,211.5,-21</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83,-87.5,-83,-32</points>
<intersection>-87.5 4</intersection>
<intersection>-39 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83,-32,0,-32</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83,-39,6,-39</points>
<connection>
<GID>572</GID>
<name>ENABLE_0</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84,-87.5,-83,-87.5</points>
<connection>
<GID>748</GID>
<name>OUT_6</name></connection>
<intersection>-83 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-24,163.5,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-20,167.5,-20</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-11,163.5,-11</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>163.5,-24,178.5,-24</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-63.5,62.5,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-59.5,66.5,-59.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-50.5,62.5,-50.5</points>
<connection>
<GID>573</GID>
<name>OUT_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62.5,-63.5,77.5,-63.5</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,-21,176.5,-21</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-60.5,75.5,-60.5</points>
<connection>
<GID>575</GID>
<name>OUT</name></connection>
<connection>
<GID>574</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-24,266.5,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-20,270.5,-20</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>264.5,-11,266.5,-11</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>266.5,-24,281.5,-24</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-63.5,27.5,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-59.5,31.5,-59.5</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-50.5,27.5,-50.5</points>
<connection>
<GID>576</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27.5,-63.5,42.5,-63.5</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276.5,-21,279.5,-21</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>23</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-60.5,40.5,-60.5</points>
<connection>
<GID>578</GID>
<name>OUT</name></connection>
<connection>
<GID>577</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-24,231.5,-11</points>
<intersection>-24 4</intersection>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231.5,-20,235.5,-20</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229.5,-11,231.5,-11</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>231.5,-24,246.5,-24</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-63.5,130.5,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-59.5,134.5,-59.5</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-50.5,130.5,-50.5</points>
<connection>
<GID>579</GID>
<name>OUT_0</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130.5,-63.5,145.5,-63.5</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241.5,-21,244.5,-21</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<connection>
<GID>26</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140.5,-60.5,143.5,-60.5</points>
<connection>
<GID>581</GID>
<name>OUT</name></connection>
<connection>
<GID>580</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-22,270.5,-22</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-63.5,95.5,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-59.5,99.5,-59.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95.5,-63.5,110.5,-63.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>93.5,-50.5,95.5,-50.5</points>
<connection>
<GID>746</GID>
<name>OUT_0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-14,258.5,-14</points>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<connection>
<GID>13</GID>
<name>clock</name></connection>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<connection>
<GID>7</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105.5,-60.5,108.5,-60.5</points>
<connection>
<GID>584</GID>
<name>OUT</name></connection>
<connection>
<GID>583</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-86.5,-84,-13</points>
<connection>
<GID>748</GID>
<name>OUT_7</name></connection>
<intersection>-20 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84,-13,-1,-13</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-84,-20,5,-20</points>
<connection>
<GID>31</GID>
<name>ENABLE_0</name></connection>
<intersection>-84 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200,-63.5,200,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200,-59.5,204,-59.5</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>200 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-50.5,200,-50.5</points>
<connection>
<GID>585</GID>
<name>OUT_0</name></connection>
<intersection>200 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>200,-63.5,215,-63.5</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>200 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>210,-60.5,213,-60.5</points>
<connection>
<GID>587</GID>
<name>OUT</name></connection>
<connection>
<GID>586</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-63.5,165,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-59.5,169,-59.5</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-50.5,165,-50.5</points>
<connection>
<GID>588</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>165,-63.5,180,-63.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175,-60.5,178,-60.5</points>
<connection>
<GID>590</GID>
<name>OUT</name></connection>
<connection>
<GID>589</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268,-63.5,268,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,-59.5,272,-59.5</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266,-50.5,268,-50.5</points>
<connection>
<GID>591</GID>
<name>OUT_0</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>268,-63.5,283,-63.5</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>268 0</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>278,-60.5,281,-60.5</points>
<connection>
<GID>593</GID>
<name>OUT</name></connection>
<connection>
<GID>592</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-63.5,233,-50.5</points>
<intersection>-63.5 4</intersection>
<intersection>-59.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,-59.5,237,-59.5</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>231,-50.5,233,-50.5</points>
<connection>
<GID>594</GID>
<name>OUT_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>233,-63.5,248,-63.5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-60.5,246,-60.5</points>
<connection>
<GID>596</GID>
<name>OUT</name></connection>
<connection>
<GID>595</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-61.5,272,-61.5</points>
<connection>
<GID>593</GID>
<name>IN_1</name></connection>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<connection>
<GID>587</GID>
<name>IN_1</name></connection>
<connection>
<GID>590</GID>
<name>IN_1</name></connection>
<connection>
<GID>581</GID>
<name>IN_1</name></connection>
<connection>
<GID>584</GID>
<name>IN_1</name></connection>
<connection>
<GID>575</GID>
<name>IN_1</name></connection>
<connection>
<GID>578</GID>
<name>IN_1</name></connection>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-53.5,260,-53.5</points>
<connection>
<GID>591</GID>
<name>clock</name></connection>
<connection>
<GID>594</GID>
<name>clock</name></connection>
<connection>
<GID>585</GID>
<name>clock</name></connection>
<connection>
<GID>588</GID>
<name>clock</name></connection>
<connection>
<GID>579</GID>
<name>clock</name></connection>
<connection>
<GID>746</GID>
<name>clock</name></connection>
<connection>
<GID>573</GID>
<name>clock</name></connection>
<connection>
<GID>576</GID>
<name>clock</name></connection>
<connection>
<GID>597</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82,-88.5,-82,-52.5</points>
<intersection>-88.5 4</intersection>
<intersection>-59.5 2</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82,-52.5,0.5,-52.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-59.5,6.5,-59.5</points>
<connection>
<GID>598</GID>
<name>ENABLE_0</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84,-88.5,-82,-88.5</points>
<connection>
<GID>748</GID>
<name>OUT_5</name></connection>
<intersection>-82 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-87,62,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-83,66,-83</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-74,62,-74</points>
<connection>
<GID>599</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62,-87,77,-87</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-84,75,-84</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<connection>
<GID>600</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-87,27,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-83,31,-83</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-74,27,-74</points>
<connection>
<GID>602</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-87,42,-87</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-84,40,-84</points>
<connection>
<GID>604</GID>
<name>OUT</name></connection>
<connection>
<GID>603</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-87,130,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-83,134,-83</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-74,130,-74</points>
<connection>
<GID>605</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-87,145,-87</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,-84,143,-84</points>
<connection>
<GID>607</GID>
<name>OUT</name></connection>
<connection>
<GID>606</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-87,95,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-83,99,-83</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-74,95,-74</points>
<connection>
<GID>608</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-87,110,-87</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-84,108,-84</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<connection>
<GID>609</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-87,199.5,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-83,203.5,-83</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197.5,-74,199.5,-74</points>
<connection>
<GID>611</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199.5,-87,214.5,-87</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-84,212.5,-84</points>
<connection>
<GID>613</GID>
<name>OUT</name></connection>
<connection>
<GID>612</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-87,164.5,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-83,168.5,-83</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-74,164.5,-74</points>
<connection>
<GID>614</GID>
<name>OUT_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-87,179.5,-87</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-84,177.5,-84</points>
<connection>
<GID>616</GID>
<name>OUT</name></connection>
<connection>
<GID>615</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-87,267.5,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-83,271.5,-83</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-74,267.5,-74</points>
<connection>
<GID>617</GID>
<name>OUT_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>267.5,-87,282.5,-87</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-84,280.5,-84</points>
<connection>
<GID>619</GID>
<name>OUT</name></connection>
<connection>
<GID>618</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-87,232.5,-74</points>
<intersection>-87 4</intersection>
<intersection>-83 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,-83,236.5,-83</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230.5,-74,232.5,-74</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>232.5,-87,247.5,-87</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,-84,245.5,-84</points>
<connection>
<GID>622</GID>
<name>OUT</name></connection>
<connection>
<GID>621</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-85,271.5,-85</points>
<connection>
<GID>619</GID>
<name>IN_1</name></connection>
<connection>
<GID>622</GID>
<name>IN_1</name></connection>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<connection>
<GID>616</GID>
<name>IN_1</name></connection>
<connection>
<GID>607</GID>
<name>IN_1</name></connection>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<connection>
<GID>604</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-77,259.5,-77</points>
<connection>
<GID>617</GID>
<name>clock</name></connection>
<connection>
<GID>620</GID>
<name>clock</name></connection>
<connection>
<GID>611</GID>
<name>clock</name></connection>
<connection>
<GID>614</GID>
<name>clock</name></connection>
<connection>
<GID>605</GID>
<name>clock</name></connection>
<connection>
<GID>608</GID>
<name>clock</name></connection>
<connection>
<GID>602</GID>
<name>clock</name></connection>
<connection>
<GID>623</GID>
<name>OUT</name></connection>
<connection>
<GID>599</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,-89.5,-81,-76</points>
<intersection>-89.5 4</intersection>
<intersection>-83 2</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81,-76,0,-76</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-81,-83,6,-83</points>
<connection>
<GID>624</GID>
<name>ENABLE_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84,-89.5,-81,-89.5</points>
<connection>
<GID>748</GID>
<name>OUT_4</name></connection>
<intersection>-81 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-111.5,62,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-107.5,66,-107.5</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-98.5,62,-98.5</points>
<connection>
<GID>625</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62,-111.5,77,-111.5</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-108.5,75,-108.5</points>
<connection>
<GID>627</GID>
<name>OUT</name></connection>
<connection>
<GID>626</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-111.5,27,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-107.5,31,-107.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-98.5,27,-98.5</points>
<connection>
<GID>628</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-111.5,42,-111.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-108.5,40,-108.5</points>
<connection>
<GID>630</GID>
<name>OUT</name></connection>
<connection>
<GID>629</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-112,130,-98.5</points>
<intersection>-112 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-107.5,134,-107.5</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-98.5,130,-98.5</points>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-112,145.5,-112</points>
<intersection>130 0</intersection>
<intersection>145.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>145.5,-112,145.5,-111.5</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>-112 4</intersection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,-108.5,143.5,-108.5</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<connection>
<GID>632</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-111.5,95,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-107.5,99,-107.5</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-98.5,95,-98.5</points>
<connection>
<GID>634</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-111.5,110,-111.5</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-108.5,108,-108.5</points>
<connection>
<GID>636</GID>
<name>OUT</name></connection>
<connection>
<GID>635</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-111.5,199.5,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-107.5,203.5,-107.5</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197.5,-98.5,199.5,-98.5</points>
<connection>
<GID>637</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199.5,-111.5,214.5,-111.5</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-108.5,212.5,-108.5</points>
<connection>
<GID>639</GID>
<name>OUT</name></connection>
<connection>
<GID>638</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-111.5,164.5,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-107.5,168.5,-107.5</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-98.5,164.5,-98.5</points>
<connection>
<GID>640</GID>
<name>OUT_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-111.5,179.5,-111.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-108.5,177.5,-108.5</points>
<connection>
<GID>642</GID>
<name>OUT</name></connection>
<connection>
<GID>641</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-111.5,267.5,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-107.5,271.5,-107.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-98.5,267.5,-98.5</points>
<connection>
<GID>643</GID>
<name>OUT_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>267.5,-111.5,282.5,-111.5</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-108.5,280.5,-108.5</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<connection>
<GID>644</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-111.5,232.5,-98.5</points>
<intersection>-111.5 4</intersection>
<intersection>-107.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,-107.5,236.5,-107.5</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230.5,-98.5,232.5,-98.5</points>
<connection>
<GID>646</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>232.5,-111.5,247.5,-111.5</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,-108.5,245.5,-108.5</points>
<connection>
<GID>648</GID>
<name>OUT</name></connection>
<connection>
<GID>647</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-109.5,271.5,-109.5</points>
<connection>
<GID>645</GID>
<name>IN_1</name></connection>
<connection>
<GID>648</GID>
<name>IN_1</name></connection>
<connection>
<GID>639</GID>
<name>IN_1</name></connection>
<connection>
<GID>642</GID>
<name>IN_1</name></connection>
<connection>
<GID>633</GID>
<name>IN_1</name></connection>
<connection>
<GID>636</GID>
<name>IN_1</name></connection>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection>
<connection>
<GID>630</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-101.5,259.5,-101.5</points>
<connection>
<GID>643</GID>
<name>clock</name></connection>
<connection>
<GID>646</GID>
<name>clock</name></connection>
<connection>
<GID>637</GID>
<name>clock</name></connection>
<connection>
<GID>640</GID>
<name>clock</name></connection>
<connection>
<GID>631</GID>
<name>clock</name></connection>
<connection>
<GID>634</GID>
<name>clock</name></connection>
<connection>
<GID>625</GID>
<name>clock</name></connection>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<connection>
<GID>628</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,-107.5,-81,-90.5</points>
<intersection>-107.5 2</intersection>
<intersection>-100.5 1</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81,-100.5,0,-100.5</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-81,-107.5,6,-107.5</points>
<connection>
<GID>650</GID>
<name>ENABLE_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-84,-90.5,-81,-90.5</points>
<connection>
<GID>748</GID>
<name>OUT_3</name></connection>
<intersection>-81 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-136,62,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-132,66,-132</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-123,62,-123</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62,-136,77,-136</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-133,75,-133</points>
<connection>
<GID>653</GID>
<name>OUT</name></connection>
<connection>
<GID>652</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-136,27,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-132,31,-132</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-123,27,-123</points>
<connection>
<GID>654</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-136,42,-136</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-133,40,-133</points>
<connection>
<GID>656</GID>
<name>OUT</name></connection>
<connection>
<GID>655</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-136,130,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-132,134,-132</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-123,130,-123</points>
<connection>
<GID>657</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-136,145,-136</points>
<intersection>130 0</intersection>
<intersection>145 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>145,-136.5,145,-136</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-136 4</intersection></vsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,-133.5,143,-133.5</points>
<connection>
<GID>658</GID>
<name>ENABLE_0</name></connection>
<intersection>140 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>140,-133.5,140,-133</points>
<connection>
<GID>659</GID>
<name>OUT</name></connection>
<intersection>-133.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-136,95,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-132,99,-132</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-123,95,-123</points>
<connection>
<GID>660</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-136,110,-136</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-133,108,-133</points>
<connection>
<GID>662</GID>
<name>OUT</name></connection>
<connection>
<GID>661</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-136,199.5,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-132,203.5,-132</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197.5,-123,199.5,-123</points>
<connection>
<GID>663</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199.5,-136,214.5,-136</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-133,212.5,-133</points>
<connection>
<GID>665</GID>
<name>OUT</name></connection>
<connection>
<GID>664</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-136,164.5,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-132,168.5,-132</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-123,164.5,-123</points>
<connection>
<GID>666</GID>
<name>OUT_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-136,179.5,-136</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-133,177.5,-133</points>
<connection>
<GID>668</GID>
<name>OUT</name></connection>
<connection>
<GID>667</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-136,267.5,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-132,271.5,-132</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-123,267.5,-123</points>
<connection>
<GID>669</GID>
<name>OUT_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>267.5,-136,282.5,-136</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-133,280.5,-133</points>
<connection>
<GID>671</GID>
<name>OUT</name></connection>
<connection>
<GID>670</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-136,232.5,-123</points>
<intersection>-136 4</intersection>
<intersection>-132 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,-132,236.5,-132</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230.5,-123,232.5,-123</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>232.5,-136,247.5,-136</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,-133,245.5,-133</points>
<connection>
<GID>674</GID>
<name>OUT</name></connection>
<connection>
<GID>673</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-134,271.5,-134</points>
<connection>
<GID>671</GID>
<name>IN_1</name></connection>
<connection>
<GID>674</GID>
<name>IN_1</name></connection>
<connection>
<GID>665</GID>
<name>IN_1</name></connection>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<connection>
<GID>659</GID>
<name>IN_1</name></connection>
<connection>
<GID>662</GID>
<name>IN_1</name></connection>
<connection>
<GID>653</GID>
<name>IN_1</name></connection>
<connection>
<GID>676</GID>
<name>OUT_0</name></connection>
<connection>
<GID>656</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-126,259.5,-126</points>
<connection>
<GID>669</GID>
<name>clock</name></connection>
<connection>
<GID>672</GID>
<name>clock</name></connection>
<connection>
<GID>663</GID>
<name>clock</name></connection>
<connection>
<GID>666</GID>
<name>clock</name></connection>
<connection>
<GID>657</GID>
<name>clock</name></connection>
<connection>
<GID>660</GID>
<name>clock</name></connection>
<connection>
<GID>651</GID>
<name>clock</name></connection>
<connection>
<GID>675</GID>
<name>OUT</name></connection>
<connection>
<GID>654</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82,-132,-82,-91.5</points>
<intersection>-132 2</intersection>
<intersection>-125 1</intersection>
<intersection>-91.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82,-125,0,-125</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-132,6,-132</points>
<connection>
<GID>676</GID>
<name>ENABLE_0</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-84,-91.5,-82,-91.5</points>
<connection>
<GID>748</GID>
<name>OUT_2</name></connection>
<intersection>-82 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-159.5,62.5,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-155.5,66.5,-155.5</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-146.5,62.5,-146.5</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62.5,-159.5,77.5,-159.5</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-156.5,75.5,-156.5</points>
<connection>
<GID>679</GID>
<name>OUT</name></connection>
<connection>
<GID>678</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-159.5,27.5,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-155.5,31.5,-155.5</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-146.5,27.5,-146.5</points>
<connection>
<GID>680</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27.5,-159.5,42.5,-159.5</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-156.5,40.5,-156.5</points>
<connection>
<GID>682</GID>
<name>OUT</name></connection>
<connection>
<GID>681</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-159.5,130.5,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-155.5,134.5,-155.5</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128.5,-146.5,130.5,-146.5</points>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130.5,-159.5,145.5,-159.5</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140.5,-156.5,143.5,-156.5</points>
<connection>
<GID>685</GID>
<name>OUT</name></connection>
<connection>
<GID>684</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-159.5,95.5,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-155.5,99.5,-155.5</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-146.5,95.5,-146.5</points>
<connection>
<GID>686</GID>
<name>OUT_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95.5,-159.5,110.5,-159.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105.5,-156.5,108.5,-156.5</points>
<connection>
<GID>688</GID>
<name>OUT</name></connection>
<connection>
<GID>687</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200,-159.5,200,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200,-155.5,204,-155.5</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>200 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-146.5,200,-146.5</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>200 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>200,-159.5,215,-159.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>200 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>210,-156.5,213,-156.5</points>
<connection>
<GID>691</GID>
<name>OUT</name></connection>
<connection>
<GID>690</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-159.5,165,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-155.5,169,-155.5</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-146.5,165,-146.5</points>
<connection>
<GID>692</GID>
<name>OUT_0</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>165,-159.5,180,-159.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175,-156.5,178,-156.5</points>
<connection>
<GID>694</GID>
<name>OUT</name></connection>
<connection>
<GID>693</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268,-159.5,268,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,-155.5,272,-155.5</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266,-146.5,268,-146.5</points>
<connection>
<GID>695</GID>
<name>OUT_0</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>268,-159.5,283,-159.5</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<intersection>268 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>278,-156.5,281,-156.5</points>
<connection>
<GID>697</GID>
<name>OUT</name></connection>
<connection>
<GID>696</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-159.5,233,-146.5</points>
<intersection>-159.5 4</intersection>
<intersection>-155.5 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,-155.5,237,-155.5</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>231,-146.5,233,-146.5</points>
<connection>
<GID>698</GID>
<name>OUT_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>233,-159.5,248,-159.5</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-156.5,246,-156.5</points>
<connection>
<GID>700</GID>
<name>OUT</name></connection>
<connection>
<GID>699</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-157.5,272,-157.5</points>
<connection>
<GID>697</GID>
<name>IN_1</name></connection>
<connection>
<GID>700</GID>
<name>IN_1</name></connection>
<connection>
<GID>691</GID>
<name>IN_1</name></connection>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<connection>
<GID>685</GID>
<name>IN_1</name></connection>
<connection>
<GID>688</GID>
<name>IN_1</name></connection>
<connection>
<GID>679</GID>
<name>IN_1</name></connection>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<connection>
<GID>682</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-149.5,260,-149.5</points>
<connection>
<GID>695</GID>
<name>clock</name></connection>
<connection>
<GID>698</GID>
<name>clock</name></connection>
<connection>
<GID>689</GID>
<name>clock</name></connection>
<connection>
<GID>692</GID>
<name>clock</name></connection>
<connection>
<GID>683</GID>
<name>clock</name></connection>
<connection>
<GID>686</GID>
<name>clock</name></connection>
<connection>
<GID>677</GID>
<name>clock</name></connection>
<connection>
<GID>701</GID>
<name>OUT</name></connection>
<connection>
<GID>680</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83,-155.5,-83,-92.5</points>
<intersection>-155.5 2</intersection>
<intersection>-148.5 1</intersection>
<intersection>-92.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83,-148.5,0.5,-148.5</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83,-155.5,6.5,-155.5</points>
<connection>
<GID>702</GID>
<name>ENABLE_0</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84,-92.5,-83,-92.5</points>
<connection>
<GID>748</GID>
<name>OUT_1</name></connection>
<intersection>-83 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-182,62,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-178,66,-178</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-169,62,-169</points>
<connection>
<GID>703</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62,-182,77,-182</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-179,75,-179</points>
<connection>
<GID>705</GID>
<name>OUT</name></connection>
<connection>
<GID>704</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-182,27,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-178,31,-178</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-169,27,-169</points>
<connection>
<GID>706</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-182,42,-182</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-179,40,-179</points>
<connection>
<GID>708</GID>
<name>OUT</name></connection>
<connection>
<GID>707</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-182,130,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-178,134,-178</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-169,130,-169</points>
<connection>
<GID>709</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-182,145,-182</points>
<intersection>130 0</intersection>
<intersection>145 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>145,-182.5,145,-182</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>-182 4</intersection></vsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,-179.5,143,-179.5</points>
<connection>
<GID>710</GID>
<name>ENABLE_0</name></connection>
<intersection>140 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>140,-179.5,140,-179</points>
<connection>
<GID>711</GID>
<name>OUT</name></connection>
<intersection>-179.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-182,95,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-178,99,-178</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-169,95,-169</points>
<connection>
<GID>712</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95,-182,110,-182</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-179,108,-179</points>
<connection>
<GID>714</GID>
<name>OUT</name></connection>
<connection>
<GID>713</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-182,199.5,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-178,203.5,-178</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197.5,-169,199.5,-169</points>
<connection>
<GID>715</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199.5,-182,214.5,-182</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-179,212.5,-179</points>
<connection>
<GID>717</GID>
<name>OUT</name></connection>
<connection>
<GID>716</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-182,164.5,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-178,168.5,-178</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-169,164.5,-169</points>
<connection>
<GID>718</GID>
<name>OUT_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-182,179.5,-182</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-179,177.5,-179</points>
<connection>
<GID>720</GID>
<name>OUT</name></connection>
<connection>
<GID>719</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-182,267.5,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-178,271.5,-178</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-169,267.5,-169</points>
<connection>
<GID>721</GID>
<name>OUT_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>267.5,-182,282.5,-182</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-179,280.5,-179</points>
<connection>
<GID>723</GID>
<name>OUT</name></connection>
<connection>
<GID>722</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-182,232.5,-169</points>
<intersection>-182 4</intersection>
<intersection>-178 1</intersection>
<intersection>-169 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,-178,236.5,-178</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230.5,-169,232.5,-169</points>
<connection>
<GID>724</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>232.5,-182,247.5,-182</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,-179,245.5,-179</points>
<connection>
<GID>726</GID>
<name>OUT</name></connection>
<connection>
<GID>725</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-180,271.5,-180</points>
<connection>
<GID>723</GID>
<name>IN_1</name></connection>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<connection>
<GID>717</GID>
<name>IN_1</name></connection>
<connection>
<GID>720</GID>
<name>IN_1</name></connection>
<connection>
<GID>711</GID>
<name>IN_1</name></connection>
<connection>
<GID>714</GID>
<name>IN_1</name></connection>
<connection>
<GID>705</GID>
<name>IN_1</name></connection>
<connection>
<GID>728</GID>
<name>OUT_0</name></connection>
<connection>
<GID>708</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-172,259.5,-172</points>
<connection>
<GID>721</GID>
<name>clock</name></connection>
<connection>
<GID>724</GID>
<name>clock</name></connection>
<connection>
<GID>715</GID>
<name>clock</name></connection>
<connection>
<GID>718</GID>
<name>clock</name></connection>
<connection>
<GID>709</GID>
<name>clock</name></connection>
<connection>
<GID>712</GID>
<name>clock</name></connection>
<connection>
<GID>703</GID>
<name>clock</name></connection>
<connection>
<GID>727</GID>
<name>OUT</name></connection>
<connection>
<GID>706</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-178,-84,-93.5</points>
<connection>
<GID>748</GID>
<name>OUT_0</name></connection>
<intersection>-178 2</intersection>
<intersection>-171 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84,-171,0,-171</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-84,-178,6,-178</points>
<connection>
<GID>728</GID>
<name>ENABLE_0</name></connection>
<intersection>-84 0</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-197.5,14.5,-6</points>
<connection>
<GID>729</GID>
<name>N_in1</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<intersection>-169 10</intersection>
<intersection>-146.5 9</intersection>
<intersection>-123 8</intersection>
<intersection>-98.5 7</intersection>
<intersection>-74 6</intersection>
<intersection>-50.5 5</intersection>
<intersection>-30 4</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-11,18,-11</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-30,19,-30</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-50.5,19.5,-50.5</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>14.5,-74,19,-74</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>14.5,-98.5,19,-98.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>14.5,-123,19,-123</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>14.5,-146.5,19.5,-146.5</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14.5,-169,19,-169</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-192.5,45,-1</points>
<connection>
<GID>730</GID>
<name>N_in1</name></connection>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<intersection>-176.5 6</intersection>
<intersection>-154 7</intersection>
<intersection>-130.5 8</intersection>
<intersection>-106 9</intersection>
<intersection>-81.5 10</intersection>
<intersection>-58 11</intersection>
<intersection>-37.5 12</intersection>
<intersection>-18.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>42,-176.5,45,-176.5</points>
<connection>
<GID>707</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>42.5,-154,45,-154</points>
<connection>
<GID>681</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>42,-130.5,45,-130.5</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42,-106,45,-106</points>
<connection>
<GID>629</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>42,-81.5,45,-81.5</points>
<connection>
<GID>603</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>42.5,-58,45,-58</points>
<connection>
<GID>577</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>42,-37.5,45,-37.5</points>
<connection>
<GID>551</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>41,-18.5,45,-18.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-197.5,50,-6</points>
<connection>
<GID>731</GID>
<name>N_in1</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<intersection>-169 10</intersection>
<intersection>-146.5 9</intersection>
<intersection>-123 8</intersection>
<intersection>-98.5 7</intersection>
<intersection>-74 6</intersection>
<intersection>-50.5 5</intersection>
<intersection>-30 4</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>50,-11,53,-11</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50,-30,54,-30</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>50,-50.5,54.5,-50.5</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>50,-74,54,-74</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>50,-98.5,54,-98.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>50,-123,54,-123</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>50,-146.5,54.5,-146.5</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>50,-169,54,-169</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-193,80,-1</points>
<connection>
<GID>732</GID>
<name>N_in1</name></connection>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<intersection>-176.5 6</intersection>
<intersection>-154 7</intersection>
<intersection>-130.5 8</intersection>
<intersection>-106 9</intersection>
<intersection>-81.5 10</intersection>
<intersection>-58 11</intersection>
<intersection>-37.5 12</intersection>
<intersection>-18.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-176.5,80,-176.5</points>
<connection>
<GID>704</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>77.5,-154,80,-154</points>
<connection>
<GID>678</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>77,-130.5,80,-130.5</points>
<connection>
<GID>652</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-106,80,-106</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>77,-81.5,80,-81.5</points>
<connection>
<GID>600</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>77.5,-58,80,-58</points>
<connection>
<GID>574</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>77,-37.5,80,-37.5</points>
<connection>
<GID>548</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>76,-18.5,80,-18.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-197.5,84,-6</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>733</GID>
<name>N_in1</name></connection>
<intersection>-169 3</intersection>
<intersection>-146.5 4</intersection>
<intersection>-123 5</intersection>
<intersection>-98.5 6</intersection>
<intersection>-74 7</intersection>
<intersection>-50.5 11</intersection>
<intersection>-30 9</intersection>
<intersection>-11 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-169,87,-169</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>84,-146.5,87.5,-146.5</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>84,-123,87,-123</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>84,-98.5,87,-98.5</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84,-74,87,-74</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>84,-30,87,-30</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84,-11,86,-11</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>84,-50.5,87.5,-50.5</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-192.5,115,-1</points>
<connection>
<GID>734</GID>
<name>N_in1</name></connection>
<connection>
<GID>65</GID>
<name>N_in0</name></connection>
<intersection>-176.5 13</intersection>
<intersection>-154 12</intersection>
<intersection>-130.5 11</intersection>
<intersection>-106 10</intersection>
<intersection>-81.5 9</intersection>
<intersection>-58 8</intersection>
<intersection>-37.5 7</intersection>
<intersection>-18.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109,-18.5,115,-18.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>110,-37.5,115,-37.5</points>
<connection>
<GID>557</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>110.5,-58,115,-58</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>110,-81.5,115,-81.5</points>
<connection>
<GID>609</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>110,-106,115,-106</points>
<connection>
<GID>635</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>110,-130.5,115,-130.5</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>110.5,-154,115,-154</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>110,-176.5,115,-176.5</points>
<connection>
<GID>713</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-197.5,118,-6</points>
<connection>
<GID>735</GID>
<name>N_in1</name></connection>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<intersection>-169 10</intersection>
<intersection>-146.5 9</intersection>
<intersection>-123 8</intersection>
<intersection>-98.5 7</intersection>
<intersection>-74 6</intersection>
<intersection>-50.5 5</intersection>
<intersection>-30 4</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,-11,121,-11</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>118,-30,122,-30</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>118,-50.5,122.5,-50.5</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>118,-74,122,-74</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>118,-98.5,122,-98.5</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118,-123,122,-123</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>118,-146.5,122.5,-146.5</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>118,-169,122,-169</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-192.5,150,-1</points>
<connection>
<GID>736</GID>
<name>N_in1</name></connection>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<intersection>-177 6</intersection>
<intersection>-154.5 7</intersection>
<intersection>-131 8</intersection>
<intersection>-106.5 9</intersection>
<intersection>-82 10</intersection>
<intersection>-58 11</intersection>
<intersection>-37 12</intersection>
<intersection>-18.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>145,-177,150,-177</points>
<connection>
<GID>710</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>145.5,-154.5,150,-154.5</points>
<intersection>145.5 19</intersection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>145,-131,150,-131</points>
<connection>
<GID>658</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>145.5,-106.5,150,-106.5</points>
<intersection>145.5 17</intersection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>145,-82,150,-82</points>
<intersection>145 16</intersection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>145.5,-58,150,-58</points>
<connection>
<GID>580</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>145,-37,150,-37</points>
<intersection>145 15</intersection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>144,-18.5,150,-18.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>145,-37.5,145,-37</points>
<connection>
<GID>554</GID>
<name>OUT_0</name></connection>
<intersection>-37 12</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>145,-82,145,-81.5</points>
<connection>
<GID>606</GID>
<name>OUT_0</name></connection>
<intersection>-82 10</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>145.5,-106.5,145.5,-106</points>
<connection>
<GID>632</GID>
<name>OUT_0</name></connection>
<intersection>-106.5 9</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>145.5,-154.5,145.5,-154</points>
<connection>
<GID>684</GID>
<name>OUT_0</name></connection>
<intersection>-154.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-197.5,153,-6</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<connection>
<GID>737</GID>
<name>N_in1</name></connection>
<intersection>-169 3</intersection>
<intersection>-146.5 4</intersection>
<intersection>-123 5</intersection>
<intersection>-98.5 6</intersection>
<intersection>-74 7</intersection>
<intersection>-50.5 8</intersection>
<intersection>-30 9</intersection>
<intersection>-11 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>153,-169,156.5,-169</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>153,-146.5,157,-146.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>153,-123,156.5,-123</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>153,-98.5,156.5,-98.5</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>153,-74,156.5,-74</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>153,-50.5,157,-50.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>153,-30,156.5,-30</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>153,-11,155.5,-11</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-192,184,-1</points>
<connection>
<GID>738</GID>
<name>N_in1</name></connection>
<connection>
<GID>69</GID>
<name>N_in0</name></connection>
<intersection>-176.5 13</intersection>
<intersection>-154 12</intersection>
<intersection>-130.5 11</intersection>
<intersection>-106 10</intersection>
<intersection>-81.5 9</intersection>
<intersection>-58 8</intersection>
<intersection>-37.5 7</intersection>
<intersection>-18.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>178.5,-18.5,184,-18.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>179.5,-37.5,184,-37.5</points>
<connection>
<GID>563</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>180,-58,184,-58</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>179.5,-81.5,184,-81.5</points>
<connection>
<GID>615</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>179.5,-106,184,-106</points>
<connection>
<GID>641</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>179.5,-130.5,184,-130.5</points>
<connection>
<GID>667</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>180,-154,184,-154</points>
<connection>
<GID>693</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>179.5,-176.5,184,-176.5</points>
<connection>
<GID>719</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-197.5,187,-6</points>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<connection>
<GID>739</GID>
<name>N_in1</name></connection>
<intersection>-169 10</intersection>
<intersection>-146.5 9</intersection>
<intersection>-123 8</intersection>
<intersection>-98.5 7</intersection>
<intersection>-74 6</intersection>
<intersection>-50.5 5</intersection>
<intersection>-30 4</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187,-11,190.5,-11</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>187,-30,191.5,-30</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>187,-50.5,192,-50.5</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>187,-74,191.5,-74</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>187,-98.5,191.5,-98.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187,-123,191.5,-123</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>187,-146.5,192,-146.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>187,-169,191.5,-169</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-192.5,219,-1</points>
<connection>
<GID>740</GID>
<name>N_in1</name></connection>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<intersection>-176.5 6</intersection>
<intersection>-154 7</intersection>
<intersection>-130.5 8</intersection>
<intersection>-106 9</intersection>
<intersection>-81.5 10</intersection>
<intersection>-58 11</intersection>
<intersection>-37.5 12</intersection>
<intersection>-18.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>214.5,-176.5,219,-176.5</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>215,-154,219,-154</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>214.5,-130.5,219,-130.5</points>
<connection>
<GID>664</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>214.5,-106,219,-106</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>214.5,-81.5,219,-81.5</points>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>215,-58,219,-58</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>214.5,-37.5,219,-37.5</points>
<connection>
<GID>560</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>213.5,-18.5,219,-18.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-197.5,222,-6</points>
<connection>
<GID>72</GID>
<name>N_in0</name></connection>
<connection>
<GID>741</GID>
<name>N_in1</name></connection>
<intersection>-169 3</intersection>
<intersection>-146.5 4</intersection>
<intersection>-123 5</intersection>
<intersection>-98.5 6</intersection>
<intersection>-74 7</intersection>
<intersection>-50.5 8</intersection>
<intersection>-30 9</intersection>
<intersection>-11 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>222,-169,224.5,-169</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>222,-146.5,225,-146.5</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>222,-123,224.5,-123</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>222,-98.5,224.5,-98.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>222,-74,224.5,-74</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>222,-50.5,225,-50.5</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>222,-30,224.5,-30</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>222,-11,223.5,-11</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-192,251,-1</points>
<connection>
<GID>73</GID>
<name>N_in0</name></connection>
<connection>
<GID>742</GID>
<name>N_in1</name></connection>
<intersection>-176.5 15</intersection>
<intersection>-154 14</intersection>
<intersection>-130.5 13</intersection>
<intersection>-106 12</intersection>
<intersection>-81.5 11</intersection>
<intersection>-58 10</intersection>
<intersection>-37.5 9</intersection>
<intersection>-18.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>246.5,-18.5,251,-18.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>247.5,-37.5,251,-37.5</points>
<connection>
<GID>569</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>248,-58,251,-58</points>
<connection>
<GID>595</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>247.5,-81.5,251,-81.5</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>247.5,-106,251,-106</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>247.5,-130.5,251,-130.5</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>248,-154,251,-154</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>247.5,-176.5,251,-176.5</points>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,-197.5,256,-6</points>
<connection>
<GID>743</GID>
<name>N_in1</name></connection>
<connection>
<GID>74</GID>
<name>N_in0</name></connection>
<intersection>-169 10</intersection>
<intersection>-146.5 9</intersection>
<intersection>-123 8</intersection>
<intersection>-98.5 7</intersection>
<intersection>-74 6</intersection>
<intersection>-50.5 5</intersection>
<intersection>-30 4</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>256,-11,258.5,-11</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>256,-30,259.5,-30</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>256,-50.5,260,-50.5</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256,-74,259.5,-74</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>256,-98.5,259.5,-98.5</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>256,-123,259.5,-123</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>256,-146.5,260,-146.5</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>256,-169,259.5,-169</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-192,288,-1</points>
<connection>
<GID>744</GID>
<name>N_in1</name></connection>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<intersection>-176.5 6</intersection>
<intersection>-154 7</intersection>
<intersection>-130.5 8</intersection>
<intersection>-106 9</intersection>
<intersection>-81.5 10</intersection>
<intersection>-58 11</intersection>
<intersection>-37.5 12</intersection>
<intersection>-18.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>282.5,-176.5,288,-176.5</points>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>283,-154,288,-154</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>282.5,-130.5,288,-130.5</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>282.5,-106,288,-106</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>282.5,-81.5,288,-81.5</points>
<connection>
<GID>618</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>283,-58,288,-58</points>
<connection>
<GID>592</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>282.5,-37.5,288,-37.5</points>
<connection>
<GID>566</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>281.5,-18.5,288,-18.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>288 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-43,62,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-39,66,-39</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-30,62,-30</points>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62,-43,77,-43</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-40,75,-40</points>
<connection>
<GID>549</GID>
<name>OUT</name></connection>
<connection>
<GID>548</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-43,27,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-39,31,-39</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-30,27,-30</points>
<connection>
<GID>550</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>27,-43,42,-43</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-40,40,-40</points>
<connection>
<GID>552</GID>
<name>OUT</name></connection>
<connection>
<GID>551</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-43,130,-30</points>
<intersection>-43 4</intersection>
<intersection>-39 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-39,134,-39</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-30,130,-30</points>
<connection>
<GID>553</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-43,145,-43</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 9></circuit>