<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-62.8331,50.2757,234.159,-96.5219</PageViewport>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>5,0</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>17,0</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>78.5,-80</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>15 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>10</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>88.5,-79.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>19 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-16</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>17,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_FULLADDER_1BIT</type>
<position>14.5,-27</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_B_0</ID>21 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>carry_in</ID>124 </input>
<output>
<ID>carry_out</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>5.5,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AE_DFF_LOW</type>
<position>18.5,-37</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>249</ID>
<type>GA_LED</type>
<position>24.5,-47</position>
<input>
<ID>N_in2</ID>15 </input>
<input>
<ID>N_in3</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_TOGGLE</type>
<position>-5,-38</position>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>28,0</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>39.5,0</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37,-27</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_B_0</ID>27 </input>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>carry_in</ID>123 </input>
<output>
<ID>carry_out</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>39.5,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>AE_DFF_LOW</type>
<position>41,-37</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>28,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>GA_LED</type>
<position>47,-47</position>
<input>
<ID>N_in2</ID>14 </input>
<input>
<ID>N_in3</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AE_DFF_LOW</type>
<position>31.5,-15</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>27 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_DFF_LOW</type>
<position>42.5,-15</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>49,0</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_TOGGLE</type>
<position>60.5,0</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_FULLADDER_1BIT</type>
<position>58,-27</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_B_0</ID>33 </input>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>carry_in</ID>122 </input>
<output>
<ID>carry_out</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>60.5,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AE_DFF_LOW</type>
<position>62,-37</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>36 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>49,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>GA_LED</type>
<position>68,-47</position>
<input>
<ID>N_in2</ID>13 </input>
<input>
<ID>N_in3</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>AA_TOGGLE</type>
<position>71.5,0</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_TOGGLE</type>
<position>83,0</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_FULLADDER_1BIT</type>
<position>80.5,-27</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_B_0</ID>39 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>carry_in</ID>121 </input>
<output>
<ID>carry_out</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>83,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>AE_DFF_LOW</type>
<position>84.5,-37</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>42 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_LABEL</type>
<position>71.5,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>GA_LED</type>
<position>90.5,-47</position>
<input>
<ID>N_in2</ID>12 </input>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>AE_DFF_LOW</type>
<position>75,-15</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>276</ID>
<type>AE_DFF_LOW</type>
<position>86,-15</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>277</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-15</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>33 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>278</ID>
<type>AE_DFF_LOW</type>
<position>63.5,-15</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_TOGGLE</type>
<position>91.5,0</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_TOGGLE</type>
<position>103,0</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_FULLADDER_1BIT</type>
<position>100.5,-27</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_B_0</ID>45 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>carry_in</ID>120 </input>
<output>
<ID>carry_out</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_LABEL</type>
<position>103,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>AE_DFF_LOW</type>
<position>104.5,-37</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>91.5,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>GA_LED</type>
<position>110.5,-47</position>
<input>
<ID>N_in2</ID>19 </input>
<input>
<ID>N_in3</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>AA_TOGGLE</type>
<position>114,0</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_TOGGLE</type>
<position>125.5,0</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_DFF_LOW</type>
<position>9,-15</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>21 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_FULLADDER_1BIT</type>
<position>123,-27</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>carry_in</ID>119 </input>
<output>
<ID>carry_out</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>125.5,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>20,-15</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_DFF_LOW</type>
<position>127,-37</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>114,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>GA_LED</type>
<position>133,-47</position>
<input>
<ID>N_in2</ID>18 </input>
<input>
<ID>N_in3</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AE_DFF_LOW</type>
<position>117.5,-15</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-15</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_TOGGLE</type>
<position>135,0</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_TOGGLE</type>
<position>146.5,0</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_FULLADDER_1BIT</type>
<position>144,-27</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_B_0</ID>57 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>carry_in</ID>118 </input>
<output>
<ID>carry_out</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_LABEL</type>
<position>146.5,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>AE_DFF_LOW</type>
<position>148,-37</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>61 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_LABEL</type>
<position>135,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>GA_LED</type>
<position>154,-47</position>
<input>
<ID>N_in2</ID>17 </input>
<input>
<ID>N_in3</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>AA_TOGGLE</type>
<position>157.5,0</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_TOGGLE</type>
<position>169,0</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_FULLADDER_1BIT</type>
<position>166.5,-27</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_B_0</ID>64 </input>
<output>
<ID>OUT_0</ID>66 </output>
<output>
<ID>carry_out</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_LABEL</type>
<position>169,2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>170.5,-37</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>107 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_LABEL</type>
<position>157,2.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>308</ID>
<type>GA_LED</type>
<position>176.5,-47</position>
<input>
<ID>N_in2</ID>16 </input>
<input>
<ID>N_in3</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>AE_DFF_LOW</type>
<position>161,-15</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>310</ID>
<type>AE_DFF_LOW</type>
<position>172,-15</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>311</ID>
<type>AE_DFF_LOW</type>
<position>138.5,-15</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>57 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>312</ID>
<type>AE_DFF_LOW</type>
<position>149.5,-15</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>313</ID>
<type>AE_DFF_LOW</type>
<position>95,-15</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>314</ID>
<type>AE_DFF_LOW</type>
<position>106,-15</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>320</ID>
<type>GA_LED</type>
<position>-9,-31</position>
<input>
<ID>N_in1</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>AE_DFF_LOW</type>
<position>-1,-29</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>130 </output>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>-10,-15.5</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>AA_LABEL</type>
<position>-11.5,-37.5</position>
<gparam>LABEL_TEXT Collect</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>AA_LABEL</type>
<position>-14.5,-30.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>330</ID>
<type>AA_LABEL</type>
<position>132,24</position>
<gparam>LABEL_TEXT X 8-bit value = 10001100</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>AA_LABEL</type>
<position>132,19.5</position>
<gparam>LABEL_TEXT Y 8-bit value = 01000011</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>334</ID>
<type>AA_LABEL</type>
<position>77,-56</position>
<gparam>LABEL_TEXT Out-put  8-bit value = 11001111</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>-40,28</position>
<gparam>LABEL_TEXT SECOND</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-13,5,-2</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-13,6,-13</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-13,17,-2</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-81,73,-48</points>
<intersection>-81 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-81,75.5,-81</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-48,90.5,-48</points>
<connection>
<GID>274</GID>
<name>N_in2</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-80,68,-48</points>
<connection>
<GID>267</GID>
<name>N_in2</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-80,75.5,-80</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-79,47,-48</points>
<connection>
<GID>258</GID>
<name>N_in2</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-79,75.5,-79</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-78,24.5,-48</points>
<connection>
<GID>249</GID>
<name>N_in2</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-78,75.5,-78</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-58.5,176.5,-48</points>
<connection>
<GID>308</GID>
<name>N_in2</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-58.5,176.5,-58.5</points>
<intersection>82.5 2</intersection>
<intersection>176.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>82.5,-80.5,82.5,-58.5</points>
<intersection>-80.5 3</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82.5,-80.5,85.5,-80.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>82.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-61,154,-48</points>
<connection>
<GID>301</GID>
<name>N_in2</name></connection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-61,154,-61</points>
<intersection>85.5 2</intersection>
<intersection>154 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>85.5,-79.5,85.5,-61</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-63.5,133,-48</points>
<connection>
<GID>292</GID>
<name>N_in2</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-63.5,133,-63.5</points>
<intersection>83.5 2</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83.5,-78.5,83.5,-63.5</points>
<intersection>-78.5 3</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83.5,-78.5,85.5,-78.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>83.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-67,110.5,-48</points>
<connection>
<GID>285</GID>
<name>N_in2</name></connection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-67,110.5,-67</points>
<intersection>81 2</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>81,-77.5,81,-67</points>
<intersection>-77.5 3</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81,-77.5,85.5,-77.5</points>
<connection>
<GID>10</GID>
<name>IN_3</name></connection>
<intersection>81 2</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-24,13.5,-13</points>
<connection>
<GID>245</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-13,13.5,-13</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-24,23.5,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>15.5,-24,23.5,-24</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>23,-13,23.5,-13</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-35,14.5,-30</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-35,15.5,-35</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-46,24.5,-35</points>
<connection>
<GID>249</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-35,24.5,-35</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-13,28,-2</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-13,28.5,-13</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-13,39.5,-2</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-24,36,-13</points>
<connection>
<GID>254</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-13,36,-13</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-24,46,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>38,-24,46,-24</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>45.5,-13,46,-13</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-35,37,-30</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-35,38,-35</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-46,47,-35</points>
<connection>
<GID>258</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-35,47,-35</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-13,49,-2</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-13,49.5,-13</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-13,60.5,-2</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-24,57,-13</points>
<connection>
<GID>263</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-13,57,-13</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-24,67,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59,-24,67,-24</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>66.5,-13,67,-13</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-35,58,-30</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-35,59,-35</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-46,68,-35</points>
<connection>
<GID>267</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-35,68,-35</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-13,71.5,-2</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-13,72,-13</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-13,83,-2</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-24,79.5,-13</points>
<connection>
<GID>270</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-13,79.5,-13</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-24,89.5,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-24,89.5,-24</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>89,-13,89.5,-13</points>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-35,80.5,-30</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-35,81.5,-35</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-46,90.5,-35</points>
<connection>
<GID>274</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-35,90.5,-35</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-13,91.5,-2</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-13,92,-13</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-13,103,-2</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-24,99.5,-13</points>
<connection>
<GID>281</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-13,99.5,-13</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-24,109.5,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>101.5,-24,109.5,-24</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>109,-13,109.5,-13</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-35,100.5,-30</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-35,101.5,-35</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-46,110.5,-35</points>
<connection>
<GID>285</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-35,110.5,-35</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-13,114,-2</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-13,114.5,-13</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-13,125.5,-2</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-24,122,-13</points>
<connection>
<GID>288</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-13,122,-13</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-24,132,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>124,-24,132,-24</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>131.5,-13,132,-13</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-35,123,-30</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-35,124,-35</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-46,133,-35</points>
<connection>
<GID>292</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-35,133,-35</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-13,135,-2</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-13,135.5,-13</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-13,146.5,-2</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-24,143,-13</points>
<connection>
<GID>297</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-13,143,-13</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-24,153,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>145,-24,153,-24</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>152.5,-13,153,-13</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-35,144,-30</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-35,145,-35</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-46,154,-35</points>
<connection>
<GID>301</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-35,154,-35</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-13,157.5,-2</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-13,158,-13</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-13,169,-2</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-24,165.5,-13</points>
<connection>
<GID>304</GID>
<name>IN_B_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164,-13,165.5,-13</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-24,175.5,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>167.5,-24,175.5,-24</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>175,-13,175.5,-13</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-35,166.5,-30</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-35,167.5,-35</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-46,176.5,-35</points>
<connection>
<GID>308</GID>
<name>N_in3</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,-35,176.5,-35</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-16,169,-16</points>
<connection>
<GID>310</GID>
<name>clock</name></connection>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<connection>
<GID>294</GID>
<name>clock</name></connection>
<connection>
<GID>293</GID>
<name>clock</name></connection>
<connection>
<GID>314</GID>
<name>clock</name></connection>
<connection>
<GID>313</GID>
<name>clock</name></connection>
<connection>
<GID>276</GID>
<name>clock</name></connection>
<connection>
<GID>275</GID>
<name>clock</name></connection>
<connection>
<GID>278</GID>
<name>clock</name></connection>
<connection>
<GID>277</GID>
<name>clock</name></connection>
<connection>
<GID>260</GID>
<name>clock</name></connection>
<connection>
<GID>259</GID>
<name>clock</name></connection>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3,-38,167.5,-38</points>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<connection>
<GID>299</GID>
<name>clock</name></connection>
<connection>
<GID>290</GID>
<name>clock</name></connection>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<connection>
<GID>272</GID>
<name>clock</name></connection>
<connection>
<GID>265</GID>
<name>clock</name></connection>
<connection>
<GID>256</GID>
<name>clock</name></connection>
<connection>
<GID>247</GID>
<name>clock</name></connection>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>3.5 37</intersection></hsegment>
<vsegment>
<ID>37</ID>
<points>3.5,-38,3.5,-28</points>
<intersection>-38 1</intersection>
<intersection>-28 38</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>2,-28,3.5,-28</points>
<connection>
<GID>322</GID>
<name>clock</name></connection>
<intersection>3.5 37</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148,-27,162.5,-27</points>
<connection>
<GID>297</GID>
<name>carry_in</name></connection>
<connection>
<GID>304</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127,-27,140,-27</points>
<connection>
<GID>288</GID>
<name>carry_in</name></connection>
<connection>
<GID>297</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-27,119,-27</points>
<connection>
<GID>281</GID>
<name>carry_in</name></connection>
<connection>
<GID>288</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-27,96.5,-27</points>
<connection>
<GID>270</GID>
<name>carry_in</name></connection>
<connection>
<GID>281</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-27,76.5,-27</points>
<connection>
<GID>263</GID>
<name>carry_in</name></connection>
<connection>
<GID>270</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-27,54,-27</points>
<connection>
<GID>254</GID>
<name>carry_in</name></connection>
<connection>
<GID>263</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-27,33,-27</points>
<connection>
<GID>245</GID>
<name>carry_in</name></connection>
<connection>
<GID>254</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-31,6,-27</points>
<intersection>-31 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-31,6,-31</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-27,10.5,-27</points>
<connection>
<GID>245</GID>
<name>carry_out</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-31,-4,-31</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<connection>
<GID>320</GID>
<name>N_in1</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>12.4661,-6.9855,137.76,-68.9159</PageViewport>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>93,-14.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>100.5,-14.5</position>
<gparam>LABEL_TEXT X2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>BA_TRI_STATE</type>
<position>93,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>BA_TRI_STATE</type>
<position>100.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_FULLADDER_1BIT</type>
<position>111,-36</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_B_0</ID>100 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>carry_in</ID>115 </input>
<output>
<ID>carry_out</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>GA_LED</type>
<position>111,-43</position>
<input>
<ID>N_in3</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_TOGGLE</type>
<position>107.5,-18</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_TOGGLE</type>
<position>115,-18</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>107.5,-14.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_LABEL</type>
<position>115,-14.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>BA_TRI_STATE</type>
<position>107.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>204</ID>
<type>BA_TRI_STATE</type>
<position>115,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_FULLADDER_1BIT</type>
<position>124.5,-36</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_B_0</ID>105 </input>
<output>
<ID>OUT_0</ID>101 </output>
<output>
<ID>carry_out</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>206</ID>
<type>GA_LED</type>
<position>124.5,-43</position>
<input>
<ID>N_in3</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>121,-18</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_TOGGLE</type>
<position>128.5,-18</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>121,-14.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>128.5,-14.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>BA_TRI_STATE</type>
<position>121,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>212</ID>
<type>BA_TRI_STATE</type>
<position>128.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>133,-49</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>220</ID>
<type>GA_LED</type>
<position>19,-50.5</position>
<input>
<ID>N_in3</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>82,0.5</position>
<gparam>LABEL_TEXT X Input Data</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>133,-51.5</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>18.5,-53</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_LABEL</type>
<position>110,0.5</position>
<gparam>LABEL_TEXT 8-bit Data = 10101011</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>110,-3.5</position>
<gparam>LABEL_TEXT 8-bit Data = 11010101</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>73.5,-47.5</position>
<gparam>LABEL_TEXT SUM   = 10000000</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>82,-3.5</position>
<gparam>LABEL_TEXT Y Input Data</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>19.5,-57</position>
<gparam>LABEL_TEXT Carry = 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_FULLADDER_1BIT</type>
<position>25,-36</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_B_0</ID>70 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>carry_in</ID>109 </input>
<output>
<ID>carry_out</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>25,-43</position>
<input>
<ID>N_in3</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>21.5,-18</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>29,-18</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>21.5,-14.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>29,-14.5</position>
<gparam>LABEL_TEXT X7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>BA_TRI_STATE</type>
<position>21.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>BA_TRI_STATE</type>
<position>29,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_FULLADDER_1BIT</type>
<position>40,-36</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_B_0</ID>75 </input>
<output>
<ID>OUT_0</ID>71 </output>
<input>
<ID>carry_in</ID>110 </input>
<output>
<ID>carry_out</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>40,-43</position>
<input>
<ID>N_in3</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>36.5,-18</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_TOGGLE</type>
<position>44,-18</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>36.5,-14.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>44,-14.5</position>
<gparam>LABEL_TEXT X6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>BA_TRI_STATE</type>
<position>36.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>BA_TRI_STATE</type>
<position>44,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_FULLADDER_1BIT</type>
<position>54.5,-36</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_B_0</ID>80 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>carry_in</ID>111 </input>
<output>
<ID>carry_out</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>GA_LED</type>
<position>54.5,-43</position>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>51,-18</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>58.5,-18</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>51,-14.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>23.5,-9.5</position>
<gparam>LABEL_TEXT FIRST</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>58.5,-14.5</position>
<gparam>LABEL_TEXT X5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>BA_TRI_STATE</type>
<position>51,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>172</ID>
<type>BA_TRI_STATE</type>
<position>58.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_FULLADDER_1BIT</type>
<position>68,-36</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_B_0</ID>85 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>carry_in</ID>112 </input>
<output>
<ID>carry_out</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>68,-43</position>
<input>
<ID>N_in3</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_TOGGLE</type>
<position>64.5,-18</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_TOGGLE</type>
<position>72,-18</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>64.5,-14.5</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>72,-14.5</position>
<gparam>LABEL_TEXT X4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>BA_TRI_STATE</type>
<position>64.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>BA_TRI_STATE</type>
<position>72,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_FULLADDER_1BIT</type>
<position>81.5,-36</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_B_0</ID>90 </input>
<output>
<ID>OUT_0</ID>86 </output>
<input>
<ID>carry_in</ID>113 </input>
<output>
<ID>carry_out</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>81.5,-43</position>
<input>
<ID>N_in3</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>78,-18</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_TOGGLE</type>
<position>85.5,-18</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>78,-14.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>85.5,-14.5</position>
<gparam>LABEL_TEXT X3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>BA_TRI_STATE</type>
<position>78,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>188</ID>
<type>BA_TRI_STATE</type>
<position>85.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_FULLADDER_1BIT</type>
<position>96.5,-36</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_B_0</ID>95 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>carry_in</ID>114 </input>
<output>
<ID>carry_out</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>190</ID>
<type>GA_LED</type>
<position>96.5,-43</position>
<input>
<ID>N_in3</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>93,-18</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>100.5,-18</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-42,25,-39</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>96</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-26,21.5,-20</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-26,29,-20</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-33,26,-32</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,-32,29,-31.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26,-32,29,-32</points>
<intersection>26 0</intersection>
<intersection>29 1</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-33,24,-32</points>
<connection>
<GID>79</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>21.5,-32,21.5,-31.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-32,24,-32</points>
<intersection>21.5 1</intersection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-42,40,-39</points>
<connection>
<GID>158</GID>
<name>N_in3</name></connection>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-26,36.5,-20</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-26,44,-20</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-33,41,-32</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44,-32,44,-31.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41,-32,44,-32</points>
<intersection>41 0</intersection>
<intersection>44 1</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-33,39,-32</points>
<connection>
<GID>157</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>36.5,-32,36.5,-31.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-32,39,-32</points>
<intersection>36.5 1</intersection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-42,54.5,-39</points>
<connection>
<GID>166</GID>
<name>N_in3</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-26,51,-20</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-26,58.5,-20</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-33,55.5,-32</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58.5,-32,58.5,-31.5</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-32,58.5,-32</points>
<intersection>55.5 0</intersection>
<intersection>58.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-33,53.5,-32</points>
<connection>
<GID>165</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51,-32,51,-31.5</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51,-32,53.5,-32</points>
<intersection>51 1</intersection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-42,68,-39</points>
<connection>
<GID>174</GID>
<name>N_in3</name></connection>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-26,64.5,-20</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-26,72,-20</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-33,69,-32</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72,-32,72,-31.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-32,72,-32</points>
<intersection>69 0</intersection>
<intersection>72 1</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-33,67,-32</points>
<connection>
<GID>173</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-32,64.5,-31.5</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-32,67,-32</points>
<intersection>64.5 1</intersection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-42,81.5,-39</points>
<connection>
<GID>182</GID>
<name>N_in3</name></connection>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-26,78,-20</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-26,85.5,-20</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-33,82.5,-32</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>85.5,-32,85.5,-31.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-32,85.5,-32</points>
<intersection>82.5 0</intersection>
<intersection>85.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-33,80.5,-32</points>
<connection>
<GID>181</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78,-32,78,-31.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-32,80.5,-32</points>
<intersection>78 1</intersection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-42,96.5,-39</points>
<connection>
<GID>190</GID>
<name>N_in3</name></connection>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-26,93,-20</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-26,100.5,-20</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<connection>
<GID>196</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-33,97.5,-32</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>100.5,-32,100.5,-31.5</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-32,100.5,-32</points>
<intersection>97.5 0</intersection>
<intersection>100.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-33,95.5,-32</points>
<connection>
<GID>189</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93,-32,93,-31.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>93,-32,95.5,-32</points>
<intersection>93 1</intersection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-42,111,-39</points>
<connection>
<GID>198</GID>
<name>N_in3</name></connection>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-26,107.5,-20</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-26,115,-20</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-33,112,-32</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>115,-32,115,-31.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112,-32,115,-32</points>
<intersection>112 0</intersection>
<intersection>115 1</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-33,110,-32</points>
<connection>
<GID>197</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>107.5,-32,107.5,-31.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-32,110,-32</points>
<intersection>107.5 1</intersection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-42,124.5,-39</points>
<connection>
<GID>206</GID>
<name>N_in3</name></connection>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-26,121,-20</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-26,128.5,-20</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-33,125.5,-32</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>128.5,-32,128.5,-31.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-32,128.5,-32</points>
<intersection>125.5 0</intersection>
<intersection>128.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-33,123.5,-32</points>
<connection>
<GID>205</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>121,-32,121,-31.5</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121,-32,123.5,-32</points>
<intersection>121 1</intersection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-29,133,-29</points>
<connection>
<GID>154</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>156</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>163</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>164</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>171</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>172</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>179</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>180</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>187</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>188</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>195</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>196</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>203</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>204</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>211</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>212</GID>
<name>ENABLE_0</name></connection>
<intersection>133 66</intersection></hsegment>
<vsegment>
<ID>66</ID>
<points>133,-47,133,-29</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-49.5,19,-36</points>
<connection>
<GID>220</GID>
<name>N_in3</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-36,21,-36</points>
<connection>
<GID>79</GID>
<name>carry_out</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-36,36,-36</points>
<connection>
<GID>79</GID>
<name>carry_in</name></connection>
<connection>
<GID>157</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-36,50.5,-36</points>
<connection>
<GID>157</GID>
<name>carry_in</name></connection>
<connection>
<GID>165</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-36,64,-36</points>
<connection>
<GID>165</GID>
<name>carry_in</name></connection>
<connection>
<GID>173</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-36,77.5,-36</points>
<connection>
<GID>173</GID>
<name>carry_in</name></connection>
<connection>
<GID>181</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-36,92.5,-36</points>
<connection>
<GID>181</GID>
<name>carry_in</name></connection>
<connection>
<GID>189</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-36,107,-36</points>
<connection>
<GID>189</GID>
<name>carry_in</name></connection>
<connection>
<GID>197</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-36,120.5,-36</points>
<connection>
<GID>197</GID>
<name>carry_in</name></connection>
<connection>
<GID>205</GID>
<name>carry_out</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>163.713,137.113,691.699,-123.86</PageViewport>
<gate>
<ID>12</ID>
<type>AI_XOR2</type>
<position>328,27.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR2</type>
<position>342,22</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>342,12.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AI_XOR2</type>
<position>286.5,22</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR2</type>
<position>352,9</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>286.5,12.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_OR2</type>
<position>296.5,9</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>246 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>GA_LED</type>
<position>293.5,22</position>
<input>
<ID>N_in0</ID>208 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_TOGGLE</type>
<position>253.5,31.5</position>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_TOGGLE</type>
<position>253.5,26.5</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>349,22</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_AND2</type>
<position>267.5,8</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>303,6.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>295.5,20</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>HA_JUNC_2</type>
<position>255,9</position>
<input>
<ID>N_in0</ID>213 </input>
<input>
<ID>N_in1</ID>206 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>308.5,31.5</position>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>229</ID>
<type>AI_XOR2</type>
<position>552.5,27</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>309,26.5</position>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>231</ID>
<type>AI_XOR2</type>
<position>566.5,21.5</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>323,8</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>566.5,12</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AI_XOR2</type>
<position>511,21.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>358.5,6.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>AE_OR2</type>
<position>576.5,8.5</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>511,12</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>239 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>351,20</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AE_OR2</type>
<position>521,8.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AI_XOR2</type>
<position>383,27.5</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>GA_LED</type>
<position>518,21.5</position>
<input>
<ID>N_in0</ID>240 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AI_XOR2</type>
<position>397,22</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>397,12.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_OR2</type>
<position>407,9</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_TOGGLE</type>
<position>478,31</position>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>404,22</position>
<input>
<ID>N_in0</ID>143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_TOGGLE</type>
<position>478,26</position>
<output>
<ID>OUT_0</ID>243 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>248</ID>
<type>GA_LED</type>
<position>573.5,21.5</position>
<input>
<ID>N_in0</ID>217 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>364,31.5</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>364,26.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>492,7.5</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND2</type>
<position>378,8</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>413.5,6.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>406,20</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AA_LABEL</type>
<position>527.5,6</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>AA_LABEL</type>
<position>520,19.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>HA_JUNC_2</type>
<position>479.5,8.5</position>
<input>
<ID>N_in0</ID>245 </input>
<input>
<ID>N_in1</ID>238 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AA_TOGGLE</type>
<position>533.5,31</position>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_TOGGLE</type>
<position>533.5,26</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_AND2</type>
<position>547.5,7.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_LABEL</type>
<position>583,6</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>AA_LABEL</type>
<position>575.5,19.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>AI_XOR2</type>
<position>607.5,27</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AI_XOR2</type>
<position>621.5,21.5</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AA_AND2</type>
<position>621.5,12</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_OR2</type>
<position>631.5,8.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>HA_JUNC_2</type>
<position>365.5,9</position>
<input>
<ID>N_in0</ID>197 </input>
<input>
<ID>N_in1</ID>141 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>GA_LED</type>
<position>628.5,21.5</position>
<input>
<ID>N_in0</ID>224 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AI_XOR2</type>
<position>217.5,27.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>GA_LED</type>
<position>637.5,8.5</position>
<input>
<ID>N_in0</ID>225 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AI_XOR2</type>
<position>231.5,22</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_TOGGLE</type>
<position>588.5,31</position>
<output>
<ID>OUT_0</ID>226 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>231.5,12.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_TOGGLE</type>
<position>588.5,26</position>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>146</ID>
<type>AE_OR2</type>
<position>241.5,9</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>602.5,7.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>238.5,22</position>
<input>
<ID>N_in0</ID>201 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>341</ID>
<type>AA_LABEL</type>
<position>638,6</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>198.5,31.5</position>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>342</ID>
<type>AA_LABEL</type>
<position>630.5,19.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>198.5,26.5</position>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>343</ID>
<type>HA_JUNC_2</type>
<position>590,8.5</position>
<input>
<ID>N_in0</ID>229 </input>
<input>
<ID>N_in1</ID>222 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>212.5,8</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>AI_XOR2</type>
<position>442,27</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>198.5,13.5</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>345</ID>
<type>AI_XOR2</type>
<position>456,21.5</position>
<input>
<ID>IN_0</ID>232 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>248,6.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>AA_AND2</type>
<position>456,12</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>240.5,20</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AE_OR2</type>
<position>466,8.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>GA_LED</type>
<position>463,21.5</position>
<input>
<ID>N_in0</ID>233 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AI_XOR2</type>
<position>272.5,27.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_TOGGLE</type>
<position>423,31</position>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_TOGGLE</type>
<position>423,26</position>
<output>
<ID>OUT_0</ID>235 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_AND2</type>
<position>437,7.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_LABEL</type>
<position>472.5,6</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>465,19.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>AI_XOR2</type>
<position>497,27</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>HA_JUNC_2</type>
<position>310,9</position>
<input>
<ID>N_in0</ID>246 </input>
<input>
<ID>N_in1</ID>133 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>359</ID>
<type>HA_JUNC_2</type>
<position>418.5,9</position>
<input>
<ID>N_in0</ID>247 </input>
<input>
<ID>N_in1</ID>231 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>361</ID>
<type>HA_JUNC_2</type>
<position>533,8.5</position>
<input>
<ID>N_in0</ID>248 </input>
<input>
<ID>N_in1</ID>215 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,9,364.5,9</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>142</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,10,236.5,12.5</points>
<intersection>10 1</intersection>
<intersection>12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,10,238.5,10</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>236.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234.5,12.5,236.5,12.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,21,228.5,21</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>227.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>227.5,13.5,227.5,21</points>
<intersection>13.5 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>200.5,13.5,228.5,13.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>227.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,27.5,225,27.5</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<intersection>225 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>225,11.5,225,27.5</points>
<intersection>11.5 5</intersection>
<intersection>23 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225,11.5,228.5,11.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>225 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>225,23,228.5,23</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>225 3</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,22,237.5,22</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<connection>
<GID>147</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,31.5,209.5,31.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,9,209.5,31.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>28.5 6</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>209.5,28.5,214.5,28.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>209.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>200.5,26.5,214.5,26.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>204.5,7,204.5,26.5</points>
<intersection>7 4</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>204.5,7,209.5,7</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215.5,8,238.5,8</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<connection>
<GID>146</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,10,291.5,12.5</points>
<intersection>10 1</intersection>
<intersection>12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,10,293.5,10</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>289.5,12.5,291.5,12.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>282.5,21,283.5,21</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>282.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>282.5,13.5,282.5,21</points>
<intersection>13.5 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256,13.5,283.5,13.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>256 7</intersection>
<intersection>282.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>256,9,256,13.5</points>
<connection>
<GID>227</GID>
<name>N_in1</name></connection>
<intersection>13.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>275.5,27.5,280,27.5</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>280 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>280,11.5,280,27.5</points>
<intersection>11.5 5</intersection>
<intersection>23 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>280,11.5,283.5,11.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>280 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>280,23,283.5,23</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>280 3</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,22,292.5,22</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<connection>
<GID>217</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>255.5,31.5,264.5,31.5</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>264.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>264.5,9,264.5,31.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>28.5 6</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>264.5,28.5,269.5,28.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>264.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>255.5,26.5,269.5,26.5</points>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>260 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>260,7,260,26.5</points>
<intersection>7 4</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260,7,264.5,7</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>260 3</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>270.5,8,293.5,8</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<connection>
<GID>215</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244.5,9,254,9</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<connection>
<GID>227</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,9.5,571.5,12</points>
<intersection>9.5 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571.5,9.5,573.5,9.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>571.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>569.5,12,571.5,12</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<intersection>571.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562.5,20.5,563.5,20.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>562.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>562.5,13,562.5,20.5</points>
<intersection>13 4</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>535.5,13,563.5,13</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>535.5 7</intersection>
<intersection>562.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>535.5,8.5,535.5,13</points>
<intersection>8.5 8</intersection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>534,8.5,535.5,8.5</points>
<connection>
<GID>361</GID>
<name>N_in1</name></connection>
<intersection>535.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>555.5,27,560,27</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>560 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>560,11,560,27</points>
<intersection>11 5</intersection>
<intersection>22.5 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>560,11,563.5,11</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>560 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>560,22.5,563.5,22.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>560 3</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>569.5,21.5,572.5,21.5</points>
<connection>
<GID>248</GID>
<name>N_in0</name></connection>
<connection>
<GID>231</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>535.5,31,544.5,31</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>544.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>544.5,8.5,544.5,31</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>28 6</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>544.5,28,549.5,28</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>544.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>535.5,26,549.5,26</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>540 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>540,6.5,540,26</points>
<intersection>6.5 4</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>540,6.5,544.5,6.5</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>540 3</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>550.5,7.5,573.5,7.5</points>
<connection>
<GID>321</GID>
<name>OUT</name></connection>
<connection>
<GID>238</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>626.5,9.5,626.5,12</points>
<intersection>9.5 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>626.5,9.5,628.5,9.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>626.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>624.5,12,626.5,12</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<intersection>626.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>617.5,20.5,618.5,20.5</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>617.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>617.5,13,617.5,20.5</points>
<intersection>13 4</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>591,13,618.5,13</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>591 7</intersection>
<intersection>617.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>591,8.5,591,13</points>
<connection>
<GID>343</GID>
<name>N_in1</name></connection>
<intersection>13 4</intersection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,27,615,27</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>615 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>615,11,615,27</points>
<intersection>11 5</intersection>
<intersection>22.5 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>615,11,618.5,11</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>615 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>615,22.5,618.5,22.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>615 3</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>624.5,21.5,627.5,21.5</points>
<connection>
<GID>336</GID>
<name>N_in0</name></connection>
<connection>
<GID>331</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>634.5,8.5,636.5,8.5</points>
<connection>
<GID>337</GID>
<name>N_in0</name></connection>
<connection>
<GID>335</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>590.5,31,599.5,31</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>599.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>599.5,8.5,599.5,31</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>28 6</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>599.5,28,604.5,28</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>599.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>590.5,26,604.5,26</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>595 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>595,6.5,595,26</points>
<intersection>6.5 4</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>595,6.5,599.5,6.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>595 3</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>605.5,7.5,628.5,7.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<connection>
<GID>335</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>579.5,8.5,589,8.5</points>
<connection>
<GID>343</GID>
<name>N_in0</name></connection>
<connection>
<GID>238</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461,9.5,461,12</points>
<intersection>9.5 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>461,9.5,463,9.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>461 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>459,12,461,12</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<intersection>461 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>452,20.5,453,20.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>452 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>452,13,452,20.5</points>
<intersection>13 4</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>419.5,13,453,13</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>419.5 7</intersection>
<intersection>452 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>419.5,9,419.5,13</points>
<connection>
<GID>359</GID>
<name>N_in1</name></connection>
<intersection>13 4</intersection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>445,27,449.5,27</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>449.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449.5,11,449.5,27</points>
<intersection>11 5</intersection>
<intersection>22.5 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>449.5,11,453,11</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>449.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>449.5,22.5,453,22.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>449.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>459,21.5,462,21.5</points>
<connection>
<GID>348</GID>
<name>N_in0</name></connection>
<connection>
<GID>345</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>425,31,434,31</points>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection>
<intersection>434 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>434,8.5,434,31</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>28 6</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>434,28,439,28</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>434 4</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>425,26,439,26</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>429 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>429,6.5,429,26</points>
<intersection>6.5 4</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>429,6.5,434,6.5</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>429 3</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440,7.5,463,7.5</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<connection>
<GID>347</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,9.5,516,12</points>
<intersection>9.5 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,9.5,518,9.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,12,516,12</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<intersection>516 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>507,20.5,508,20.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>507 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>507,13,507,20.5</points>
<intersection>13 4</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>480.5,13,508,13</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>480.5 7</intersection>
<intersection>507 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>480.5,8.5,480.5,13</points>
<connection>
<GID>317</GID>
<name>N_in1</name></connection>
<intersection>13 4</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>500,27,504.5,27</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<intersection>504.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>504.5,11,504.5,27</points>
<intersection>11 5</intersection>
<intersection>22.5 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>504.5,11,508,11</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<intersection>504.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>504.5,22.5,508,22.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>504.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>514,21.5,517,21.5</points>
<connection>
<GID>241</GID>
<name>N_in0</name></connection>
<connection>
<GID>237</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>480,31,489,31</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>489 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>489,8.5,489,31</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>28 6</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>489,28,494,28</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>489 4</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>480,26,494,26</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>484.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>484.5,6.5,484.5,26</points>
<intersection>6.5 4</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>484.5,6.5,489,6.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>484.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>495,7.5,518,7.5</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<connection>
<GID>240</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>469,8.5,478.5,8.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<connection>
<GID>317</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>299.5,9,309,9</points>
<connection>
<GID>357</GID>
<name>N_in0</name></connection>
<connection>
<GID>215</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410,9,417.5,9</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<connection>
<GID>359</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524,8.5,532,8.5</points>
<connection>
<GID>361</GID>
<name>N_in0</name></connection>
<connection>
<GID>240</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,10,347,12.5</points>
<intersection>10 1</intersection>
<intersection>12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,10,349,10</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>347 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>345,12.5,347,12.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>347 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>338,21,339,21</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>338 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>338,13.5,338,21</points>
<intersection>13.5 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>311,13.5,339,13.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>311 10</intersection>
<intersection>338 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>311,9,311,13.5</points>
<connection>
<GID>357</GID>
<name>N_in1</name></connection>
<intersection>13.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>331,27.5,335.5,27.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>335.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335.5,11.5,335.5,27.5</points>
<intersection>11.5 5</intersection>
<intersection>23 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>335.5,11.5,339,11.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>335.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>335.5,23,339,23</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>335.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>345,22,348,22</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>310.5,31.5,320,31.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>320 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>320,9,320,31.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>28.5 6</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>320,28.5,325,28.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>320 4</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>311,26.5,325,26.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>315.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>315.5,7,315.5,26.5</points>
<intersection>7 4</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>315.5,7,320,7</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>315.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>326,8,349,8</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402,10,402,12.5</points>
<intersection>10 1</intersection>
<intersection>12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,10,404,10</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400,12.5,402,12.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>402 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>393,21,394,21</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>393 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>393,13.5,393,21</points>
<intersection>13.5 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>366.5,13.5,394,13.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>366.5 7</intersection>
<intersection>393 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>366.5,9,366.5,13.5</points>
<connection>
<GID>142</GID>
<name>N_in1</name></connection>
<intersection>13.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>386,27.5,390.5,27.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>390.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>390.5,11.5,390.5,27.5</points>
<intersection>11.5 5</intersection>
<intersection>23 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>390.5,11.5,394,11.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>390.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>390.5,23,394,23</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>390.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>400,22,403,22</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366,31.5,375,31.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>375 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375,9,375,31.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>28.5 6</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>375,28.5,380,28.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>375 4</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>366,26.5,380,26.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>370.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>370.5,7,370.5,26.5</points>
<intersection>7 4</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>370.5,7,375,7</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>370.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381,8,404,8</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 3>
<page 4>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 4>
<page 5>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 5>
<page 6>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 6>
<page 7>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 7>
<page 8>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 8>
<page 9>
<PageViewport>-3.20813e-005,126.574,938.642,-337.379</PageViewport></page 9></circuit>