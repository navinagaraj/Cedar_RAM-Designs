<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-432.832,512.756,791.168,-92.2437</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-60.5,-975.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>BE_DECODER_3x8</type>
<position>-266.5,-1337</position>
<output>
<ID>OUT_0</ID>1555 </output>
<output>
<ID>OUT_1</ID>1554 </output>
<output>
<ID>OUT_2</ID>1553 </output>
<output>
<ID>OUT_3</ID>5 </output>
<output>
<ID>OUT_4</ID>4 </output>
<output>
<ID>OUT_5</ID>3 </output>
<output>
<ID>OUT_6</ID>2 </output>
<output>
<ID>OUT_7</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1552</ID>
<type>AE_DFF_LOW</type>
<position>-26.5,-122</position>
<output>
<ID>OUT_0</ID>888 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1553</ID>
<type>AA_AND2</type>
<position>-16.5,-127.5</position>
<input>
<ID>IN_0</ID>888 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1554</ID>
<type>AE_DFF_LOW</type>
<position>23,-122</position>
<output>
<ID>OUT_0</ID>889 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1555</ID>
<type>AA_AND2</type>
<position>32,-128.5</position>
<input>
<ID>IN_0</ID>889 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1556</ID>
<type>AE_DFF_LOW</type>
<position>71,-122</position>
<output>
<ID>OUT_0</ID>891 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1557</ID>
<type>AA_AND2</type>
<position>78.5,-127.5</position>
<input>
<ID>IN_0</ID>891 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1558</ID>
<type>AE_DFF_LOW</type>
<position>120.5,-122</position>
<output>
<ID>OUT_0</ID>892 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1559</ID>
<type>AA_AND2</type>
<position>129,-127.5</position>
<input>
<ID>IN_0</ID>892 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1560</ID>
<type>AE_DFF_LOW</type>
<position>168.5,-122</position>
<output>
<ID>OUT_0</ID>893 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1561</ID>
<type>AA_AND2</type>
<position>177,-127</position>
<input>
<ID>IN_0</ID>893 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1562</ID>
<type>AE_DFF_LOW</type>
<position>226,-122</position>
<output>
<ID>OUT_0</ID>894 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1563</ID>
<type>AA_AND2</type>
<position>235.5,-129</position>
<input>
<ID>IN_0</ID>894 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1564</ID>
<type>AE_DFF_LOW</type>
<position>281,-122</position>
<output>
<ID>OUT_0</ID>895 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1565</ID>
<type>AA_AND2</type>
<position>289,-128</position>
<input>
<ID>IN_0</ID>895 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1566</ID>
<type>AE_DFF_LOW</type>
<position>338,-122</position>
<output>
<ID>OUT_0</ID>896 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1567</ID>
<type>AA_AND2</type>
<position>347.5,-128.5</position>
<input>
<ID>IN_0</ID>896 </input>
<input>
<ID>IN_1</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1568</ID>
<type>AA_AND2</type>
<position>-58,-121</position>
<input>
<ID>IN_0</ID>897 </input>
<output>
<ID>OUT</ID>890 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1569</ID>
<type>AE_DFF_LOW</type>
<position>-26.5,-136</position>
<output>
<ID>OUT_0</ID>898 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1570</ID>
<type>AA_AND2</type>
<position>-16.5,-141.5</position>
<input>
<ID>IN_0</ID>898 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1571</ID>
<type>AE_DFF_LOW</type>
<position>23,-136</position>
<output>
<ID>OUT_0</ID>899 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1572</ID>
<type>AA_AND2</type>
<position>32,-142.5</position>
<input>
<ID>IN_0</ID>899 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1573</ID>
<type>AE_DFF_LOW</type>
<position>71,-136</position>
<output>
<ID>OUT_0</ID>901 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1574</ID>
<type>AA_AND2</type>
<position>78.5,-141.5</position>
<input>
<ID>IN_0</ID>901 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1575</ID>
<type>AE_DFF_LOW</type>
<position>120.5,-136</position>
<output>
<ID>OUT_0</ID>902 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1576</ID>
<type>AA_AND2</type>
<position>129,-141.5</position>
<input>
<ID>IN_0</ID>902 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1577</ID>
<type>AE_DFF_LOW</type>
<position>168.5,-136</position>
<output>
<ID>OUT_0</ID>903 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1578</ID>
<type>AA_AND2</type>
<position>177,-141</position>
<input>
<ID>IN_0</ID>903 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1579</ID>
<type>AE_DFF_LOW</type>
<position>226,-136</position>
<output>
<ID>OUT_0</ID>904 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1580</ID>
<type>AA_AND2</type>
<position>235.5,-143</position>
<input>
<ID>IN_0</ID>904 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1581</ID>
<type>AE_DFF_LOW</type>
<position>281,-136</position>
<output>
<ID>OUT_0</ID>905 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1582</ID>
<type>AA_AND2</type>
<position>289,-142</position>
<input>
<ID>IN_0</ID>905 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1583</ID>
<type>AE_DFF_LOW</type>
<position>338,-136</position>
<output>
<ID>OUT_0</ID>906 </output>
<input>
<ID>clock</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1584</ID>
<type>AA_AND2</type>
<position>347.5,-142.5</position>
<input>
<ID>IN_0</ID>906 </input>
<input>
<ID>IN_1</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1585</ID>
<type>AA_AND2</type>
<position>-58,-135</position>
<input>
<ID>IN_0</ID>907 </input>
<output>
<ID>OUT</ID>900 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1586</ID>
<type>AE_DFF_LOW</type>
<position>-27,-153.5</position>
<output>
<ID>OUT_0</ID>908 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1587</ID>
<type>AA_AND2</type>
<position>-17,-159</position>
<input>
<ID>IN_0</ID>908 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1588</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-153.5</position>
<output>
<ID>OUT_0</ID>909 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1589</ID>
<type>AA_AND2</type>
<position>31.5,-160</position>
<input>
<ID>IN_0</ID>909 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1590</ID>
<type>AE_DFF_LOW</type>
<position>70.5,-153.5</position>
<output>
<ID>OUT_0</ID>911 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1591</ID>
<type>AA_AND2</type>
<position>78,-159</position>
<input>
<ID>IN_0</ID>911 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1592</ID>
<type>AE_DFF_LOW</type>
<position>120,-153.5</position>
<output>
<ID>OUT_0</ID>912 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1593</ID>
<type>AA_AND2</type>
<position>128.5,-159</position>
<input>
<ID>IN_0</ID>912 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1594</ID>
<type>AE_DFF_LOW</type>
<position>168,-153.5</position>
<output>
<ID>OUT_0</ID>913 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1595</ID>
<type>AA_AND2</type>
<position>176.5,-158.5</position>
<input>
<ID>IN_0</ID>913 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1596</ID>
<type>AE_DFF_LOW</type>
<position>225.5,-153.5</position>
<output>
<ID>OUT_0</ID>914 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1597</ID>
<type>AA_AND2</type>
<position>235,-160.5</position>
<input>
<ID>IN_0</ID>914 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1598</ID>
<type>AE_DFF_LOW</type>
<position>280.5,-153.5</position>
<output>
<ID>OUT_0</ID>915 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1599</ID>
<type>AA_AND2</type>
<position>288.5,-159.5</position>
<input>
<ID>IN_0</ID>915 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1600</ID>
<type>AE_DFF_LOW</type>
<position>337.5,-153.5</position>
<output>
<ID>OUT_0</ID>916 </output>
<input>
<ID>clock</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>57</ID>
<type>BE_DECODER_3x8</type>
<position>-85,-88</position>
<input>
<ID>ENABLE</ID>1 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>917 </output>
<output>
<ID>OUT_1</ID>907 </output>
<output>
<ID>OUT_2</ID>897 </output>
<output>
<ID>OUT_3</ID>878 </output>
<output>
<ID>OUT_4</ID>868 </output>
<output>
<ID>OUT_5</ID>858 </output>
<output>
<ID>OUT_6</ID>848 </output>
<output>
<ID>OUT_7</ID>838 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1601</ID>
<type>AA_AND2</type>
<position>347,-160</position>
<input>
<ID>IN_0</ID>916 </input>
<input>
<ID>IN_1</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1602</ID>
<type>AA_AND2</type>
<position>-58.5,-152.5</position>
<input>
<ID>IN_0</ID>917 </input>
<output>
<ID>OUT</ID>910 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1603</ID>
<type>AE_DFF_LOW</type>
<position>-1.5,-355</position>
<output>
<ID>OUT_0</ID>963 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1604</ID>
<type>AA_AND2</type>
<position>8.5,-360.5</position>
<input>
<ID>IN_0</ID>963 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1605</ID>
<type>AE_DFF_LOW</type>
<position>48,-355</position>
<output>
<ID>OUT_0</ID>964 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1606</ID>
<type>AA_AND2</type>
<position>57,-361.5</position>
<input>
<ID>IN_0</ID>964 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1607</ID>
<type>AE_DFF_LOW</type>
<position>96,-355</position>
<output>
<ID>OUT_0</ID>966 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1608</ID>
<type>AA_AND2</type>
<position>103.5,-360.5</position>
<input>
<ID>IN_0</ID>966 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1609</ID>
<type>AE_DFF_LOW</type>
<position>145.5,-355</position>
<output>
<ID>OUT_0</ID>967 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1610</ID>
<type>AA_AND2</type>
<position>154,-360.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1611</ID>
<type>AE_DFF_LOW</type>
<position>193.5,-355</position>
<output>
<ID>OUT_0</ID>968 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1612</ID>
<type>AA_AND2</type>
<position>202,-360</position>
<input>
<ID>IN_0</ID>968 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1613</ID>
<type>AE_DFF_LOW</type>
<position>251,-355</position>
<output>
<ID>OUT_0</ID>969 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1614</ID>
<type>AA_AND2</type>
<position>260.5,-362</position>
<input>
<ID>IN_0</ID>969 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1615</ID>
<type>AE_DFF_LOW</type>
<position>306,-355</position>
<output>
<ID>OUT_0</ID>970 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1616</ID>
<type>AA_AND2</type>
<position>314,-361</position>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1617</ID>
<type>AE_DFF_LOW</type>
<position>363,-355</position>
<output>
<ID>OUT_0</ID>971 </output>
<input>
<ID>clock</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1618</ID>
<type>AA_AND2</type>
<position>372.5,-361.5</position>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1619</ID>
<type>AA_AND2</type>
<position>-33,-354</position>
<input>
<ID>IN_0</ID>995 </input>
<output>
<ID>OUT</ID>965 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1620</ID>
<type>AE_DFF_LOW</type>
<position>-1.5,-369</position>
<output>
<ID>OUT_0</ID>972 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1621</ID>
<type>AA_AND2</type>
<position>8.5,-374.5</position>
<input>
<ID>IN_0</ID>972 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1622</ID>
<type>AE_DFF_LOW</type>
<position>48,-369</position>
<output>
<ID>OUT_0</ID>973 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1623</ID>
<type>AA_AND2</type>
<position>57,-375.5</position>
<input>
<ID>IN_0</ID>973 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1624</ID>
<type>AE_DFF_LOW</type>
<position>96,-369</position>
<output>
<ID>OUT_0</ID>975 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1625</ID>
<type>AA_AND2</type>
<position>103.5,-374.5</position>
<input>
<ID>IN_0</ID>975 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1626</ID>
<type>AE_DFF_LOW</type>
<position>145.5,-369</position>
<output>
<ID>OUT_0</ID>976 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1627</ID>
<type>AA_AND2</type>
<position>154,-374.5</position>
<input>
<ID>IN_0</ID>976 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1628</ID>
<type>AE_DFF_LOW</type>
<position>193.5,-369</position>
<output>
<ID>OUT_0</ID>977 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1629</ID>
<type>AA_AND2</type>
<position>202,-374</position>
<input>
<ID>IN_0</ID>977 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1630</ID>
<type>AE_DFF_LOW</type>
<position>251,-369</position>
<output>
<ID>OUT_0</ID>978 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1631</ID>
<type>AA_AND2</type>
<position>260.5,-376</position>
<input>
<ID>IN_0</ID>978 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1632</ID>
<type>AE_DFF_LOW</type>
<position>306,-369</position>
<output>
<ID>OUT_0</ID>979 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1633</ID>
<type>AA_AND2</type>
<position>314,-375</position>
<input>
<ID>IN_0</ID>979 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1634</ID>
<type>AE_DFF_LOW</type>
<position>363,-369</position>
<output>
<ID>OUT_0</ID>980 </output>
<input>
<ID>clock</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1635</ID>
<type>AA_AND2</type>
<position>372.5,-375.5</position>
<input>
<ID>IN_0</ID>980 </input>
<input>
<ID>IN_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1636</ID>
<type>AA_AND2</type>
<position>-33,-368</position>
<input>
<ID>IN_0</ID>996 </input>
<output>
<ID>OUT</ID>974 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1637</ID>
<type>AE_DFF_LOW</type>
<position>-2,-386.5</position>
<output>
<ID>OUT_0</ID>981 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1638</ID>
<type>AA_AND2</type>
<position>8,-392</position>
<input>
<ID>IN_0</ID>981 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1639</ID>
<type>AE_DFF_LOW</type>
<position>47.5,-386.5</position>
<output>
<ID>OUT_0</ID>982 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1640</ID>
<type>AA_AND2</type>
<position>56.5,-393</position>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1641</ID>
<type>AE_DFF_LOW</type>
<position>95.5,-386.5</position>
<output>
<ID>OUT_0</ID>984 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1642</ID>
<type>AA_AND2</type>
<position>103,-392</position>
<input>
<ID>IN_0</ID>984 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1643</ID>
<type>AE_DFF_LOW</type>
<position>145,-386.5</position>
<output>
<ID>OUT_0</ID>985 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1644</ID>
<type>AA_AND2</type>
<position>153.5,-392</position>
<input>
<ID>IN_0</ID>985 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1645</ID>
<type>AE_DFF_LOW</type>
<position>193,-386.5</position>
<output>
<ID>OUT_0</ID>986 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1646</ID>
<type>AA_AND2</type>
<position>201.5,-391.5</position>
<input>
<ID>IN_0</ID>986 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1647</ID>
<type>AE_DFF_LOW</type>
<position>250.5,-386.5</position>
<output>
<ID>OUT_0</ID>987 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1648</ID>
<type>AA_AND2</type>
<position>260,-393.5</position>
<input>
<ID>IN_0</ID>987 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1649</ID>
<type>AE_DFF_LOW</type>
<position>305.5,-386.5</position>
<output>
<ID>OUT_0</ID>988 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1650</ID>
<type>AA_AND2</type>
<position>313.5,-392.5</position>
<input>
<ID>IN_0</ID>988 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1651</ID>
<type>AE_DFF_LOW</type>
<position>362.5,-386.5</position>
<output>
<ID>OUT_0</ID>989 </output>
<input>
<ID>clock</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1652</ID>
<type>AA_AND2</type>
<position>372,-393</position>
<input>
<ID>IN_0</ID>989 </input>
<input>
<ID>IN_1</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1653</ID>
<type>AA_AND2</type>
<position>-33.5,-385.5</position>
<input>
<ID>IN_0</ID>997 </input>
<output>
<ID>OUT</ID>983 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1654</ID>
<type>AE_DFF_LOW</type>
<position>-0.5,-287</position>
<output>
<ID>OUT_0</ID>918 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1655</ID>
<type>AA_AND2</type>
<position>9.5,-292.5</position>
<input>
<ID>IN_0</ID>918 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1656</ID>
<type>AE_DFF_LOW</type>
<position>49,-287</position>
<output>
<ID>OUT_0</ID>919 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1657</ID>
<type>AA_AND2</type>
<position>58,-293.5</position>
<input>
<ID>IN_0</ID>919 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1658</ID>
<type>AE_DFF_LOW</type>
<position>97,-287</position>
<output>
<ID>OUT_0</ID>921 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1659</ID>
<type>AA_AND2</type>
<position>104.5,-292.5</position>
<input>
<ID>IN_0</ID>921 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1660</ID>
<type>AE_DFF_LOW</type>
<position>146.5,-287</position>
<output>
<ID>OUT_0</ID>922 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1661</ID>
<type>AA_AND2</type>
<position>155,-292.5</position>
<input>
<ID>IN_0</ID>922 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1662</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-287</position>
<output>
<ID>OUT_0</ID>923 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1663</ID>
<type>AA_AND2</type>
<position>203,-292</position>
<input>
<ID>IN_0</ID>923 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1664</ID>
<type>AE_DFF_LOW</type>
<position>252,-287</position>
<output>
<ID>OUT_0</ID>924 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1665</ID>
<type>AA_AND2</type>
<position>261.5,-294</position>
<input>
<ID>IN_0</ID>924 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1666</ID>
<type>AE_DFF_LOW</type>
<position>307,-287</position>
<output>
<ID>OUT_0</ID>925 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1667</ID>
<type>AA_AND2</type>
<position>315,-293</position>
<input>
<ID>IN_0</ID>925 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1668</ID>
<type>AE_DFF_LOW</type>
<position>364,-287</position>
<output>
<ID>OUT_0</ID>926 </output>
<input>
<ID>clock</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1669</ID>
<type>AA_AND2</type>
<position>373.5,-293.5</position>
<input>
<ID>IN_0</ID>926 </input>
<input>
<ID>IN_1</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1670</ID>
<type>AA_AND2</type>
<position>-32,-286</position>
<input>
<ID>IN_0</ID>990 </input>
<output>
<ID>OUT</ID>920 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1671</ID>
<type>AE_DFF_LOW</type>
<position>-0.5,-300</position>
<output>
<ID>OUT_0</ID>927 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1672</ID>
<type>AA_AND2</type>
<position>9.5,-305.5</position>
<input>
<ID>IN_0</ID>927 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1673</ID>
<type>AE_DFF_LOW</type>
<position>49,-300</position>
<output>
<ID>OUT_0</ID>928 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1674</ID>
<type>AA_AND2</type>
<position>58,-306.5</position>
<input>
<ID>IN_0</ID>928 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1675</ID>
<type>AE_DFF_LOW</type>
<position>97,-300</position>
<output>
<ID>OUT_0</ID>930 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1676</ID>
<type>AA_AND2</type>
<position>104.5,-305.5</position>
<input>
<ID>IN_0</ID>930 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1677</ID>
<type>AE_DFF_LOW</type>
<position>146.5,-300</position>
<output>
<ID>OUT_0</ID>931 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1678</ID>
<type>AA_AND2</type>
<position>155,-305.5</position>
<input>
<ID>IN_0</ID>931 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1679</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-300</position>
<output>
<ID>OUT_0</ID>932 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1680</ID>
<type>AA_AND2</type>
<position>203,-305</position>
<input>
<ID>IN_0</ID>932 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1681</ID>
<type>AE_DFF_LOW</type>
<position>252,-300</position>
<output>
<ID>OUT_0</ID>933 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1682</ID>
<type>AA_AND2</type>
<position>261.5,-307</position>
<input>
<ID>IN_0</ID>933 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1683</ID>
<type>AE_DFF_LOW</type>
<position>307,-300</position>
<output>
<ID>OUT_0</ID>934 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1684</ID>
<type>AA_AND2</type>
<position>315,-306</position>
<input>
<ID>IN_0</ID>934 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1685</ID>
<type>AE_DFF_LOW</type>
<position>364,-300</position>
<output>
<ID>OUT_0</ID>935 </output>
<input>
<ID>clock</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1686</ID>
<type>AA_AND2</type>
<position>373.5,-306.5</position>
<input>
<ID>IN_0</ID>935 </input>
<input>
<ID>IN_1</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1687</ID>
<type>AA_AND2</type>
<position>-32,-299</position>
<input>
<ID>IN_0</ID>991 </input>
<output>
<ID>OUT</ID>929 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1688</ID>
<type>AE_DFF_LOW</type>
<position>-0.5,-314.5</position>
<output>
<ID>OUT_0</ID>936 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1689</ID>
<type>AA_AND2</type>
<position>9.5,-320</position>
<input>
<ID>IN_0</ID>936 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1690</ID>
<type>AE_DFF_LOW</type>
<position>49,-314.5</position>
<output>
<ID>OUT_0</ID>937 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1691</ID>
<type>AA_AND2</type>
<position>58,-321</position>
<input>
<ID>IN_0</ID>937 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1692</ID>
<type>AE_DFF_LOW</type>
<position>97,-314.5</position>
<output>
<ID>OUT_0</ID>939 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1693</ID>
<type>AA_AND2</type>
<position>104.5,-320</position>
<input>
<ID>IN_0</ID>939 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1694</ID>
<type>AE_DFF_LOW</type>
<position>146.5,-314.5</position>
<output>
<ID>OUT_0</ID>940 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1695</ID>
<type>AA_AND2</type>
<position>155,-320</position>
<input>
<ID>IN_0</ID>940 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1696</ID>
<type>AE_DFF_LOW</type>
<position>194.5,-314.5</position>
<output>
<ID>OUT_0</ID>941 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1697</ID>
<type>AA_AND2</type>
<position>203,-319.5</position>
<input>
<ID>IN_0</ID>941 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1698</ID>
<type>AE_DFF_LOW</type>
<position>252,-314.5</position>
<output>
<ID>OUT_0</ID>942 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1699</ID>
<type>AA_AND2</type>
<position>261.5,-321.5</position>
<input>
<ID>IN_0</ID>942 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1700</ID>
<type>AE_DFF_LOW</type>
<position>307,-314.5</position>
<output>
<ID>OUT_0</ID>943 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1701</ID>
<type>AA_AND2</type>
<position>315,-320.5</position>
<input>
<ID>IN_0</ID>943 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1702</ID>
<type>AE_DFF_LOW</type>
<position>364,-314.5</position>
<output>
<ID>OUT_0</ID>944 </output>
<input>
<ID>clock</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1703</ID>
<type>AA_AND2</type>
<position>373.5,-321</position>
<input>
<ID>IN_0</ID>944 </input>
<input>
<ID>IN_1</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1704</ID>
<type>AA_AND2</type>
<position>-32,-313.5</position>
<input>
<ID>IN_0</ID>992 </input>
<output>
<ID>OUT</ID>938 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1705</ID>
<type>AE_DFF_LOW</type>
<position>-1,-327</position>
<output>
<ID>OUT_0</ID>945 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1706</ID>
<type>AA_AND2</type>
<position>9,-332.5</position>
<input>
<ID>IN_0</ID>945 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1707</ID>
<type>AE_DFF_LOW</type>
<position>48.5,-327</position>
<output>
<ID>OUT_0</ID>946 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1708</ID>
<type>AA_AND2</type>
<position>57.5,-333.5</position>
<input>
<ID>IN_0</ID>946 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1709</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-327</position>
<output>
<ID>OUT_0</ID>948 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1710</ID>
<type>AA_AND2</type>
<position>104,-332.5</position>
<input>
<ID>IN_0</ID>948 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1711</ID>
<type>AE_DFF_LOW</type>
<position>146,-327</position>
<output>
<ID>OUT_0</ID>949 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1712</ID>
<type>AA_AND2</type>
<position>154.5,-332.5</position>
<input>
<ID>IN_0</ID>949 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1713</ID>
<type>AE_DFF_LOW</type>
<position>194,-327</position>
<output>
<ID>OUT_0</ID>950 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1714</ID>
<type>AA_AND2</type>
<position>202.5,-332</position>
<input>
<ID>IN_0</ID>950 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1715</ID>
<type>AE_DFF_LOW</type>
<position>251.5,-327</position>
<output>
<ID>OUT_0</ID>951 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1716</ID>
<type>AA_AND2</type>
<position>261,-334</position>
<input>
<ID>IN_0</ID>951 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1717</ID>
<type>AE_DFF_LOW</type>
<position>306.5,-327</position>
<output>
<ID>OUT_0</ID>952 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1718</ID>
<type>AA_AND2</type>
<position>314.5,-333</position>
<input>
<ID>IN_0</ID>952 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1719</ID>
<type>AE_DFF_LOW</type>
<position>363.5,-327</position>
<output>
<ID>OUT_0</ID>953 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1720</ID>
<type>AA_AND2</type>
<position>373,-333.5</position>
<input>
<ID>IN_0</ID>953 </input>
<input>
<ID>IN_1</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1721</ID>
<type>AA_AND2</type>
<position>-32.5,-326</position>
<input>
<ID>IN_0</ID>993 </input>
<output>
<ID>OUT</ID>947 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1722</ID>
<type>AE_DFF_LOW</type>
<position>-1.5,-340</position>
<output>
<ID>OUT_0</ID>954 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1723</ID>
<type>AA_AND2</type>
<position>8.5,-345.5</position>
<input>
<ID>IN_0</ID>954 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1724</ID>
<type>AE_DFF_LOW</type>
<position>48,-340</position>
<output>
<ID>OUT_0</ID>955 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1725</ID>
<type>AA_AND2</type>
<position>57,-346.5</position>
<input>
<ID>IN_0</ID>955 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1726</ID>
<type>AE_DFF_LOW</type>
<position>96,-340</position>
<output>
<ID>OUT_0</ID>957 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1727</ID>
<type>AA_AND2</type>
<position>103.5,-345.5</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1728</ID>
<type>AE_DFF_LOW</type>
<position>145.5,-340</position>
<output>
<ID>OUT_0</ID>958 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1729</ID>
<type>AA_AND2</type>
<position>154,-345.5</position>
<input>
<ID>IN_0</ID>958 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1730</ID>
<type>AE_DFF_LOW</type>
<position>193.5,-340</position>
<output>
<ID>OUT_0</ID>959 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1731</ID>
<type>AA_AND2</type>
<position>202,-345</position>
<input>
<ID>IN_0</ID>959 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1732</ID>
<type>AE_DFF_LOW</type>
<position>251,-340</position>
<output>
<ID>OUT_0</ID>960 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1733</ID>
<type>AA_AND2</type>
<position>260.5,-347</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1734</ID>
<type>AE_DFF_LOW</type>
<position>306,-340</position>
<output>
<ID>OUT_0</ID>961 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1735</ID>
<type>AA_AND2</type>
<position>314,-346</position>
<input>
<ID>IN_0</ID>961 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1736</ID>
<type>AE_DFF_LOW</type>
<position>363,-340</position>
<output>
<ID>OUT_0</ID>962 </output>
<input>
<ID>clock</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1737</ID>
<type>AA_AND2</type>
<position>372.5,-346.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1738</ID>
<type>AA_AND2</type>
<position>-33,-339</position>
<input>
<ID>IN_0</ID>994 </input>
<output>
<ID>OUT</ID>956 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>BE_DECODER_3x8</type>
<position>-81.5,-326.5</position>
<input>
<ID>ENABLE</ID>2 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>997 </output>
<output>
<ID>OUT_1</ID>996 </output>
<output>
<ID>OUT_2</ID>995 </output>
<output>
<ID>OUT_3</ID>994 </output>
<output>
<ID>OUT_4</ID>993 </output>
<output>
<ID>OUT_5</ID>992 </output>
<output>
<ID>OUT_6</ID>991 </output>
<output>
<ID>OUT_7</ID>990 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1739</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-641.5</position>
<output>
<ID>OUT_0</ID>1043 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1740</ID>
<type>AA_AND2</type>
<position>-8.5,-647</position>
<input>
<ID>IN_0</ID>1043 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1741</ID>
<type>AE_DFF_LOW</type>
<position>31,-641.5</position>
<output>
<ID>OUT_0</ID>1044 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1742</ID>
<type>AA_AND2</type>
<position>40,-648</position>
<input>
<ID>IN_0</ID>1044 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1743</ID>
<type>AE_DFF_LOW</type>
<position>79,-641.5</position>
<output>
<ID>OUT_0</ID>1046 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1744</ID>
<type>AA_AND2</type>
<position>86.5,-647</position>
<input>
<ID>IN_0</ID>1046 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1745</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-641.5</position>
<output>
<ID>OUT_0</ID>1047 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1746</ID>
<type>AA_AND2</type>
<position>137,-647</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1747</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-641.5</position>
<output>
<ID>OUT_0</ID>1048 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1748</ID>
<type>AA_AND2</type>
<position>185,-646.5</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1749</ID>
<type>AE_DFF_LOW</type>
<position>234,-641.5</position>
<output>
<ID>OUT_0</ID>1049 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1750</ID>
<type>AA_AND2</type>
<position>243.5,-648.5</position>
<input>
<ID>IN_0</ID>1049 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1751</ID>
<type>AE_DFF_LOW</type>
<position>289,-641.5</position>
<output>
<ID>OUT_0</ID>1050 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1752</ID>
<type>AA_AND2</type>
<position>297,-647.5</position>
<input>
<ID>IN_0</ID>1050 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1753</ID>
<type>AE_DFF_LOW</type>
<position>346,-641.5</position>
<output>
<ID>OUT_0</ID>1051 </output>
<input>
<ID>clock</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1754</ID>
<type>AA_AND2</type>
<position>355.5,-648</position>
<input>
<ID>IN_0</ID>1051 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1755</ID>
<type>AA_AND2</type>
<position>-50,-640.5</position>
<input>
<ID>IN_0</ID>1075 </input>
<output>
<ID>OUT</ID>1045 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1756</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-655.5</position>
<output>
<ID>OUT_0</ID>1052 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1757</ID>
<type>AA_AND2</type>
<position>-8.5,-661</position>
<input>
<ID>IN_0</ID>1052 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1758</ID>
<type>AE_DFF_LOW</type>
<position>31,-655.5</position>
<output>
<ID>OUT_0</ID>1053 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1759</ID>
<type>AA_AND2</type>
<position>40,-662</position>
<input>
<ID>IN_0</ID>1053 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1760</ID>
<type>AE_DFF_LOW</type>
<position>79,-655.5</position>
<output>
<ID>OUT_0</ID>1055 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1761</ID>
<type>AA_AND2</type>
<position>86.5,-661</position>
<input>
<ID>IN_0</ID>1055 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1762</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-655.5</position>
<output>
<ID>OUT_0</ID>1056 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1763</ID>
<type>AA_AND2</type>
<position>137,-661</position>
<input>
<ID>IN_0</ID>1056 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1764</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-655.5</position>
<output>
<ID>OUT_0</ID>1057 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1765</ID>
<type>AA_AND2</type>
<position>185,-660.5</position>
<input>
<ID>IN_0</ID>1057 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1766</ID>
<type>AE_DFF_LOW</type>
<position>234,-655.5</position>
<output>
<ID>OUT_0</ID>1058 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1767</ID>
<type>AA_AND2</type>
<position>243.5,-662.5</position>
<input>
<ID>IN_0</ID>1058 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1768</ID>
<type>AE_DFF_LOW</type>
<position>289,-655.5</position>
<output>
<ID>OUT_0</ID>1059 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1769</ID>
<type>AA_AND2</type>
<position>297,-661.5</position>
<input>
<ID>IN_0</ID>1059 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1770</ID>
<type>AE_DFF_LOW</type>
<position>346,-655.5</position>
<output>
<ID>OUT_0</ID>1060 </output>
<input>
<ID>clock</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1771</ID>
<type>AA_AND2</type>
<position>355.5,-662</position>
<input>
<ID>IN_0</ID>1060 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1772</ID>
<type>AA_AND2</type>
<position>-50,-654.5</position>
<input>
<ID>IN_0</ID>1076 </input>
<output>
<ID>OUT</ID>1054 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1773</ID>
<type>AE_DFF_LOW</type>
<position>-19,-673</position>
<output>
<ID>OUT_0</ID>1061 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1774</ID>
<type>AA_AND2</type>
<position>-9,-678.5</position>
<input>
<ID>IN_0</ID>1061 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1775</ID>
<type>AE_DFF_LOW</type>
<position>30.5,-673</position>
<output>
<ID>OUT_0</ID>1062 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1776</ID>
<type>AA_AND2</type>
<position>39.5,-679.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1777</ID>
<type>AE_DFF_LOW</type>
<position>78.5,-673</position>
<output>
<ID>OUT_0</ID>1064 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1778</ID>
<type>AA_AND2</type>
<position>86,-678.5</position>
<input>
<ID>IN_0</ID>1064 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1779</ID>
<type>AE_DFF_LOW</type>
<position>128,-673</position>
<output>
<ID>OUT_0</ID>1065 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1780</ID>
<type>AA_AND2</type>
<position>136.5,-678.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1781</ID>
<type>AE_DFF_LOW</type>
<position>176,-673</position>
<output>
<ID>OUT_0</ID>1066 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1782</ID>
<type>AA_AND2</type>
<position>184.5,-678</position>
<input>
<ID>IN_0</ID>1066 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1783</ID>
<type>AE_DFF_LOW</type>
<position>233.5,-673</position>
<output>
<ID>OUT_0</ID>1067 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1784</ID>
<type>AA_AND2</type>
<position>243,-680</position>
<input>
<ID>IN_0</ID>1067 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1785</ID>
<type>AE_DFF_LOW</type>
<position>288.5,-673</position>
<output>
<ID>OUT_0</ID>1068 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1786</ID>
<type>AA_AND2</type>
<position>296.5,-679</position>
<input>
<ID>IN_0</ID>1068 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1787</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-673</position>
<output>
<ID>OUT_0</ID>1069 </output>
<input>
<ID>clock</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1788</ID>
<type>AA_AND2</type>
<position>355,-679.5</position>
<input>
<ID>IN_0</ID>1069 </input>
<input>
<ID>IN_1</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1789</ID>
<type>AA_AND2</type>
<position>-50.5,-672</position>
<input>
<ID>IN_0</ID>1077 </input>
<output>
<ID>OUT</ID>1063 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1790</ID>
<type>AE_DFF_LOW</type>
<position>-17.5,-573.5</position>
<output>
<ID>OUT_0</ID>998 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1791</ID>
<type>AA_AND2</type>
<position>-7.5,-579</position>
<input>
<ID>IN_0</ID>998 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1792</ID>
<type>AE_DFF_LOW</type>
<position>32,-573.5</position>
<output>
<ID>OUT_0</ID>999 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1793</ID>
<type>AA_AND2</type>
<position>41,-580</position>
<input>
<ID>IN_0</ID>999 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1794</ID>
<type>AE_DFF_LOW</type>
<position>80,-573.5</position>
<output>
<ID>OUT_0</ID>1001 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1795</ID>
<type>AA_AND2</type>
<position>87.5,-579</position>
<input>
<ID>IN_0</ID>1001 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1796</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-573.5</position>
<output>
<ID>OUT_0</ID>1002 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1797</ID>
<type>AA_AND2</type>
<position>138,-579</position>
<input>
<ID>IN_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1798</ID>
<type>AE_DFF_LOW</type>
<position>177.5,-573.5</position>
<output>
<ID>OUT_0</ID>1003 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1799</ID>
<type>AA_AND2</type>
<position>186,-578.5</position>
<input>
<ID>IN_0</ID>1003 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1800</ID>
<type>AE_DFF_LOW</type>
<position>235,-573.5</position>
<output>
<ID>OUT_0</ID>1004 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1801</ID>
<type>AA_AND2</type>
<position>244.5,-580.5</position>
<input>
<ID>IN_0</ID>1004 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1802</ID>
<type>AE_DFF_LOW</type>
<position>290,-573.5</position>
<output>
<ID>OUT_0</ID>1005 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1803</ID>
<type>AA_AND2</type>
<position>298,-579.5</position>
<input>
<ID>IN_0</ID>1005 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1804</ID>
<type>AE_DFF_LOW</type>
<position>347,-573.5</position>
<output>
<ID>OUT_0</ID>1006 </output>
<input>
<ID>clock</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1805</ID>
<type>AA_AND2</type>
<position>356.5,-580</position>
<input>
<ID>IN_0</ID>1006 </input>
<input>
<ID>IN_1</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1806</ID>
<type>AA_AND2</type>
<position>-49,-572.5</position>
<input>
<ID>IN_0</ID>1070 </input>
<output>
<ID>OUT</ID>1000 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1807</ID>
<type>AE_DFF_LOW</type>
<position>-17.5,-586.5</position>
<output>
<ID>OUT_0</ID>1007 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1808</ID>
<type>AA_AND2</type>
<position>-7.5,-592</position>
<input>
<ID>IN_0</ID>1007 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1809</ID>
<type>AE_DFF_LOW</type>
<position>32,-586.5</position>
<output>
<ID>OUT_0</ID>1008 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1810</ID>
<type>AA_AND2</type>
<position>41,-593</position>
<input>
<ID>IN_0</ID>1008 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1811</ID>
<type>AE_DFF_LOW</type>
<position>80,-586.5</position>
<output>
<ID>OUT_0</ID>1010 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1812</ID>
<type>AA_AND2</type>
<position>87.5,-592</position>
<input>
<ID>IN_0</ID>1010 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1813</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-586.5</position>
<output>
<ID>OUT_0</ID>1011 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1814</ID>
<type>AA_AND2</type>
<position>138,-592</position>
<input>
<ID>IN_0</ID>1011 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1815</ID>
<type>AE_DFF_LOW</type>
<position>177.5,-586.5</position>
<output>
<ID>OUT_0</ID>1012 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1816</ID>
<type>AA_AND2</type>
<position>186,-591.5</position>
<input>
<ID>IN_0</ID>1012 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1817</ID>
<type>AE_DFF_LOW</type>
<position>235,-586.5</position>
<output>
<ID>OUT_0</ID>1013 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1818</ID>
<type>AA_AND2</type>
<position>244.5,-593.5</position>
<input>
<ID>IN_0</ID>1013 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1819</ID>
<type>AE_DFF_LOW</type>
<position>290,-586.5</position>
<output>
<ID>OUT_0</ID>1014 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1820</ID>
<type>AA_AND2</type>
<position>298,-592.5</position>
<input>
<ID>IN_0</ID>1014 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1821</ID>
<type>AE_DFF_LOW</type>
<position>347,-586.5</position>
<output>
<ID>OUT_0</ID>1015 </output>
<input>
<ID>clock</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1822</ID>
<type>AA_AND2</type>
<position>356.5,-593</position>
<input>
<ID>IN_0</ID>1015 </input>
<input>
<ID>IN_1</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1823</ID>
<type>AA_AND2</type>
<position>-49,-585.5</position>
<input>
<ID>IN_0</ID>1071 </input>
<output>
<ID>OUT</ID>1009 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1824</ID>
<type>AE_DFF_LOW</type>
<position>-17.5,-601</position>
<output>
<ID>OUT_0</ID>1016 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1825</ID>
<type>AA_AND2</type>
<position>-7.5,-606.5</position>
<input>
<ID>IN_0</ID>1016 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1826</ID>
<type>AE_DFF_LOW</type>
<position>32,-601</position>
<output>
<ID>OUT_0</ID>1017 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1827</ID>
<type>AA_AND2</type>
<position>41,-607.5</position>
<input>
<ID>IN_0</ID>1017 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1828</ID>
<type>AE_DFF_LOW</type>
<position>80,-601</position>
<output>
<ID>OUT_0</ID>1019 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1829</ID>
<type>AA_AND2</type>
<position>87.5,-606.5</position>
<input>
<ID>IN_0</ID>1019 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1830</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-601</position>
<output>
<ID>OUT_0</ID>1020 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1831</ID>
<type>AA_AND2</type>
<position>138,-606.5</position>
<input>
<ID>IN_0</ID>1020 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1832</ID>
<type>AE_DFF_LOW</type>
<position>177.5,-601</position>
<output>
<ID>OUT_0</ID>1021 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1833</ID>
<type>AA_AND2</type>
<position>186,-606</position>
<input>
<ID>IN_0</ID>1021 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1834</ID>
<type>AE_DFF_LOW</type>
<position>235,-601</position>
<output>
<ID>OUT_0</ID>1022 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1835</ID>
<type>AA_AND2</type>
<position>244.5,-608</position>
<input>
<ID>IN_0</ID>1022 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1836</ID>
<type>AE_DFF_LOW</type>
<position>290,-601</position>
<output>
<ID>OUT_0</ID>1023 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1837</ID>
<type>AA_AND2</type>
<position>298,-607</position>
<input>
<ID>IN_0</ID>1023 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1838</ID>
<type>AE_DFF_LOW</type>
<position>347,-601</position>
<output>
<ID>OUT_0</ID>1024 </output>
<input>
<ID>clock</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1839</ID>
<type>AA_AND2</type>
<position>356.5,-607.5</position>
<input>
<ID>IN_0</ID>1024 </input>
<input>
<ID>IN_1</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1840</ID>
<type>AA_AND2</type>
<position>-49,-600</position>
<input>
<ID>IN_0</ID>1072 </input>
<output>
<ID>OUT</ID>1018 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1841</ID>
<type>AE_DFF_LOW</type>
<position>-18,-613.5</position>
<output>
<ID>OUT_0</ID>1025 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1842</ID>
<type>AA_AND2</type>
<position>-8,-619</position>
<input>
<ID>IN_0</ID>1025 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1843</ID>
<type>AE_DFF_LOW</type>
<position>31.5,-613.5</position>
<output>
<ID>OUT_0</ID>1026 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1844</ID>
<type>AA_AND2</type>
<position>40.5,-620</position>
<input>
<ID>IN_0</ID>1026 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1845</ID>
<type>AE_DFF_LOW</type>
<position>79.5,-613.5</position>
<output>
<ID>OUT_0</ID>1028 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1846</ID>
<type>AA_AND2</type>
<position>87,-619</position>
<input>
<ID>IN_0</ID>1028 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1847</ID>
<type>AE_DFF_LOW</type>
<position>129,-613.5</position>
<output>
<ID>OUT_0</ID>1029 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1848</ID>
<type>AA_AND2</type>
<position>137.5,-619</position>
<input>
<ID>IN_0</ID>1029 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1849</ID>
<type>AE_DFF_LOW</type>
<position>177,-613.5</position>
<output>
<ID>OUT_0</ID>1030 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1850</ID>
<type>AA_AND2</type>
<position>185.5,-618.5</position>
<input>
<ID>IN_0</ID>1030 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1851</ID>
<type>AE_DFF_LOW</type>
<position>234.5,-613.5</position>
<output>
<ID>OUT_0</ID>1031 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1852</ID>
<type>AA_AND2</type>
<position>244,-620.5</position>
<input>
<ID>IN_0</ID>1031 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1853</ID>
<type>AE_DFF_LOW</type>
<position>289.5,-613.5</position>
<output>
<ID>OUT_0</ID>1032 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1854</ID>
<type>AA_AND2</type>
<position>297.5,-619.5</position>
<input>
<ID>IN_0</ID>1032 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1855</ID>
<type>AE_DFF_LOW</type>
<position>346.5,-613.5</position>
<output>
<ID>OUT_0</ID>1033 </output>
<input>
<ID>clock</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1856</ID>
<type>AA_AND2</type>
<position>356,-620</position>
<input>
<ID>IN_0</ID>1033 </input>
<input>
<ID>IN_1</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1857</ID>
<type>AA_AND2</type>
<position>-49.5,-612.5</position>
<input>
<ID>IN_0</ID>1073 </input>
<output>
<ID>OUT</ID>1027 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1858</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-626.5</position>
<output>
<ID>OUT_0</ID>1034 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1859</ID>
<type>AA_AND2</type>
<position>-8.5,-632</position>
<input>
<ID>IN_0</ID>1034 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1860</ID>
<type>AE_DFF_LOW</type>
<position>31,-626.5</position>
<output>
<ID>OUT_0</ID>1035 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1861</ID>
<type>AA_AND2</type>
<position>40,-633</position>
<input>
<ID>IN_0</ID>1035 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1862</ID>
<type>AE_DFF_LOW</type>
<position>79,-626.5</position>
<output>
<ID>OUT_0</ID>1037 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1863</ID>
<type>AA_AND2</type>
<position>86.5,-632</position>
<input>
<ID>IN_0</ID>1037 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1864</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-626.5</position>
<output>
<ID>OUT_0</ID>1038 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1865</ID>
<type>AA_AND2</type>
<position>137,-632</position>
<input>
<ID>IN_0</ID>1038 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1866</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-626.5</position>
<output>
<ID>OUT_0</ID>1039 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1867</ID>
<type>AA_AND2</type>
<position>185,-631.5</position>
<input>
<ID>IN_0</ID>1039 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1868</ID>
<type>AE_DFF_LOW</type>
<position>234,-626.5</position>
<output>
<ID>OUT_0</ID>1040 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1869</ID>
<type>AA_AND2</type>
<position>243.5,-633.5</position>
<input>
<ID>IN_0</ID>1040 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1870</ID>
<type>AE_DFF_LOW</type>
<position>289,-626.5</position>
<output>
<ID>OUT_0</ID>1041 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1871</ID>
<type>AA_AND2</type>
<position>297,-632.5</position>
<input>
<ID>IN_0</ID>1041 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1872</ID>
<type>AE_DFF_LOW</type>
<position>346,-626.5</position>
<output>
<ID>OUT_0</ID>1042 </output>
<input>
<ID>clock</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1873</ID>
<type>AA_AND2</type>
<position>355.5,-633</position>
<input>
<ID>IN_0</ID>1042 </input>
<input>
<ID>IN_1</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1874</ID>
<type>AA_AND2</type>
<position>-50,-625.5</position>
<input>
<ID>IN_0</ID>1074 </input>
<output>
<ID>OUT</ID>1036 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1875</ID>
<type>AE_DFF_LOW</type>
<position>-14.5,-930</position>
<output>
<ID>OUT_0</ID>1123 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>332</ID>
<type>BE_DECODER_3x8</type>
<position>-89,-621.5</position>
<input>
<ID>ENABLE</ID>3 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>1077 </output>
<output>
<ID>OUT_1</ID>1076 </output>
<output>
<ID>OUT_2</ID>1075 </output>
<output>
<ID>OUT_3</ID>1074 </output>
<output>
<ID>OUT_4</ID>1073 </output>
<output>
<ID>OUT_5</ID>1072 </output>
<output>
<ID>OUT_6</ID>1071 </output>
<output>
<ID>OUT_7</ID>1070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1876</ID>
<type>AA_AND2</type>
<position>-4.5,-935.5</position>
<input>
<ID>IN_0</ID>1123 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1877</ID>
<type>AE_DFF_LOW</type>
<position>35,-930</position>
<output>
<ID>OUT_0</ID>1124 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1878</ID>
<type>AA_AND2</type>
<position>44,-936.5</position>
<input>
<ID>IN_0</ID>1124 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1879</ID>
<type>AE_DFF_LOW</type>
<position>83,-930</position>
<output>
<ID>OUT_0</ID>1126 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1880</ID>
<type>AA_AND2</type>
<position>90.5,-935.5</position>
<input>
<ID>IN_0</ID>1126 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1881</ID>
<type>AE_DFF_LOW</type>
<position>132.5,-930</position>
<output>
<ID>OUT_0</ID>1127 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1882</ID>
<type>AA_AND2</type>
<position>141,-935.5</position>
<input>
<ID>IN_0</ID>1127 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1883</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-930</position>
<output>
<ID>OUT_0</ID>1128 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1884</ID>
<type>AA_AND2</type>
<position>189,-935</position>
<input>
<ID>IN_0</ID>1128 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1885</ID>
<type>AE_DFF_LOW</type>
<position>238,-930</position>
<output>
<ID>OUT_0</ID>1129 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1886</ID>
<type>AA_AND2</type>
<position>247.5,-937</position>
<input>
<ID>IN_0</ID>1129 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1887</ID>
<type>AE_DFF_LOW</type>
<position>293,-930</position>
<output>
<ID>OUT_0</ID>1130 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1888</ID>
<type>AA_AND2</type>
<position>301,-936</position>
<input>
<ID>IN_0</ID>1130 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1889</ID>
<type>AE_DFF_LOW</type>
<position>350,-930</position>
<output>
<ID>OUT_0</ID>1131 </output>
<input>
<ID>clock</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1890</ID>
<type>AA_AND2</type>
<position>359.5,-936.5</position>
<input>
<ID>IN_0</ID>1131 </input>
<input>
<ID>IN_1</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1891</ID>
<type>AA_AND2</type>
<position>-46,-929</position>
<input>
<ID>IN_0</ID>1155 </input>
<output>
<ID>OUT</ID>1125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1892</ID>
<type>AE_DFF_LOW</type>
<position>-14.5,-944</position>
<output>
<ID>OUT_0</ID>1132 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1893</ID>
<type>AA_AND2</type>
<position>-4.5,-949.5</position>
<input>
<ID>IN_0</ID>1132 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1894</ID>
<type>AE_DFF_LOW</type>
<position>35,-944</position>
<output>
<ID>OUT_0</ID>1133 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1895</ID>
<type>AA_AND2</type>
<position>44,-950.5</position>
<input>
<ID>IN_0</ID>1133 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1896</ID>
<type>AE_DFF_LOW</type>
<position>83,-944</position>
<output>
<ID>OUT_0</ID>1135 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1897</ID>
<type>AA_AND2</type>
<position>90.5,-949.5</position>
<input>
<ID>IN_0</ID>1135 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1898</ID>
<type>AE_DFF_LOW</type>
<position>132.5,-944</position>
<output>
<ID>OUT_0</ID>1136 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1899</ID>
<type>AA_AND2</type>
<position>141,-949.5</position>
<input>
<ID>IN_0</ID>1136 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1900</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-944</position>
<output>
<ID>OUT_0</ID>1137 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1901</ID>
<type>AA_AND2</type>
<position>189,-949</position>
<input>
<ID>IN_0</ID>1137 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1902</ID>
<type>AE_DFF_LOW</type>
<position>238,-944</position>
<output>
<ID>OUT_0</ID>1138 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1903</ID>
<type>AA_AND2</type>
<position>247.5,-951</position>
<input>
<ID>IN_0</ID>1138 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1904</ID>
<type>AE_DFF_LOW</type>
<position>293,-944</position>
<output>
<ID>OUT_0</ID>1139 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1905</ID>
<type>AA_AND2</type>
<position>301,-950</position>
<input>
<ID>IN_0</ID>1139 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1906</ID>
<type>AE_DFF_LOW</type>
<position>350,-944</position>
<output>
<ID>OUT_0</ID>1140 </output>
<input>
<ID>clock</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1907</ID>
<type>AA_AND2</type>
<position>359.5,-950.5</position>
<input>
<ID>IN_0</ID>1140 </input>
<input>
<ID>IN_1</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1908</ID>
<type>AA_AND2</type>
<position>-46,-943</position>
<input>
<ID>IN_0</ID>1156 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>1134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1909</ID>
<type>AE_DFF_LOW</type>
<position>-15,-961.5</position>
<output>
<ID>OUT_0</ID>1141 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1910</ID>
<type>AA_AND2</type>
<position>-5,-967</position>
<input>
<ID>IN_0</ID>1141 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1911</ID>
<type>AE_DFF_LOW</type>
<position>34.5,-961.5</position>
<output>
<ID>OUT_0</ID>1142 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1912</ID>
<type>AA_AND2</type>
<position>43.5,-968</position>
<input>
<ID>IN_0</ID>1142 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1913</ID>
<type>AE_DFF_LOW</type>
<position>82.5,-961.5</position>
<output>
<ID>OUT_0</ID>1144 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1914</ID>
<type>AA_AND2</type>
<position>90,-967</position>
<input>
<ID>IN_0</ID>1144 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1915</ID>
<type>AE_DFF_LOW</type>
<position>132,-961.5</position>
<output>
<ID>OUT_0</ID>1145 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1916</ID>
<type>AA_AND2</type>
<position>140.5,-967</position>
<input>
<ID>IN_0</ID>1145 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1917</ID>
<type>AE_DFF_LOW</type>
<position>180,-961.5</position>
<output>
<ID>OUT_0</ID>1146 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1918</ID>
<type>AA_AND2</type>
<position>188.5,-966.5</position>
<input>
<ID>IN_0</ID>1146 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1919</ID>
<type>AE_DFF_LOW</type>
<position>237.5,-961.5</position>
<output>
<ID>OUT_0</ID>1147 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1920</ID>
<type>AA_AND2</type>
<position>247,-968.5</position>
<input>
<ID>IN_0</ID>1147 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1921</ID>
<type>AE_DFF_LOW</type>
<position>292.5,-961.5</position>
<output>
<ID>OUT_0</ID>1148 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1922</ID>
<type>AA_AND2</type>
<position>300.5,-967.5</position>
<input>
<ID>IN_0</ID>1148 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1923</ID>
<type>AE_DFF_LOW</type>
<position>349.5,-961.5</position>
<output>
<ID>OUT_0</ID>1149 </output>
<input>
<ID>clock</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1924</ID>
<type>AA_AND2</type>
<position>359,-968</position>
<input>
<ID>IN_0</ID>1149 </input>
<input>
<ID>IN_1</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1925</ID>
<type>AA_AND2</type>
<position>-46.5,-960.5</position>
<input>
<ID>IN_0</ID>1157 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>1143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1926</ID>
<type>AE_DFF_LOW</type>
<position>-13.5,-862</position>
<output>
<ID>OUT_0</ID>1078 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1927</ID>
<type>AA_AND2</type>
<position>-3.5,-867.5</position>
<input>
<ID>IN_0</ID>1078 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1928</ID>
<type>AE_DFF_LOW</type>
<position>36,-862</position>
<output>
<ID>OUT_0</ID>1079 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1929</ID>
<type>AA_AND2</type>
<position>45,-868.5</position>
<input>
<ID>IN_0</ID>1079 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1930</ID>
<type>AE_DFF_LOW</type>
<position>84,-862</position>
<output>
<ID>OUT_0</ID>1081 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1931</ID>
<type>AA_AND2</type>
<position>91.5,-867.5</position>
<input>
<ID>IN_0</ID>1081 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1932</ID>
<type>AE_DFF_LOW</type>
<position>133.5,-862</position>
<output>
<ID>OUT_0</ID>1082 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1933</ID>
<type>AA_AND2</type>
<position>142,-867.5</position>
<input>
<ID>IN_0</ID>1082 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1934</ID>
<type>AE_DFF_LOW</type>
<position>181.5,-862</position>
<output>
<ID>OUT_0</ID>1083 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1935</ID>
<type>AA_AND2</type>
<position>190,-867</position>
<input>
<ID>IN_0</ID>1083 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1936</ID>
<type>AE_DFF_LOW</type>
<position>239,-862</position>
<output>
<ID>OUT_0</ID>1084 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1937</ID>
<type>AA_AND2</type>
<position>248.5,-869</position>
<input>
<ID>IN_0</ID>1084 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1938</ID>
<type>AE_DFF_LOW</type>
<position>294,-862</position>
<output>
<ID>OUT_0</ID>1085 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1939</ID>
<type>AA_AND2</type>
<position>302,-868</position>
<input>
<ID>IN_0</ID>1085 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1940</ID>
<type>AE_DFF_LOW</type>
<position>351,-862</position>
<output>
<ID>OUT_0</ID>1086 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1941</ID>
<type>AA_AND2</type>
<position>360.5,-868.5</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1942</ID>
<type>AA_AND2</type>
<position>-45,-861</position>
<input>
<ID>IN_0</ID>1150 </input>
<output>
<ID>OUT</ID>1080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1943</ID>
<type>AE_DFF_LOW</type>
<position>-13.5,-875</position>
<output>
<ID>OUT_0</ID>1087 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1944</ID>
<type>AA_AND2</type>
<position>-3.5,-880.5</position>
<input>
<ID>IN_0</ID>1087 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1945</ID>
<type>AE_DFF_LOW</type>
<position>36,-875</position>
<output>
<ID>OUT_0</ID>1088 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1946</ID>
<type>AA_AND2</type>
<position>45,-881.5</position>
<input>
<ID>IN_0</ID>1088 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1947</ID>
<type>AE_DFF_LOW</type>
<position>84,-875</position>
<output>
<ID>OUT_0</ID>1090 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1948</ID>
<type>AA_AND2</type>
<position>91.5,-880.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1949</ID>
<type>AE_DFF_LOW</type>
<position>133.5,-875</position>
<output>
<ID>OUT_0</ID>1091 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1950</ID>
<type>AA_AND2</type>
<position>142,-880.5</position>
<input>
<ID>IN_0</ID>1091 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1951</ID>
<type>AE_DFF_LOW</type>
<position>181.5,-875</position>
<output>
<ID>OUT_0</ID>1092 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1952</ID>
<type>AA_AND2</type>
<position>190,-880</position>
<input>
<ID>IN_0</ID>1092 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1953</ID>
<type>AE_DFF_LOW</type>
<position>239,-875</position>
<output>
<ID>OUT_0</ID>1093 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1954</ID>
<type>AA_AND2</type>
<position>248.5,-882</position>
<input>
<ID>IN_0</ID>1093 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1955</ID>
<type>AE_DFF_LOW</type>
<position>294,-875</position>
<output>
<ID>OUT_0</ID>1094 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1956</ID>
<type>AA_AND2</type>
<position>302,-881</position>
<input>
<ID>IN_0</ID>1094 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1957</ID>
<type>AE_DFF_LOW</type>
<position>351,-875</position>
<output>
<ID>OUT_0</ID>1095 </output>
<input>
<ID>clock</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1958</ID>
<type>AA_AND2</type>
<position>360.5,-881.5</position>
<input>
<ID>IN_0</ID>1095 </input>
<input>
<ID>IN_1</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1959</ID>
<type>AA_AND2</type>
<position>-45,-874</position>
<input>
<ID>IN_0</ID>1151 </input>
<output>
<ID>OUT</ID>1089 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1960</ID>
<type>AE_DFF_LOW</type>
<position>-13.5,-889.5</position>
<output>
<ID>OUT_0</ID>1096 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1961</ID>
<type>AA_AND2</type>
<position>-3.5,-895</position>
<input>
<ID>IN_0</ID>1096 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1962</ID>
<type>AE_DFF_LOW</type>
<position>36,-889.5</position>
<output>
<ID>OUT_0</ID>1097 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1963</ID>
<type>AA_AND2</type>
<position>45,-896</position>
<input>
<ID>IN_0</ID>1097 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1964</ID>
<type>AE_DFF_LOW</type>
<position>84,-889.5</position>
<output>
<ID>OUT_0</ID>1099 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1965</ID>
<type>AA_AND2</type>
<position>91.5,-895</position>
<input>
<ID>IN_0</ID>1099 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1966</ID>
<type>AE_DFF_LOW</type>
<position>133.5,-889.5</position>
<output>
<ID>OUT_0</ID>1100 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1967</ID>
<type>AA_AND2</type>
<position>142,-895</position>
<input>
<ID>IN_0</ID>1100 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1968</ID>
<type>AE_DFF_LOW</type>
<position>181.5,-889.5</position>
<output>
<ID>OUT_0</ID>1101 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1969</ID>
<type>AA_AND2</type>
<position>190,-894.5</position>
<input>
<ID>IN_0</ID>1101 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1970</ID>
<type>AE_DFF_LOW</type>
<position>239,-889.5</position>
<output>
<ID>OUT_0</ID>1102 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1971</ID>
<type>AA_AND2</type>
<position>248.5,-896.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1972</ID>
<type>AE_DFF_LOW</type>
<position>294,-889.5</position>
<output>
<ID>OUT_0</ID>1103 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1973</ID>
<type>AA_AND2</type>
<position>302,-895.5</position>
<input>
<ID>IN_0</ID>1103 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1974</ID>
<type>AE_DFF_LOW</type>
<position>351,-889.5</position>
<output>
<ID>OUT_0</ID>1104 </output>
<input>
<ID>clock</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1975</ID>
<type>AA_AND2</type>
<position>360.5,-896</position>
<input>
<ID>IN_0</ID>1104 </input>
<input>
<ID>IN_1</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1976</ID>
<type>AA_AND2</type>
<position>-45,-888.5</position>
<input>
<ID>IN_0</ID>1152 </input>
<output>
<ID>OUT</ID>1098 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1977</ID>
<type>AE_DFF_LOW</type>
<position>-14,-902</position>
<output>
<ID>OUT_0</ID>1105 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1978</ID>
<type>AA_AND2</type>
<position>-4,-907.5</position>
<input>
<ID>IN_0</ID>1105 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1979</ID>
<type>AE_DFF_LOW</type>
<position>35.5,-902</position>
<output>
<ID>OUT_0</ID>1106 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1980</ID>
<type>AA_AND2</type>
<position>44.5,-908.5</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1981</ID>
<type>AE_DFF_LOW</type>
<position>83.5,-902</position>
<output>
<ID>OUT_0</ID>1108 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1982</ID>
<type>AA_AND2</type>
<position>91,-907.5</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1983</ID>
<type>AE_DFF_LOW</type>
<position>133,-902</position>
<output>
<ID>OUT_0</ID>1109 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1984</ID>
<type>AA_AND2</type>
<position>141.5,-907.5</position>
<input>
<ID>IN_0</ID>1109 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1985</ID>
<type>AE_DFF_LOW</type>
<position>181,-902</position>
<output>
<ID>OUT_0</ID>1110 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1986</ID>
<type>AA_AND2</type>
<position>189.5,-907</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1987</ID>
<type>AE_DFF_LOW</type>
<position>238.5,-902</position>
<output>
<ID>OUT_0</ID>1111 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1988</ID>
<type>AA_AND2</type>
<position>248,-909</position>
<input>
<ID>IN_0</ID>1111 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1989</ID>
<type>AE_DFF_LOW</type>
<position>293.5,-902</position>
<output>
<ID>OUT_0</ID>1112 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1990</ID>
<type>AA_AND2</type>
<position>301.5,-908</position>
<input>
<ID>IN_0</ID>1112 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1991</ID>
<type>AE_DFF_LOW</type>
<position>350.5,-902</position>
<output>
<ID>OUT_0</ID>1113 </output>
<input>
<ID>clock</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1992</ID>
<type>AA_AND2</type>
<position>360,-908.5</position>
<input>
<ID>IN_0</ID>1113 </input>
<input>
<ID>IN_1</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1993</ID>
<type>AA_AND2</type>
<position>-45.5,-901</position>
<input>
<ID>IN_0</ID>1153 </input>
<output>
<ID>OUT</ID>1107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1994</ID>
<type>AE_DFF_LOW</type>
<position>-14.5,-915</position>
<output>
<ID>OUT_0</ID>1114 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1995</ID>
<type>AA_AND2</type>
<position>-4.5,-920.5</position>
<input>
<ID>IN_0</ID>1114 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1996</ID>
<type>AE_DFF_LOW</type>
<position>35,-915</position>
<output>
<ID>OUT_0</ID>1115 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1997</ID>
<type>AA_AND2</type>
<position>44,-921.5</position>
<input>
<ID>IN_0</ID>1115 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1998</ID>
<type>AE_DFF_LOW</type>
<position>83,-915</position>
<output>
<ID>OUT_0</ID>1117 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1999</ID>
<type>AA_AND2</type>
<position>90.5,-920.5</position>
<input>
<ID>IN_0</ID>1117 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2000</ID>
<type>AE_DFF_LOW</type>
<position>132.5,-915</position>
<output>
<ID>OUT_0</ID>1118 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2001</ID>
<type>AA_AND2</type>
<position>141,-920.5</position>
<input>
<ID>IN_0</ID>1118 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2002</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-915</position>
<output>
<ID>OUT_0</ID>1119 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2003</ID>
<type>AA_AND2</type>
<position>189,-920</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2004</ID>
<type>AE_DFF_LOW</type>
<position>238,-915</position>
<output>
<ID>OUT_0</ID>1120 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2005</ID>
<type>AA_AND2</type>
<position>247.5,-922</position>
<input>
<ID>IN_0</ID>1120 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2006</ID>
<type>AE_DFF_LOW</type>
<position>293,-915</position>
<output>
<ID>OUT_0</ID>1121 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2007</ID>
<type>AA_AND2</type>
<position>301,-921</position>
<input>
<ID>IN_0</ID>1121 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2008</ID>
<type>AE_DFF_LOW</type>
<position>350,-915</position>
<output>
<ID>OUT_0</ID>1122 </output>
<input>
<ID>clock</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2009</ID>
<type>AA_AND2</type>
<position>359.5,-921.5</position>
<input>
<ID>IN_0</ID>1122 </input>
<input>
<ID>IN_1</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2010</ID>
<type>AA_AND2</type>
<position>-46,-914</position>
<input>
<ID>IN_0</ID>1154 </input>
<output>
<ID>OUT</ID>1116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2011</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-1255.5</position>
<output>
<ID>OUT_0</ID>1203 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2012</ID>
<type>AA_AND2</type>
<position>-8.5,-1261</position>
<input>
<ID>IN_0</ID>1203 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>BE_DECODER_3x8</type>
<position>-82,-920.5</position>
<input>
<ID>ENABLE</ID>4 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>1157 </output>
<output>
<ID>OUT_1</ID>1156 </output>
<output>
<ID>OUT_2</ID>1155 </output>
<output>
<ID>OUT_3</ID>1154 </output>
<output>
<ID>OUT_4</ID>1153 </output>
<output>
<ID>OUT_5</ID>1152 </output>
<output>
<ID>OUT_6</ID>1151 </output>
<output>
<ID>OUT_7</ID>1150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2013</ID>
<type>AE_DFF_LOW</type>
<position>31,-1255.5</position>
<output>
<ID>OUT_0</ID>1204 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2014</ID>
<type>AA_AND2</type>
<position>40,-1262</position>
<input>
<ID>IN_0</ID>1204 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2015</ID>
<type>AE_DFF_LOW</type>
<position>79,-1255.5</position>
<output>
<ID>OUT_0</ID>1206 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2016</ID>
<type>AA_AND2</type>
<position>86.5,-1261</position>
<input>
<ID>IN_0</ID>1206 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2017</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-1255.5</position>
<output>
<ID>OUT_0</ID>1207 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2018</ID>
<type>AA_AND2</type>
<position>137,-1261</position>
<input>
<ID>IN_0</ID>1207 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2019</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-1255.5</position>
<output>
<ID>OUT_0</ID>1208 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2020</ID>
<type>AA_AND2</type>
<position>185,-1260.5</position>
<input>
<ID>IN_0</ID>1208 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2021</ID>
<type>AE_DFF_LOW</type>
<position>234,-1255.5</position>
<output>
<ID>OUT_0</ID>1209 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2022</ID>
<type>AA_AND2</type>
<position>243.5,-1262.5</position>
<input>
<ID>IN_0</ID>1209 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2023</ID>
<type>AE_DFF_LOW</type>
<position>289,-1255.5</position>
<output>
<ID>OUT_0</ID>1210 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2024</ID>
<type>AA_AND2</type>
<position>297,-1261.5</position>
<input>
<ID>IN_0</ID>1210 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2025</ID>
<type>AE_DFF_LOW</type>
<position>346,-1255.5</position>
<output>
<ID>OUT_0</ID>1211 </output>
<input>
<ID>clock</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2026</ID>
<type>AA_AND2</type>
<position>355.5,-1262</position>
<input>
<ID>IN_0</ID>1211 </input>
<input>
<ID>IN_1</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2027</ID>
<type>AA_AND2</type>
<position>-50,-1254.5</position>
<input>
<ID>IN_0</ID>1237 </input>
<output>
<ID>OUT</ID>1205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2028</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-1269.5</position>
<output>
<ID>OUT_0</ID>1212 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2029</ID>
<type>AA_AND2</type>
<position>-8.5,-1275</position>
<input>
<ID>IN_0</ID>1212 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2030</ID>
<type>AE_DFF_LOW</type>
<position>31,-1269.5</position>
<output>
<ID>OUT_0</ID>1213 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2031</ID>
<type>AA_AND2</type>
<position>40,-1276</position>
<input>
<ID>IN_0</ID>1213 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2032</ID>
<type>AE_DFF_LOW</type>
<position>79,-1269.5</position>
<output>
<ID>OUT_0</ID>1215 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2033</ID>
<type>AA_AND2</type>
<position>86.5,-1275</position>
<input>
<ID>IN_0</ID>1215 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2034</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-1269.5</position>
<output>
<ID>OUT_0</ID>1216 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2035</ID>
<type>AA_AND2</type>
<position>137,-1275</position>
<input>
<ID>IN_0</ID>1216 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2036</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-1269.5</position>
<output>
<ID>OUT_0</ID>1217 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2037</ID>
<type>AA_AND2</type>
<position>185,-1274.5</position>
<input>
<ID>IN_0</ID>1217 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2038</ID>
<type>AE_DFF_LOW</type>
<position>234,-1269.5</position>
<output>
<ID>OUT_0</ID>1218 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2039</ID>
<type>AA_AND2</type>
<position>243.5,-1276.5</position>
<input>
<ID>IN_0</ID>1218 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2040</ID>
<type>AE_DFF_LOW</type>
<position>289,-1269.5</position>
<output>
<ID>OUT_0</ID>1219 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2041</ID>
<type>AA_AND2</type>
<position>297,-1275.5</position>
<input>
<ID>IN_0</ID>1219 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2042</ID>
<type>AE_DFF_LOW</type>
<position>346,-1269.5</position>
<output>
<ID>OUT_0</ID>1220 </output>
<input>
<ID>clock</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2043</ID>
<type>AA_AND2</type>
<position>355.5,-1276</position>
<input>
<ID>IN_0</ID>1220 </input>
<input>
<ID>IN_1</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2044</ID>
<type>AA_AND2</type>
<position>-50,-1268.5</position>
<input>
<ID>IN_0</ID>1238 </input>
<output>
<ID>OUT</ID>1214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2045</ID>
<type>AE_DFF_LOW</type>
<position>-19,-1287</position>
<output>
<ID>OUT_0</ID>1221 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2046</ID>
<type>AA_AND2</type>
<position>-9,-1292.5</position>
<input>
<ID>IN_0</ID>1221 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2047</ID>
<type>AE_DFF_LOW</type>
<position>30.5,-1287</position>
<output>
<ID>OUT_0</ID>1222 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2048</ID>
<type>AA_AND2</type>
<position>39.5,-1293.5</position>
<input>
<ID>IN_0</ID>1222 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2049</ID>
<type>AE_DFF_LOW</type>
<position>78.5,-1287</position>
<output>
<ID>OUT_0</ID>1224 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2050</ID>
<type>AA_AND2</type>
<position>86,-1292.5</position>
<input>
<ID>IN_0</ID>1224 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2051</ID>
<type>AE_DFF_LOW</type>
<position>128,-1287</position>
<output>
<ID>OUT_0</ID>1225 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2052</ID>
<type>AA_AND2</type>
<position>136.5,-1292.5</position>
<input>
<ID>IN_0</ID>1225 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2053</ID>
<type>AE_DFF_LOW</type>
<position>176,-1287</position>
<output>
<ID>OUT_0</ID>1226 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2054</ID>
<type>AA_AND2</type>
<position>184.5,-1292</position>
<input>
<ID>IN_0</ID>1226 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2055</ID>
<type>AE_DFF_LOW</type>
<position>233.5,-1287</position>
<output>
<ID>OUT_0</ID>1227 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2056</ID>
<type>AA_AND2</type>
<position>243,-1294</position>
<input>
<ID>IN_0</ID>1227 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2057</ID>
<type>AE_DFF_LOW</type>
<position>288.5,-1287</position>
<output>
<ID>OUT_0</ID>1228 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2058</ID>
<type>AA_AND2</type>
<position>296.5,-1293</position>
<input>
<ID>IN_0</ID>1228 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2059</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-1287</position>
<output>
<ID>OUT_0</ID>1229 </output>
<input>
<ID>clock</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2060</ID>
<type>AA_AND2</type>
<position>355,-1293.5</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2061</ID>
<type>AA_AND2</type>
<position>-50.5,-1286</position>
<input>
<ID>IN_0</ID>1239 </input>
<output>
<ID>OUT</ID>1223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2062</ID>
<type>AE_DFF_LOW</type>
<position>-17.5,-1187.5</position>
<output>
<ID>OUT_0</ID>1158 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2063</ID>
<type>AA_AND2</type>
<position>-7.5,-1193</position>
<input>
<ID>IN_0</ID>1158 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2064</ID>
<type>AE_DFF_LOW</type>
<position>32,-1187.5</position>
<output>
<ID>OUT_0</ID>1159 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2065</ID>
<type>AA_AND2</type>
<position>41,-1194</position>
<input>
<ID>IN_0</ID>1159 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2066</ID>
<type>AE_DFF_LOW</type>
<position>80,-1187.5</position>
<output>
<ID>OUT_0</ID>1161 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2067</ID>
<type>AA_AND2</type>
<position>87.5,-1193</position>
<input>
<ID>IN_0</ID>1161 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2068</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-1187.5</position>
<output>
<ID>OUT_0</ID>1162 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2069</ID>
<type>AA_AND2</type>
<position>138,-1193</position>
<input>
<ID>IN_0</ID>1162 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2070</ID>
<type>AE_DFF_LOW</type>
<position>177.5,-1187.5</position>
<output>
<ID>OUT_0</ID>1163 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2071</ID>
<type>AA_AND2</type>
<position>186,-1192.5</position>
<input>
<ID>IN_0</ID>1163 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2072</ID>
<type>AE_DFF_LOW</type>
<position>235,-1187.5</position>
<output>
<ID>OUT_0</ID>1164 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2073</ID>
<type>AA_AND2</type>
<position>244.5,-1194.5</position>
<input>
<ID>IN_0</ID>1164 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2074</ID>
<type>AE_DFF_LOW</type>
<position>290,-1187.5</position>
<output>
<ID>OUT_0</ID>1165 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2075</ID>
<type>AA_AND2</type>
<position>298,-1193.5</position>
<input>
<ID>IN_0</ID>1165 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2076</ID>
<type>AE_DFF_LOW</type>
<position>347,-1187.5</position>
<output>
<ID>OUT_0</ID>1166 </output>
<input>
<ID>clock</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2077</ID>
<type>AA_AND2</type>
<position>356.5,-1194</position>
<input>
<ID>IN_0</ID>1166 </input>
<input>
<ID>IN_1</ID>1160 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2078</ID>
<type>AA_AND2</type>
<position>-49,-1186.5</position>
<input>
<ID>IN_0</ID>1230 </input>
<output>
<ID>OUT</ID>1160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2079</ID>
<type>AE_DFF_LOW</type>
<position>-17.5,-1200.5</position>
<output>
<ID>OUT_0</ID>1167 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2080</ID>
<type>AA_AND2</type>
<position>-7.5,-1206</position>
<input>
<ID>IN_0</ID>1167 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2081</ID>
<type>AE_DFF_LOW</type>
<position>32,-1200.5</position>
<output>
<ID>OUT_0</ID>1168 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2082</ID>
<type>AA_AND2</type>
<position>41,-1207</position>
<input>
<ID>IN_0</ID>1168 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2083</ID>
<type>AE_DFF_LOW</type>
<position>80,-1200.5</position>
<output>
<ID>OUT_0</ID>1170 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2084</ID>
<type>AA_AND2</type>
<position>87.5,-1206</position>
<input>
<ID>IN_0</ID>1170 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2085</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-1200.5</position>
<output>
<ID>OUT_0</ID>1171 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2086</ID>
<type>AA_AND2</type>
<position>138,-1206</position>
<input>
<ID>IN_0</ID>1171 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2087</ID>
<type>AE_DFF_LOW</type>
<position>177.5,-1200.5</position>
<output>
<ID>OUT_0</ID>1172 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2088</ID>
<type>AA_AND2</type>
<position>186,-1205.5</position>
<input>
<ID>IN_0</ID>1172 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2089</ID>
<type>AE_DFF_LOW</type>
<position>235,-1200.5</position>
<output>
<ID>OUT_0</ID>1173 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2090</ID>
<type>AA_AND2</type>
<position>244.5,-1207.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2091</ID>
<type>AE_DFF_LOW</type>
<position>290,-1200.5</position>
<output>
<ID>OUT_0</ID>1174 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2092</ID>
<type>AA_AND2</type>
<position>298,-1206.5</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2093</ID>
<type>AE_DFF_LOW</type>
<position>347,-1200.5</position>
<output>
<ID>OUT_0</ID>1175 </output>
<input>
<ID>clock</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2094</ID>
<type>AA_AND2</type>
<position>356.5,-1207</position>
<input>
<ID>IN_0</ID>1175 </input>
<input>
<ID>IN_1</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2095</ID>
<type>AA_AND2</type>
<position>-49,-1199.5</position>
<input>
<ID>IN_0</ID>1231 </input>
<output>
<ID>OUT</ID>1169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2096</ID>
<type>AE_DFF_LOW</type>
<position>-17.5,-1215</position>
<output>
<ID>OUT_0</ID>1176 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2097</ID>
<type>AA_AND2</type>
<position>-7.5,-1220.5</position>
<input>
<ID>IN_0</ID>1176 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2098</ID>
<type>AE_DFF_LOW</type>
<position>32,-1215</position>
<output>
<ID>OUT_0</ID>1177 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2099</ID>
<type>AA_AND2</type>
<position>41,-1221.5</position>
<input>
<ID>IN_0</ID>1177 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2100</ID>
<type>AE_DFF_LOW</type>
<position>80,-1215</position>
<output>
<ID>OUT_0</ID>1179 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2101</ID>
<type>AA_AND2</type>
<position>87.5,-1220.5</position>
<input>
<ID>IN_0</ID>1179 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2102</ID>
<type>AE_DFF_LOW</type>
<position>129.5,-1215</position>
<output>
<ID>OUT_0</ID>1180 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2103</ID>
<type>AA_AND2</type>
<position>138,-1220.5</position>
<input>
<ID>IN_0</ID>1180 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2104</ID>
<type>AE_DFF_LOW</type>
<position>177.5,-1215</position>
<output>
<ID>OUT_0</ID>1181 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2105</ID>
<type>AA_AND2</type>
<position>186,-1220</position>
<input>
<ID>IN_0</ID>1181 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2106</ID>
<type>AE_DFF_LOW</type>
<position>235,-1215</position>
<output>
<ID>OUT_0</ID>1182 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2107</ID>
<type>AA_AND2</type>
<position>244.5,-1222</position>
<input>
<ID>IN_0</ID>1182 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2108</ID>
<type>AE_DFF_LOW</type>
<position>290,-1215</position>
<output>
<ID>OUT_0</ID>1183 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2109</ID>
<type>AA_AND2</type>
<position>298,-1221</position>
<input>
<ID>IN_0</ID>1183 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2110</ID>
<type>AE_DFF_LOW</type>
<position>347,-1215</position>
<output>
<ID>OUT_0</ID>1184 </output>
<input>
<ID>clock</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2111</ID>
<type>AA_AND2</type>
<position>356.5,-1221.5</position>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1178 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2112</ID>
<type>AA_AND2</type>
<position>-49,-1214</position>
<input>
<ID>IN_0</ID>1232 </input>
<output>
<ID>OUT</ID>1178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2113</ID>
<type>AE_DFF_LOW</type>
<position>-18,-1227.5</position>
<output>
<ID>OUT_0</ID>1185 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2114</ID>
<type>AA_AND2</type>
<position>-8,-1233</position>
<input>
<ID>IN_0</ID>1185 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2115</ID>
<type>AE_DFF_LOW</type>
<position>31.5,-1227.5</position>
<output>
<ID>OUT_0</ID>1186 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2116</ID>
<type>AA_AND2</type>
<position>40.5,-1234</position>
<input>
<ID>IN_0</ID>1186 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2117</ID>
<type>AE_DFF_LOW</type>
<position>79.5,-1227.5</position>
<output>
<ID>OUT_0</ID>1188 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2118</ID>
<type>AA_AND2</type>
<position>87,-1233</position>
<input>
<ID>IN_0</ID>1188 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2119</ID>
<type>AE_DFF_LOW</type>
<position>129,-1227.5</position>
<output>
<ID>OUT_0</ID>1189 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2120</ID>
<type>AA_AND2</type>
<position>137.5,-1233</position>
<input>
<ID>IN_0</ID>1189 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2121</ID>
<type>AE_DFF_LOW</type>
<position>177,-1227.5</position>
<output>
<ID>OUT_0</ID>1190 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2122</ID>
<type>AA_AND2</type>
<position>185.5,-1232.5</position>
<input>
<ID>IN_0</ID>1190 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2123</ID>
<type>AE_DFF_LOW</type>
<position>234.5,-1227.5</position>
<output>
<ID>OUT_0</ID>1191 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2124</ID>
<type>AA_AND2</type>
<position>244,-1234.5</position>
<input>
<ID>IN_0</ID>1191 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2125</ID>
<type>AE_DFF_LOW</type>
<position>289.5,-1227.5</position>
<output>
<ID>OUT_0</ID>1192 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2126</ID>
<type>AA_AND2</type>
<position>297.5,-1233.5</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2127</ID>
<type>AE_DFF_LOW</type>
<position>346.5,-1227.5</position>
<output>
<ID>OUT_0</ID>1193 </output>
<input>
<ID>clock</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2128</ID>
<type>AA_AND2</type>
<position>356,-1234</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2129</ID>
<type>AA_AND2</type>
<position>-49.5,-1226.5</position>
<input>
<ID>IN_0</ID>1233 </input>
<output>
<ID>OUT</ID>1187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2130</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-1240.5</position>
<output>
<ID>OUT_0</ID>1194 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2131</ID>
<type>AA_AND2</type>
<position>-8.5,-1246</position>
<input>
<ID>IN_0</ID>1194 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2132</ID>
<type>AE_DFF_LOW</type>
<position>31,-1240.5</position>
<output>
<ID>OUT_0</ID>1195 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2133</ID>
<type>AA_AND2</type>
<position>40,-1247</position>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2134</ID>
<type>AE_DFF_LOW</type>
<position>79,-1240.5</position>
<output>
<ID>OUT_0</ID>1197 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2135</ID>
<type>AA_AND2</type>
<position>86.5,-1246</position>
<input>
<ID>IN_0</ID>1197 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2136</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-1240.5</position>
<output>
<ID>OUT_0</ID>1198 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2137</ID>
<type>AA_AND2</type>
<position>137,-1246</position>
<input>
<ID>IN_0</ID>1198 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2138</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-1240.5</position>
<output>
<ID>OUT_0</ID>1199 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2139</ID>
<type>AA_AND2</type>
<position>185,-1245.5</position>
<input>
<ID>IN_0</ID>1199 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2140</ID>
<type>AE_DFF_LOW</type>
<position>234,-1240.5</position>
<output>
<ID>OUT_0</ID>1200 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2141</ID>
<type>AA_AND2</type>
<position>243.5,-1247.5</position>
<input>
<ID>IN_0</ID>1200 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2142</ID>
<type>AE_DFF_LOW</type>
<position>289,-1240.5</position>
<output>
<ID>OUT_0</ID>1201 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2143</ID>
<type>AA_AND2</type>
<position>297,-1246.5</position>
<input>
<ID>IN_0</ID>1201 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2144</ID>
<type>AE_DFF_LOW</type>
<position>346,-1240.5</position>
<output>
<ID>OUT_0</ID>1202 </output>
<input>
<ID>clock</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2145</ID>
<type>AA_AND2</type>
<position>355.5,-1247</position>
<input>
<ID>IN_0</ID>1202 </input>
<input>
<ID>IN_1</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2146</ID>
<type>AA_AND2</type>
<position>-50,-1239.5</position>
<input>
<ID>IN_0</ID>1234 </input>
<output>
<ID>OUT</ID>1196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>606</ID>
<type>BE_DECODER_3x8</type>
<position>-89,-1238</position>
<input>
<ID>ENABLE</ID>5 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>1239 </output>
<output>
<ID>OUT_1</ID>1238 </output>
<output>
<ID>OUT_2</ID>1237 </output>
<output>
<ID>OUT_3</ID>1234 </output>
<output>
<ID>OUT_4</ID>1233 </output>
<output>
<ID>OUT_5</ID>1232 </output>
<output>
<ID>OUT_6</ID>1231 </output>
<output>
<ID>OUT_7</ID>1230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2283</ID>
<type>AE_DFF_LOW</type>
<position>-19.5,-1498.5</position>
<output>
<ID>OUT_0</ID>1357 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2284</ID>
<type>AA_AND2</type>
<position>-9.5,-1504</position>
<input>
<ID>IN_0</ID>1357 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2285</ID>
<type>AE_DFF_LOW</type>
<position>30,-1498.5</position>
<output>
<ID>OUT_0</ID>1358 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2286</ID>
<type>AA_AND2</type>
<position>39,-1505</position>
<input>
<ID>IN_0</ID>1358 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>743</ID>
<type>BE_DECODER_3x8</type>
<position>-85.5,-1474.5</position>
<input>
<ID>ENABLE</ID>1553 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>1391 </output>
<output>
<ID>OUT_1</ID>1390 </output>
<output>
<ID>OUT_2</ID>1389 </output>
<output>
<ID>OUT_3</ID>1388 </output>
<output>
<ID>OUT_4</ID>1387 </output>
<output>
<ID>OUT_5</ID>1386 </output>
<output>
<ID>OUT_6</ID>1385 </output>
<output>
<ID>OUT_7</ID>1384 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2287</ID>
<type>AE_DFF_LOW</type>
<position>78,-1498.5</position>
<output>
<ID>OUT_0</ID>1360 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2288</ID>
<type>AA_AND2</type>
<position>85.5,-1504</position>
<input>
<ID>IN_0</ID>1360 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2289</ID>
<type>AE_DFF_LOW</type>
<position>127.5,-1498.5</position>
<output>
<ID>OUT_0</ID>1361 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2290</ID>
<type>AA_AND2</type>
<position>136,-1504</position>
<input>
<ID>IN_0</ID>1361 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2291</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-1498.5</position>
<output>
<ID>OUT_0</ID>1362 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2292</ID>
<type>AA_AND2</type>
<position>184,-1503.5</position>
<input>
<ID>IN_0</ID>1362 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2293</ID>
<type>AE_DFF_LOW</type>
<position>233,-1498.5</position>
<output>
<ID>OUT_0</ID>1363 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2294</ID>
<type>AA_AND2</type>
<position>242.5,-1505.5</position>
<input>
<ID>IN_0</ID>1363 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2295</ID>
<type>AE_DFF_LOW</type>
<position>288,-1498.5</position>
<output>
<ID>OUT_0</ID>1364 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2296</ID>
<type>AA_AND2</type>
<position>296,-1504.5</position>
<input>
<ID>IN_0</ID>1364 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2297</ID>
<type>AE_DFF_LOW</type>
<position>345,-1498.5</position>
<output>
<ID>OUT_0</ID>1365 </output>
<input>
<ID>clock</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2298</ID>
<type>AA_AND2</type>
<position>354.5,-1505</position>
<input>
<ID>IN_0</ID>1365 </input>
<input>
<ID>IN_1</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2299</ID>
<type>AA_AND2</type>
<position>-51,-1497.5</position>
<input>
<ID>IN_0</ID>1389 </input>
<output>
<ID>OUT</ID>1359 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2300</ID>
<type>AE_DFF_LOW</type>
<position>-19.5,-1512.5</position>
<output>
<ID>OUT_0</ID>1366 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2301</ID>
<type>AA_AND2</type>
<position>-9.5,-1518</position>
<input>
<ID>IN_0</ID>1366 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2302</ID>
<type>AE_DFF_LOW</type>
<position>30,-1512.5</position>
<output>
<ID>OUT_0</ID>1367 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2303</ID>
<type>AA_AND2</type>
<position>39,-1519</position>
<input>
<ID>IN_0</ID>1367 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2304</ID>
<type>AE_DFF_LOW</type>
<position>78,-1512.5</position>
<output>
<ID>OUT_0</ID>1369 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2305</ID>
<type>AA_AND2</type>
<position>85.5,-1518</position>
<input>
<ID>IN_0</ID>1369 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2306</ID>
<type>AE_DFF_LOW</type>
<position>127.5,-1512.5</position>
<output>
<ID>OUT_0</ID>1370 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2307</ID>
<type>AA_AND2</type>
<position>136,-1518</position>
<input>
<ID>IN_0</ID>1370 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2308</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-1512.5</position>
<output>
<ID>OUT_0</ID>1371 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2309</ID>
<type>AA_AND2</type>
<position>184,-1517.5</position>
<input>
<ID>IN_0</ID>1371 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2310</ID>
<type>AE_DFF_LOW</type>
<position>233,-1512.5</position>
<output>
<ID>OUT_0</ID>1372 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2311</ID>
<type>AA_AND2</type>
<position>242.5,-1519.5</position>
<input>
<ID>IN_0</ID>1372 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2312</ID>
<type>AE_DFF_LOW</type>
<position>288,-1512.5</position>
<output>
<ID>OUT_0</ID>1373 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2313</ID>
<type>AA_AND2</type>
<position>296,-1518.5</position>
<input>
<ID>IN_0</ID>1373 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2314</ID>
<type>AE_DFF_LOW</type>
<position>345,-1512.5</position>
<output>
<ID>OUT_0</ID>1374 </output>
<input>
<ID>clock</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2315</ID>
<type>AA_AND2</type>
<position>354.5,-1519</position>
<input>
<ID>IN_0</ID>1374 </input>
<input>
<ID>IN_1</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2316</ID>
<type>AA_AND2</type>
<position>-51,-1511.5</position>
<input>
<ID>IN_0</ID>1390 </input>
<output>
<ID>OUT</ID>1368 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2317</ID>
<type>AE_DFF_LOW</type>
<position>-20,-1530</position>
<output>
<ID>OUT_0</ID>1375 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2318</ID>
<type>AA_AND2</type>
<position>-10,-1535.5</position>
<input>
<ID>IN_0</ID>1375 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2319</ID>
<type>AE_DFF_LOW</type>
<position>29.5,-1530</position>
<output>
<ID>OUT_0</ID>1376 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2320</ID>
<type>AA_AND2</type>
<position>38.5,-1536.5</position>
<input>
<ID>IN_0</ID>1376 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2321</ID>
<type>AE_DFF_LOW</type>
<position>77.5,-1530</position>
<output>
<ID>OUT_0</ID>1378 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2322</ID>
<type>AA_AND2</type>
<position>85,-1535.5</position>
<input>
<ID>IN_0</ID>1378 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2323</ID>
<type>AE_DFF_LOW</type>
<position>127,-1530</position>
<output>
<ID>OUT_0</ID>1379 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2324</ID>
<type>AA_AND2</type>
<position>135.5,-1535.5</position>
<input>
<ID>IN_0</ID>1379 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2325</ID>
<type>AE_DFF_LOW</type>
<position>175,-1530</position>
<output>
<ID>OUT_0</ID>1380 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2326</ID>
<type>AA_AND2</type>
<position>183.5,-1535</position>
<input>
<ID>IN_0</ID>1380 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2327</ID>
<type>AE_DFF_LOW</type>
<position>232.5,-1530</position>
<output>
<ID>OUT_0</ID>1381 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2328</ID>
<type>AA_AND2</type>
<position>242,-1537</position>
<input>
<ID>IN_0</ID>1381 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2329</ID>
<type>AE_DFF_LOW</type>
<position>287.5,-1530</position>
<output>
<ID>OUT_0</ID>1382 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2330</ID>
<type>AA_AND2</type>
<position>295.5,-1536</position>
<input>
<ID>IN_0</ID>1382 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2331</ID>
<type>AE_DFF_LOW</type>
<position>344.5,-1530</position>
<output>
<ID>OUT_0</ID>1383 </output>
<input>
<ID>clock</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2332</ID>
<type>AA_AND2</type>
<position>354,-1536.5</position>
<input>
<ID>IN_0</ID>1383 </input>
<input>
<ID>IN_1</ID>1377 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2333</ID>
<type>AA_AND2</type>
<position>-51.5,-1529</position>
<input>
<ID>IN_0</ID>1391 </input>
<output>
<ID>OUT</ID>1377 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2334</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-1430.5</position>
<output>
<ID>OUT_0</ID>1312 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2335</ID>
<type>AA_AND2</type>
<position>-8.5,-1436</position>
<input>
<ID>IN_0</ID>1312 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2336</ID>
<type>AE_DFF_LOW</type>
<position>31,-1430.5</position>
<output>
<ID>OUT_0</ID>1313 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2337</ID>
<type>AA_AND2</type>
<position>40,-1437</position>
<input>
<ID>IN_0</ID>1313 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2338</ID>
<type>AE_DFF_LOW</type>
<position>79,-1430.5</position>
<output>
<ID>OUT_0</ID>1315 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2339</ID>
<type>AA_AND2</type>
<position>86.5,-1436</position>
<input>
<ID>IN_0</ID>1315 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2340</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-1430.5</position>
<output>
<ID>OUT_0</ID>1316 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2341</ID>
<type>AA_AND2</type>
<position>137,-1436</position>
<input>
<ID>IN_0</ID>1316 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2342</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-1430.5</position>
<output>
<ID>OUT_0</ID>1317 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2343</ID>
<type>AA_AND2</type>
<position>185,-1435.5</position>
<input>
<ID>IN_0</ID>1317 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2344</ID>
<type>AE_DFF_LOW</type>
<position>234,-1430.5</position>
<output>
<ID>OUT_0</ID>1318 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2345</ID>
<type>AA_AND2</type>
<position>243.5,-1437.5</position>
<input>
<ID>IN_0</ID>1318 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2346</ID>
<type>AE_DFF_LOW</type>
<position>289,-1430.5</position>
<output>
<ID>OUT_0</ID>1319 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2347</ID>
<type>AA_AND2</type>
<position>297,-1436.5</position>
<input>
<ID>IN_0</ID>1319 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2348</ID>
<type>AE_DFF_LOW</type>
<position>346,-1430.5</position>
<output>
<ID>OUT_0</ID>1320 </output>
<input>
<ID>clock</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2349</ID>
<type>AA_AND2</type>
<position>355.5,-1437</position>
<input>
<ID>IN_0</ID>1320 </input>
<input>
<ID>IN_1</ID>1314 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2350</ID>
<type>AA_AND2</type>
<position>-50,-1429.5</position>
<input>
<ID>IN_0</ID>1384 </input>
<output>
<ID>OUT</ID>1314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2351</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-1443.5</position>
<output>
<ID>OUT_0</ID>1321 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2352</ID>
<type>AA_AND2</type>
<position>-8.5,-1449</position>
<input>
<ID>IN_0</ID>1321 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2353</ID>
<type>AE_DFF_LOW</type>
<position>31,-1443.5</position>
<output>
<ID>OUT_0</ID>1322 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2354</ID>
<type>AA_AND2</type>
<position>40,-1450</position>
<input>
<ID>IN_0</ID>1322 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2355</ID>
<type>AE_DFF_LOW</type>
<position>79,-1443.5</position>
<output>
<ID>OUT_0</ID>1324 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2356</ID>
<type>AA_AND2</type>
<position>86.5,-1449</position>
<input>
<ID>IN_0</ID>1324 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2357</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-1443.5</position>
<output>
<ID>OUT_0</ID>1325 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2358</ID>
<type>AA_AND2</type>
<position>137,-1449</position>
<input>
<ID>IN_0</ID>1325 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2359</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-1443.5</position>
<output>
<ID>OUT_0</ID>1326 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2360</ID>
<type>AA_AND2</type>
<position>185,-1448.5</position>
<input>
<ID>IN_0</ID>1326 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2361</ID>
<type>AE_DFF_LOW</type>
<position>234,-1443.5</position>
<output>
<ID>OUT_0</ID>1327 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2362</ID>
<type>AA_AND2</type>
<position>243.5,-1450.5</position>
<input>
<ID>IN_0</ID>1327 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2363</ID>
<type>AE_DFF_LOW</type>
<position>289,-1443.5</position>
<output>
<ID>OUT_0</ID>1328 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2364</ID>
<type>AA_AND2</type>
<position>297,-1449.5</position>
<input>
<ID>IN_0</ID>1328 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2365</ID>
<type>AE_DFF_LOW</type>
<position>346,-1443.5</position>
<output>
<ID>OUT_0</ID>1329 </output>
<input>
<ID>clock</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2366</ID>
<type>AA_AND2</type>
<position>355.5,-1450</position>
<input>
<ID>IN_0</ID>1329 </input>
<input>
<ID>IN_1</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2367</ID>
<type>AA_AND2</type>
<position>-50,-1442.5</position>
<input>
<ID>IN_0</ID>1385 </input>
<output>
<ID>OUT</ID>1323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2368</ID>
<type>AE_DFF_LOW</type>
<position>-18.5,-1458</position>
<output>
<ID>OUT_0</ID>1330 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2369</ID>
<type>AA_AND2</type>
<position>-8.5,-1463.5</position>
<input>
<ID>IN_0</ID>1330 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2370</ID>
<type>AE_DFF_LOW</type>
<position>31,-1458</position>
<output>
<ID>OUT_0</ID>1331 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2371</ID>
<type>AA_AND2</type>
<position>40,-1464.5</position>
<input>
<ID>IN_0</ID>1331 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2372</ID>
<type>AE_DFF_LOW</type>
<position>79,-1458</position>
<output>
<ID>OUT_0</ID>1333 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2373</ID>
<type>AA_AND2</type>
<position>86.5,-1463.5</position>
<input>
<ID>IN_0</ID>1333 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2374</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-1458</position>
<output>
<ID>OUT_0</ID>1334 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2375</ID>
<type>AA_AND2</type>
<position>137,-1463.5</position>
<input>
<ID>IN_0</ID>1334 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2376</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-1458</position>
<output>
<ID>OUT_0</ID>1335 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2377</ID>
<type>AA_AND2</type>
<position>185,-1463</position>
<input>
<ID>IN_0</ID>1335 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2378</ID>
<type>AE_DFF_LOW</type>
<position>234,-1458</position>
<output>
<ID>OUT_0</ID>1336 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2379</ID>
<type>AA_AND2</type>
<position>243.5,-1465</position>
<input>
<ID>IN_0</ID>1336 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2380</ID>
<type>AE_DFF_LOW</type>
<position>289,-1458</position>
<output>
<ID>OUT_0</ID>1337 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2381</ID>
<type>AA_AND2</type>
<position>297,-1464</position>
<input>
<ID>IN_0</ID>1337 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2382</ID>
<type>AE_DFF_LOW</type>
<position>346,-1458</position>
<output>
<ID>OUT_0</ID>1338 </output>
<input>
<ID>clock</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2383</ID>
<type>AA_AND2</type>
<position>355.5,-1464.5</position>
<input>
<ID>IN_0</ID>1338 </input>
<input>
<ID>IN_1</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2384</ID>
<type>AA_AND2</type>
<position>-50,-1457</position>
<input>
<ID>IN_0</ID>1386 </input>
<output>
<ID>OUT</ID>1332 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2385</ID>
<type>AE_DFF_LOW</type>
<position>-19,-1470.5</position>
<output>
<ID>OUT_0</ID>1339 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2386</ID>
<type>AA_AND2</type>
<position>-9,-1476</position>
<input>
<ID>IN_0</ID>1339 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2387</ID>
<type>AE_DFF_LOW</type>
<position>30.5,-1470.5</position>
<output>
<ID>OUT_0</ID>1340 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2388</ID>
<type>AA_AND2</type>
<position>39.5,-1477</position>
<input>
<ID>IN_0</ID>1340 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2389</ID>
<type>AE_DFF_LOW</type>
<position>78.5,-1470.5</position>
<output>
<ID>OUT_0</ID>1342 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2390</ID>
<type>AA_AND2</type>
<position>86,-1476</position>
<input>
<ID>IN_0</ID>1342 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2391</ID>
<type>AE_DFF_LOW</type>
<position>128,-1470.5</position>
<output>
<ID>OUT_0</ID>1343 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2392</ID>
<type>AA_AND2</type>
<position>136.5,-1476</position>
<input>
<ID>IN_0</ID>1343 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2393</ID>
<type>AE_DFF_LOW</type>
<position>176,-1470.5</position>
<output>
<ID>OUT_0</ID>1344 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2394</ID>
<type>AA_AND2</type>
<position>184.5,-1475.5</position>
<input>
<ID>IN_0</ID>1344 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2395</ID>
<type>AE_DFF_LOW</type>
<position>233.5,-1470.5</position>
<output>
<ID>OUT_0</ID>1345 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2396</ID>
<type>AA_AND2</type>
<position>243,-1477.5</position>
<input>
<ID>IN_0</ID>1345 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2397</ID>
<type>AE_DFF_LOW</type>
<position>288.5,-1470.5</position>
<output>
<ID>OUT_0</ID>1346 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2398</ID>
<type>AA_AND2</type>
<position>296.5,-1476.5</position>
<input>
<ID>IN_0</ID>1346 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2399</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-1470.5</position>
<output>
<ID>OUT_0</ID>1347 </output>
<input>
<ID>clock</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2400</ID>
<type>AA_AND2</type>
<position>355,-1477</position>
<input>
<ID>IN_0</ID>1347 </input>
<input>
<ID>IN_1</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2401</ID>
<type>AA_AND2</type>
<position>-50.5,-1469.5</position>
<input>
<ID>IN_0</ID>1387 </input>
<output>
<ID>OUT</ID>1341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2402</ID>
<type>AE_DFF_LOW</type>
<position>-19.5,-1483.5</position>
<output>
<ID>OUT_0</ID>1348 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2403</ID>
<type>AA_AND2</type>
<position>-9.5,-1489</position>
<input>
<ID>IN_0</ID>1348 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2404</ID>
<type>AE_DFF_LOW</type>
<position>30,-1483.5</position>
<output>
<ID>OUT_0</ID>1349 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2405</ID>
<type>AA_AND2</type>
<position>39,-1490</position>
<input>
<ID>IN_0</ID>1349 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2406</ID>
<type>AE_DFF_LOW</type>
<position>78,-1483.5</position>
<output>
<ID>OUT_0</ID>1351 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2407</ID>
<type>AA_AND2</type>
<position>85.5,-1489</position>
<input>
<ID>IN_0</ID>1351 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2408</ID>
<type>AE_DFF_LOW</type>
<position>127.5,-1483.5</position>
<output>
<ID>OUT_0</ID>1352 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2409</ID>
<type>AA_AND2</type>
<position>136,-1489</position>
<input>
<ID>IN_0</ID>1352 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2410</ID>
<type>AE_DFF_LOW</type>
<position>175.5,-1483.5</position>
<output>
<ID>OUT_0</ID>1353 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2411</ID>
<type>AA_AND2</type>
<position>184,-1488.5</position>
<input>
<ID>IN_0</ID>1353 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2412</ID>
<type>AE_DFF_LOW</type>
<position>233,-1483.5</position>
<output>
<ID>OUT_0</ID>1354 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2413</ID>
<type>AA_AND2</type>
<position>242.5,-1490.5</position>
<input>
<ID>IN_0</ID>1354 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2414</ID>
<type>AE_DFF_LOW</type>
<position>288,-1483.5</position>
<output>
<ID>OUT_0</ID>1355 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2415</ID>
<type>AA_AND2</type>
<position>296,-1489.5</position>
<input>
<ID>IN_0</ID>1355 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2416</ID>
<type>AE_DFF_LOW</type>
<position>345,-1483.5</position>
<output>
<ID>OUT_0</ID>1356 </output>
<input>
<ID>clock</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2417</ID>
<type>AA_AND2</type>
<position>354.5,-1490</position>
<input>
<ID>IN_0</ID>1356 </input>
<input>
<ID>IN_1</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2418</ID>
<type>AA_AND2</type>
<position>-51,-1482.5</position>
<input>
<ID>IN_0</ID>1388 </input>
<output>
<ID>OUT</ID>1350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2419</ID>
<type>AE_DFF_LOW</type>
<position>-21.5,-1790</position>
<output>
<ID>OUT_0</ID>1437 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2420</ID>
<type>AA_AND2</type>
<position>-11.5,-1795.5</position>
<input>
<ID>IN_0</ID>1437 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2421</ID>
<type>AE_DFF_LOW</type>
<position>28,-1790</position>
<output>
<ID>OUT_0</ID>1438 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2422</ID>
<type>AA_AND2</type>
<position>37,-1796.5</position>
<input>
<ID>IN_0</ID>1438 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2423</ID>
<type>AE_DFF_LOW</type>
<position>76,-1790</position>
<output>
<ID>OUT_0</ID>1440 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>880</ID>
<type>BE_DECODER_3x8</type>
<position>-89.5,-1769</position>
<input>
<ID>ENABLE</ID>1554 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>1471 </output>
<output>
<ID>OUT_1</ID>1470 </output>
<output>
<ID>OUT_2</ID>1469 </output>
<output>
<ID>OUT_3</ID>1468 </output>
<output>
<ID>OUT_4</ID>1467 </output>
<output>
<ID>OUT_5</ID>1466 </output>
<output>
<ID>OUT_6</ID>1465 </output>
<output>
<ID>OUT_7</ID>1464 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2424</ID>
<type>AA_AND2</type>
<position>83.5,-1795.5</position>
<input>
<ID>IN_0</ID>1440 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2425</ID>
<type>AE_DFF_LOW</type>
<position>125.5,-1790</position>
<output>
<ID>OUT_0</ID>1441 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2426</ID>
<type>AA_AND2</type>
<position>134,-1795.5</position>
<input>
<ID>IN_0</ID>1441 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2427</ID>
<type>AE_DFF_LOW</type>
<position>173.5,-1790</position>
<output>
<ID>OUT_0</ID>1442 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2428</ID>
<type>AA_AND2</type>
<position>182,-1795</position>
<input>
<ID>IN_0</ID>1442 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2429</ID>
<type>AE_DFF_LOW</type>
<position>231,-1790</position>
<output>
<ID>OUT_0</ID>1443 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2430</ID>
<type>AA_AND2</type>
<position>240.5,-1797</position>
<input>
<ID>IN_0</ID>1443 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2431</ID>
<type>AE_DFF_LOW</type>
<position>286,-1790</position>
<output>
<ID>OUT_0</ID>1444 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2432</ID>
<type>AA_AND2</type>
<position>294,-1796</position>
<input>
<ID>IN_0</ID>1444 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2433</ID>
<type>AE_DFF_LOW</type>
<position>343,-1790</position>
<output>
<ID>OUT_0</ID>1445 </output>
<input>
<ID>clock</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2434</ID>
<type>AA_AND2</type>
<position>352.5,-1796.5</position>
<input>
<ID>IN_0</ID>1445 </input>
<input>
<ID>IN_1</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2435</ID>
<type>AA_AND2</type>
<position>-53,-1789</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT</ID>1439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2436</ID>
<type>AE_DFF_LOW</type>
<position>-21.5,-1804</position>
<output>
<ID>OUT_0</ID>1446 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2437</ID>
<type>AA_AND2</type>
<position>-11.5,-1809.5</position>
<input>
<ID>IN_0</ID>1446 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2438</ID>
<type>AE_DFF_LOW</type>
<position>28,-1804</position>
<output>
<ID>OUT_0</ID>1447 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2439</ID>
<type>AA_AND2</type>
<position>37,-1810.5</position>
<input>
<ID>IN_0</ID>1447 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2440</ID>
<type>AE_DFF_LOW</type>
<position>76,-1804</position>
<output>
<ID>OUT_0</ID>1449 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2441</ID>
<type>AA_AND2</type>
<position>83.5,-1809.5</position>
<input>
<ID>IN_0</ID>1449 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2442</ID>
<type>AE_DFF_LOW</type>
<position>125.5,-1804</position>
<output>
<ID>OUT_0</ID>1450 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2443</ID>
<type>AA_AND2</type>
<position>134,-1809.5</position>
<input>
<ID>IN_0</ID>1450 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2444</ID>
<type>AE_DFF_LOW</type>
<position>173.5,-1804</position>
<output>
<ID>OUT_0</ID>1451 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2445</ID>
<type>AA_AND2</type>
<position>182,-1809</position>
<input>
<ID>IN_0</ID>1451 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2446</ID>
<type>AE_DFF_LOW</type>
<position>231,-1804</position>
<output>
<ID>OUT_0</ID>1452 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2447</ID>
<type>AA_AND2</type>
<position>240.5,-1811</position>
<input>
<ID>IN_0</ID>1452 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2448</ID>
<type>AE_DFF_LOW</type>
<position>286,-1804</position>
<output>
<ID>OUT_0</ID>1453 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2449</ID>
<type>AA_AND2</type>
<position>294,-1810</position>
<input>
<ID>IN_0</ID>1453 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2450</ID>
<type>AE_DFF_LOW</type>
<position>343,-1804</position>
<output>
<ID>OUT_0</ID>1454 </output>
<input>
<ID>clock</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2451</ID>
<type>AA_AND2</type>
<position>352.5,-1810.5</position>
<input>
<ID>IN_0</ID>1454 </input>
<input>
<ID>IN_1</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2452</ID>
<type>AA_AND2</type>
<position>-53,-1803</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT</ID>1448 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2453</ID>
<type>AE_DFF_LOW</type>
<position>-22,-1821.5</position>
<output>
<ID>OUT_0</ID>1455 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2454</ID>
<type>AA_AND2</type>
<position>-12,-1827</position>
<input>
<ID>IN_0</ID>1455 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2455</ID>
<type>AE_DFF_LOW</type>
<position>27.5,-1821.5</position>
<output>
<ID>OUT_0</ID>1456 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2456</ID>
<type>AA_AND2</type>
<position>36.5,-1828</position>
<input>
<ID>IN_0</ID>1456 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2457</ID>
<type>AE_DFF_LOW</type>
<position>75.5,-1821.5</position>
<output>
<ID>OUT_0</ID>1458 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2458</ID>
<type>AA_AND2</type>
<position>83,-1827</position>
<input>
<ID>IN_0</ID>1458 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2459</ID>
<type>AE_DFF_LOW</type>
<position>125,-1821.5</position>
<output>
<ID>OUT_0</ID>1459 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2460</ID>
<type>AA_AND2</type>
<position>133.5,-1827</position>
<input>
<ID>IN_0</ID>1459 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2461</ID>
<type>AE_DFF_LOW</type>
<position>173,-1821.5</position>
<output>
<ID>OUT_0</ID>1460 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2462</ID>
<type>AA_AND2</type>
<position>181.5,-1826.5</position>
<input>
<ID>IN_0</ID>1460 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2463</ID>
<type>AE_DFF_LOW</type>
<position>230.5,-1821.5</position>
<output>
<ID>OUT_0</ID>1461 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2464</ID>
<type>AA_AND2</type>
<position>240,-1828.5</position>
<input>
<ID>IN_0</ID>1461 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2465</ID>
<type>AE_DFF_LOW</type>
<position>285.5,-1821.5</position>
<output>
<ID>OUT_0</ID>1462 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2466</ID>
<type>AA_AND2</type>
<position>293.5,-1827.5</position>
<input>
<ID>IN_0</ID>1462 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2467</ID>
<type>AE_DFF_LOW</type>
<position>342.5,-1821.5</position>
<output>
<ID>OUT_0</ID>1463 </output>
<input>
<ID>clock</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2468</ID>
<type>AA_AND2</type>
<position>352,-1828</position>
<input>
<ID>IN_0</ID>1463 </input>
<input>
<ID>IN_1</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2469</ID>
<type>AA_AND2</type>
<position>-53.5,-1820.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT</ID>1457 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2470</ID>
<type>AE_DFF_LOW</type>
<position>-20.5,-1722</position>
<output>
<ID>OUT_0</ID>1392 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2471</ID>
<type>AA_AND2</type>
<position>-10.5,-1727.5</position>
<input>
<ID>IN_0</ID>1392 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2472</ID>
<type>AE_DFF_LOW</type>
<position>29,-1722</position>
<output>
<ID>OUT_0</ID>1393 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2473</ID>
<type>AA_AND2</type>
<position>38,-1728.5</position>
<input>
<ID>IN_0</ID>1393 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2474</ID>
<type>AE_DFF_LOW</type>
<position>77,-1722</position>
<output>
<ID>OUT_0</ID>1395 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2475</ID>
<type>AA_AND2</type>
<position>84.5,-1727.5</position>
<input>
<ID>IN_0</ID>1395 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2476</ID>
<type>AE_DFF_LOW</type>
<position>126.5,-1722</position>
<output>
<ID>OUT_0</ID>1396 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2477</ID>
<type>AA_AND2</type>
<position>135,-1727.5</position>
<input>
<ID>IN_0</ID>1396 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2478</ID>
<type>AE_DFF_LOW</type>
<position>174.5,-1722</position>
<output>
<ID>OUT_0</ID>1397 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2479</ID>
<type>AA_AND2</type>
<position>183,-1727</position>
<input>
<ID>IN_0</ID>1397 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2480</ID>
<type>AE_DFF_LOW</type>
<position>232,-1722</position>
<output>
<ID>OUT_0</ID>1398 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2481</ID>
<type>AA_AND2</type>
<position>241.5,-1729</position>
<input>
<ID>IN_0</ID>1398 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2482</ID>
<type>AE_DFF_LOW</type>
<position>287,-1722</position>
<output>
<ID>OUT_0</ID>1399 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2483</ID>
<type>AA_AND2</type>
<position>295,-1728</position>
<input>
<ID>IN_0</ID>1399 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2484</ID>
<type>AE_DFF_LOW</type>
<position>344,-1722</position>
<output>
<ID>OUT_0</ID>1400 </output>
<input>
<ID>clock</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2485</ID>
<type>AA_AND2</type>
<position>353.5,-1728.5</position>
<input>
<ID>IN_0</ID>1400 </input>
<input>
<ID>IN_1</ID>1394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2486</ID>
<type>AA_AND2</type>
<position>-52,-1721</position>
<input>
<ID>IN_0</ID>1464 </input>
<output>
<ID>OUT</ID>1394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2487</ID>
<type>AE_DFF_LOW</type>
<position>-20.5,-1735</position>
<output>
<ID>OUT_0</ID>1401 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2488</ID>
<type>AA_AND2</type>
<position>-10.5,-1740.5</position>
<input>
<ID>IN_0</ID>1401 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2489</ID>
<type>AE_DFF_LOW</type>
<position>29,-1735</position>
<output>
<ID>OUT_0</ID>1402 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2490</ID>
<type>AA_AND2</type>
<position>38,-1741.5</position>
<input>
<ID>IN_0</ID>1402 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2491</ID>
<type>AE_DFF_LOW</type>
<position>77,-1735</position>
<output>
<ID>OUT_0</ID>1404 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2492</ID>
<type>AA_AND2</type>
<position>84.5,-1740.5</position>
<input>
<ID>IN_0</ID>1404 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2493</ID>
<type>AE_DFF_LOW</type>
<position>126.5,-1735</position>
<output>
<ID>OUT_0</ID>1405 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2494</ID>
<type>AA_AND2</type>
<position>135,-1740.5</position>
<input>
<ID>IN_0</ID>1405 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2495</ID>
<type>AE_DFF_LOW</type>
<position>174.5,-1735</position>
<output>
<ID>OUT_0</ID>1406 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2496</ID>
<type>AA_AND2</type>
<position>183,-1740</position>
<input>
<ID>IN_0</ID>1406 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2497</ID>
<type>AE_DFF_LOW</type>
<position>232,-1735</position>
<output>
<ID>OUT_0</ID>1407 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2498</ID>
<type>AA_AND2</type>
<position>241.5,-1742</position>
<input>
<ID>IN_0</ID>1407 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2499</ID>
<type>AE_DFF_LOW</type>
<position>287,-1735</position>
<output>
<ID>OUT_0</ID>1408 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2500</ID>
<type>AA_AND2</type>
<position>295,-1741</position>
<input>
<ID>IN_0</ID>1408 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2501</ID>
<type>AE_DFF_LOW</type>
<position>344,-1735</position>
<output>
<ID>OUT_0</ID>1409 </output>
<input>
<ID>clock</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2502</ID>
<type>AA_AND2</type>
<position>353.5,-1741.5</position>
<input>
<ID>IN_0</ID>1409 </input>
<input>
<ID>IN_1</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2503</ID>
<type>AA_AND2</type>
<position>-52,-1734</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT</ID>1403 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2504</ID>
<type>AE_DFF_LOW</type>
<position>-20.5,-1749.5</position>
<output>
<ID>OUT_0</ID>1410 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2505</ID>
<type>AA_AND2</type>
<position>-10.5,-1755</position>
<input>
<ID>IN_0</ID>1410 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2506</ID>
<type>AE_DFF_LOW</type>
<position>29,-1749.5</position>
<output>
<ID>OUT_0</ID>1411 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2507</ID>
<type>AA_AND2</type>
<position>38,-1756</position>
<input>
<ID>IN_0</ID>1411 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2508</ID>
<type>AE_DFF_LOW</type>
<position>77,-1749.5</position>
<output>
<ID>OUT_0</ID>1413 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2509</ID>
<type>AA_AND2</type>
<position>84.5,-1755</position>
<input>
<ID>IN_0</ID>1413 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2510</ID>
<type>AE_DFF_LOW</type>
<position>126.5,-1749.5</position>
<output>
<ID>OUT_0</ID>1414 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2511</ID>
<type>AA_AND2</type>
<position>135,-1755</position>
<input>
<ID>IN_0</ID>1414 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2512</ID>
<type>AE_DFF_LOW</type>
<position>174.5,-1749.5</position>
<output>
<ID>OUT_0</ID>1415 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2513</ID>
<type>AA_AND2</type>
<position>183,-1754.5</position>
<input>
<ID>IN_0</ID>1415 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2514</ID>
<type>AE_DFF_LOW</type>
<position>232,-1749.5</position>
<output>
<ID>OUT_0</ID>1416 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2515</ID>
<type>AA_AND2</type>
<position>241.5,-1756.5</position>
<input>
<ID>IN_0</ID>1416 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2516</ID>
<type>AE_DFF_LOW</type>
<position>287,-1749.5</position>
<output>
<ID>OUT_0</ID>1417 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2517</ID>
<type>AA_AND2</type>
<position>295,-1755.5</position>
<input>
<ID>IN_0</ID>1417 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2518</ID>
<type>AE_DFF_LOW</type>
<position>344,-1749.5</position>
<output>
<ID>OUT_0</ID>1418 </output>
<input>
<ID>clock</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2519</ID>
<type>AA_AND2</type>
<position>353.5,-1756</position>
<input>
<ID>IN_0</ID>1418 </input>
<input>
<ID>IN_1</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2520</ID>
<type>AA_AND2</type>
<position>-52,-1748.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT</ID>1412 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2521</ID>
<type>AE_DFF_LOW</type>
<position>-21,-1762</position>
<output>
<ID>OUT_0</ID>1419 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2522</ID>
<type>AA_AND2</type>
<position>-11,-1767.5</position>
<input>
<ID>IN_0</ID>1419 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2523</ID>
<type>AE_DFF_LOW</type>
<position>28.5,-1762</position>
<output>
<ID>OUT_0</ID>1420 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2524</ID>
<type>AA_AND2</type>
<position>37.5,-1768.5</position>
<input>
<ID>IN_0</ID>1420 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2525</ID>
<type>AE_DFF_LOW</type>
<position>76.5,-1762</position>
<output>
<ID>OUT_0</ID>1422 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2526</ID>
<type>AA_AND2</type>
<position>84,-1767.5</position>
<input>
<ID>IN_0</ID>1422 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2527</ID>
<type>AE_DFF_LOW</type>
<position>126,-1762</position>
<output>
<ID>OUT_0</ID>1423 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2528</ID>
<type>AA_AND2</type>
<position>134.5,-1767.5</position>
<input>
<ID>IN_0</ID>1423 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2529</ID>
<type>AE_DFF_LOW</type>
<position>174,-1762</position>
<output>
<ID>OUT_0</ID>1424 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2530</ID>
<type>AA_AND2</type>
<position>182.5,-1767</position>
<input>
<ID>IN_0</ID>1424 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2531</ID>
<type>AE_DFF_LOW</type>
<position>231.5,-1762</position>
<output>
<ID>OUT_0</ID>1425 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2532</ID>
<type>AA_AND2</type>
<position>241,-1769</position>
<input>
<ID>IN_0</ID>1425 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2533</ID>
<type>AE_DFF_LOW</type>
<position>286.5,-1762</position>
<output>
<ID>OUT_0</ID>1426 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2534</ID>
<type>AA_AND2</type>
<position>294.5,-1768</position>
<input>
<ID>IN_0</ID>1426 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2535</ID>
<type>AE_DFF_LOW</type>
<position>343.5,-1762</position>
<output>
<ID>OUT_0</ID>1427 </output>
<input>
<ID>clock</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2536</ID>
<type>AA_AND2</type>
<position>353,-1768.5</position>
<input>
<ID>IN_0</ID>1427 </input>
<input>
<ID>IN_1</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2537</ID>
<type>AA_AND2</type>
<position>-52.5,-1761</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT</ID>1421 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2538</ID>
<type>AE_DFF_LOW</type>
<position>-21.5,-1775</position>
<output>
<ID>OUT_0</ID>1428 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2539</ID>
<type>AA_AND2</type>
<position>-11.5,-1780.5</position>
<input>
<ID>IN_0</ID>1428 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2540</ID>
<type>AE_DFF_LOW</type>
<position>28,-1775</position>
<output>
<ID>OUT_0</ID>1429 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2541</ID>
<type>AA_AND2</type>
<position>37,-1781.5</position>
<input>
<ID>IN_0</ID>1429 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2542</ID>
<type>AE_DFF_LOW</type>
<position>76,-1775</position>
<output>
<ID>OUT_0</ID>1431 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2543</ID>
<type>AA_AND2</type>
<position>83.5,-1780.5</position>
<input>
<ID>IN_0</ID>1431 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2544</ID>
<type>AE_DFF_LOW</type>
<position>125.5,-1775</position>
<output>
<ID>OUT_0</ID>1432 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2545</ID>
<type>AA_AND2</type>
<position>134,-1780.5</position>
<input>
<ID>IN_0</ID>1432 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2546</ID>
<type>AE_DFF_LOW</type>
<position>173.5,-1775</position>
<output>
<ID>OUT_0</ID>1433 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2547</ID>
<type>AA_AND2</type>
<position>182,-1780</position>
<input>
<ID>IN_0</ID>1433 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2548</ID>
<type>AE_DFF_LOW</type>
<position>231,-1775</position>
<output>
<ID>OUT_0</ID>1434 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2549</ID>
<type>AA_AND2</type>
<position>240.5,-1782</position>
<input>
<ID>IN_0</ID>1434 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2550</ID>
<type>AE_DFF_LOW</type>
<position>286,-1775</position>
<output>
<ID>OUT_0</ID>1435 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2551</ID>
<type>AA_AND2</type>
<position>294,-1781</position>
<input>
<ID>IN_0</ID>1435 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2552</ID>
<type>AE_DFF_LOW</type>
<position>343,-1775</position>
<output>
<ID>OUT_0</ID>1436 </output>
<input>
<ID>clock</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2553</ID>
<type>AA_AND2</type>
<position>352.5,-1781.5</position>
<input>
<ID>IN_0</ID>1436 </input>
<input>
<ID>IN_1</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2554</ID>
<type>AA_AND2</type>
<position>-53,-1774</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT</ID>1430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2555</ID>
<type>AE_DFF_LOW</type>
<position>-16.5,-2083.5</position>
<output>
<ID>OUT_0</ID>1517 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2556</ID>
<type>AA_AND2</type>
<position>-6.5,-2089</position>
<input>
<ID>IN_0</ID>1517 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2557</ID>
<type>AE_DFF_LOW</type>
<position>33,-2083.5</position>
<output>
<ID>OUT_0</ID>1518 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2558</ID>
<type>AA_AND2</type>
<position>42,-2090</position>
<input>
<ID>IN_0</ID>1518 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2559</ID>
<type>AE_DFF_LOW</type>
<position>81,-2083.5</position>
<output>
<ID>OUT_0</ID>1520 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2560</ID>
<type>AA_AND2</type>
<position>88.5,-2089</position>
<input>
<ID>IN_0</ID>1520 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1017</ID>
<type>BE_DECODER_3x8</type>
<position>-86.5,-2067</position>
<input>
<ID>ENABLE</ID>1555 </input>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>671 </input>
<output>
<ID>OUT_0</ID>1551 </output>
<output>
<ID>OUT_1</ID>1550 </output>
<output>
<ID>OUT_2</ID>1549 </output>
<output>
<ID>OUT_3</ID>1548 </output>
<output>
<ID>OUT_4</ID>1547 </output>
<output>
<ID>OUT_5</ID>1546 </output>
<output>
<ID>OUT_6</ID>1545 </output>
<output>
<ID>OUT_7</ID>1544 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2561</ID>
<type>AE_DFF_LOW</type>
<position>130.5,-2083.5</position>
<output>
<ID>OUT_0</ID>1521 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2562</ID>
<type>AA_AND2</type>
<position>139,-2089</position>
<input>
<ID>IN_0</ID>1521 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2563</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-2083.5</position>
<output>
<ID>OUT_0</ID>1522 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2564</ID>
<type>AA_AND2</type>
<position>187,-2088.5</position>
<input>
<ID>IN_0</ID>1522 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2565</ID>
<type>AE_DFF_LOW</type>
<position>236,-2083.5</position>
<output>
<ID>OUT_0</ID>1523 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2566</ID>
<type>AA_AND2</type>
<position>245.5,-2090.5</position>
<input>
<ID>IN_0</ID>1523 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2567</ID>
<type>AE_DFF_LOW</type>
<position>291,-2083.5</position>
<output>
<ID>OUT_0</ID>1524 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2568</ID>
<type>AA_AND2</type>
<position>299,-2089.5</position>
<input>
<ID>IN_0</ID>1524 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2569</ID>
<type>AE_DFF_LOW</type>
<position>348,-2083.5</position>
<output>
<ID>OUT_0</ID>1525 </output>
<input>
<ID>clock</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2570</ID>
<type>AA_AND2</type>
<position>357.5,-2090</position>
<input>
<ID>IN_0</ID>1525 </input>
<input>
<ID>IN_1</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2571</ID>
<type>AA_AND2</type>
<position>-48,-2082.5</position>
<input>
<ID>IN_0</ID>1549 </input>
<output>
<ID>OUT</ID>1519 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2572</ID>
<type>AE_DFF_LOW</type>
<position>-16.5,-2097.5</position>
<output>
<ID>OUT_0</ID>1526 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2573</ID>
<type>AA_AND2</type>
<position>-6.5,-2103</position>
<input>
<ID>IN_0</ID>1526 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2574</ID>
<type>AE_DFF_LOW</type>
<position>33,-2097.5</position>
<output>
<ID>OUT_0</ID>1527 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2575</ID>
<type>AA_AND2</type>
<position>42,-2104</position>
<input>
<ID>IN_0</ID>1527 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2576</ID>
<type>AE_DFF_LOW</type>
<position>81,-2097.5</position>
<output>
<ID>OUT_0</ID>1529 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2577</ID>
<type>AA_AND2</type>
<position>88.5,-2103</position>
<input>
<ID>IN_0</ID>1529 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2578</ID>
<type>AE_DFF_LOW</type>
<position>130.5,-2097.5</position>
<output>
<ID>OUT_0</ID>1530 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2579</ID>
<type>AA_AND2</type>
<position>139,-2103</position>
<input>
<ID>IN_0</ID>1530 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2580</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-2097.5</position>
<output>
<ID>OUT_0</ID>1531 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2581</ID>
<type>AA_AND2</type>
<position>187,-2102.5</position>
<input>
<ID>IN_0</ID>1531 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2582</ID>
<type>AE_DFF_LOW</type>
<position>236,-2097.5</position>
<output>
<ID>OUT_0</ID>1532 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2583</ID>
<type>AA_AND2</type>
<position>245.5,-2104.5</position>
<input>
<ID>IN_0</ID>1532 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2584</ID>
<type>AE_DFF_LOW</type>
<position>291,-2097.5</position>
<output>
<ID>OUT_0</ID>1533 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2585</ID>
<type>AA_AND2</type>
<position>299,-2103.5</position>
<input>
<ID>IN_0</ID>1533 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2586</ID>
<type>AE_DFF_LOW</type>
<position>348,-2097.5</position>
<output>
<ID>OUT_0</ID>1534 </output>
<input>
<ID>clock</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2587</ID>
<type>AA_AND2</type>
<position>357.5,-2104</position>
<input>
<ID>IN_0</ID>1534 </input>
<input>
<ID>IN_1</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2588</ID>
<type>AA_AND2</type>
<position>-48,-2096.5</position>
<input>
<ID>IN_0</ID>1550 </input>
<output>
<ID>OUT</ID>1528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2589</ID>
<type>AE_DFF_LOW</type>
<position>-17,-2115</position>
<output>
<ID>OUT_0</ID>1535 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2590</ID>
<type>AA_AND2</type>
<position>-7,-2120.5</position>
<input>
<ID>IN_0</ID>1535 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2591</ID>
<type>AE_DFF_LOW</type>
<position>32.5,-2115</position>
<output>
<ID>OUT_0</ID>1536 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2592</ID>
<type>AA_AND2</type>
<position>41.5,-2121.5</position>
<input>
<ID>IN_0</ID>1536 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2593</ID>
<type>AE_DFF_LOW</type>
<position>80.5,-2115</position>
<output>
<ID>OUT_0</ID>1538 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2594</ID>
<type>AA_AND2</type>
<position>88,-2120.5</position>
<input>
<ID>IN_0</ID>1538 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2595</ID>
<type>AE_DFF_LOW</type>
<position>130,-2115</position>
<output>
<ID>OUT_0</ID>1539 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2596</ID>
<type>AA_AND2</type>
<position>138.5,-2120.5</position>
<input>
<ID>IN_0</ID>1539 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2597</ID>
<type>AE_DFF_LOW</type>
<position>178,-2115</position>
<output>
<ID>OUT_0</ID>1540 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2598</ID>
<type>AA_AND2</type>
<position>186.5,-2120</position>
<input>
<ID>IN_0</ID>1540 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2599</ID>
<type>AE_DFF_LOW</type>
<position>235.5,-2115</position>
<output>
<ID>OUT_0</ID>1541 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2600</ID>
<type>AA_AND2</type>
<position>245,-2122</position>
<input>
<ID>IN_0</ID>1541 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2601</ID>
<type>AE_DFF_LOW</type>
<position>290.5,-2115</position>
<output>
<ID>OUT_0</ID>1542 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2602</ID>
<type>AA_AND2</type>
<position>298.5,-2121</position>
<input>
<ID>IN_0</ID>1542 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2603</ID>
<type>AE_DFF_LOW</type>
<position>347.5,-2115</position>
<output>
<ID>OUT_0</ID>1543 </output>
<input>
<ID>clock</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2604</ID>
<type>AA_AND2</type>
<position>357,-2121.5</position>
<input>
<ID>IN_0</ID>1543 </input>
<input>
<ID>IN_1</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2605</ID>
<type>AA_AND2</type>
<position>-48.5,-2114</position>
<input>
<ID>IN_0</ID>1551 </input>
<output>
<ID>OUT</ID>1537 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2606</ID>
<type>AE_DFF_LOW</type>
<position>-15.5,-2015.5</position>
<output>
<ID>OUT_0</ID>1472 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2607</ID>
<type>AA_AND2</type>
<position>-5.5,-2021</position>
<input>
<ID>IN_0</ID>1472 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2608</ID>
<type>AE_DFF_LOW</type>
<position>34,-2015.5</position>
<output>
<ID>OUT_0</ID>1473 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2609</ID>
<type>AA_AND2</type>
<position>43,-2022</position>
<input>
<ID>IN_0</ID>1473 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2610</ID>
<type>AE_DFF_LOW</type>
<position>82,-2015.5</position>
<output>
<ID>OUT_0</ID>1475 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2611</ID>
<type>AA_AND2</type>
<position>89.5,-2021</position>
<input>
<ID>IN_0</ID>1475 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2612</ID>
<type>AE_DFF_LOW</type>
<position>131.5,-2015.5</position>
<output>
<ID>OUT_0</ID>1476 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2613</ID>
<type>AA_AND2</type>
<position>140,-2021</position>
<input>
<ID>IN_0</ID>1476 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2614</ID>
<type>AE_DFF_LOW</type>
<position>179.5,-2015.5</position>
<output>
<ID>OUT_0</ID>1477 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2615</ID>
<type>AA_AND2</type>
<position>188,-2020.5</position>
<input>
<ID>IN_0</ID>1477 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2616</ID>
<type>AE_DFF_LOW</type>
<position>237,-2015.5</position>
<output>
<ID>OUT_0</ID>1478 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2617</ID>
<type>AA_AND2</type>
<position>246.5,-2022.5</position>
<input>
<ID>IN_0</ID>1478 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2618</ID>
<type>AE_DFF_LOW</type>
<position>292,-2015.5</position>
<output>
<ID>OUT_0</ID>1479 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2619</ID>
<type>AA_AND2</type>
<position>300,-2021.5</position>
<input>
<ID>IN_0</ID>1479 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2620</ID>
<type>AE_DFF_LOW</type>
<position>349,-2015.5</position>
<output>
<ID>OUT_0</ID>1480 </output>
<input>
<ID>clock</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2621</ID>
<type>AA_AND2</type>
<position>358.5,-2022</position>
<input>
<ID>IN_0</ID>1480 </input>
<input>
<ID>IN_1</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2622</ID>
<type>AA_AND2</type>
<position>-47,-2014.5</position>
<input>
<ID>IN_0</ID>1544 </input>
<output>
<ID>OUT</ID>1474 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2623</ID>
<type>AE_DFF_LOW</type>
<position>-15.5,-2028.5</position>
<output>
<ID>OUT_0</ID>1481 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2624</ID>
<type>AA_AND2</type>
<position>-5.5,-2034</position>
<input>
<ID>IN_0</ID>1481 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2625</ID>
<type>AE_DFF_LOW</type>
<position>34,-2028.5</position>
<output>
<ID>OUT_0</ID>1482 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2626</ID>
<type>AA_AND2</type>
<position>43,-2035</position>
<input>
<ID>IN_0</ID>1482 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2627</ID>
<type>AE_DFF_LOW</type>
<position>82,-2028.5</position>
<output>
<ID>OUT_0</ID>1484 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2628</ID>
<type>AA_AND2</type>
<position>89.5,-2034</position>
<input>
<ID>IN_0</ID>1484 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2629</ID>
<type>AE_DFF_LOW</type>
<position>131.5,-2028.5</position>
<output>
<ID>OUT_0</ID>1485 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2630</ID>
<type>AA_AND2</type>
<position>140,-2034</position>
<input>
<ID>IN_0</ID>1485 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2631</ID>
<type>AE_DFF_LOW</type>
<position>179.5,-2028.5</position>
<output>
<ID>OUT_0</ID>1486 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2632</ID>
<type>AA_AND2</type>
<position>188,-2033.5</position>
<input>
<ID>IN_0</ID>1486 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2633</ID>
<type>AE_DFF_LOW</type>
<position>237,-2028.5</position>
<output>
<ID>OUT_0</ID>1487 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2634</ID>
<type>AA_AND2</type>
<position>246.5,-2035.5</position>
<input>
<ID>IN_0</ID>1487 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2635</ID>
<type>AE_DFF_LOW</type>
<position>292,-2028.5</position>
<output>
<ID>OUT_0</ID>1488 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2636</ID>
<type>AA_AND2</type>
<position>300,-2034.5</position>
<input>
<ID>IN_0</ID>1488 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2637</ID>
<type>AE_DFF_LOW</type>
<position>349,-2028.5</position>
<output>
<ID>OUT_0</ID>1489 </output>
<input>
<ID>clock</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2638</ID>
<type>AA_AND2</type>
<position>358.5,-2035</position>
<input>
<ID>IN_0</ID>1489 </input>
<input>
<ID>IN_1</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2639</ID>
<type>AA_AND2</type>
<position>-47,-2027.5</position>
<input>
<ID>IN_0</ID>1545 </input>
<output>
<ID>OUT</ID>1483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2640</ID>
<type>AE_DFF_LOW</type>
<position>-15.5,-2043</position>
<output>
<ID>OUT_0</ID>1490 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2641</ID>
<type>AA_AND2</type>
<position>-5.5,-2048.5</position>
<input>
<ID>IN_0</ID>1490 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2642</ID>
<type>AE_DFF_LOW</type>
<position>34,-2043</position>
<output>
<ID>OUT_0</ID>1491 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2643</ID>
<type>AA_AND2</type>
<position>43,-2049.5</position>
<input>
<ID>IN_0</ID>1491 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2644</ID>
<type>AE_DFF_LOW</type>
<position>82,-2043</position>
<output>
<ID>OUT_0</ID>1493 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2645</ID>
<type>AA_AND2</type>
<position>89.5,-2048.5</position>
<input>
<ID>IN_0</ID>1493 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2646</ID>
<type>AE_DFF_LOW</type>
<position>131.5,-2043</position>
<output>
<ID>OUT_0</ID>1494 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2647</ID>
<type>AA_AND2</type>
<position>140,-2048.5</position>
<input>
<ID>IN_0</ID>1494 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2648</ID>
<type>AE_DFF_LOW</type>
<position>179.5,-2043</position>
<output>
<ID>OUT_0</ID>1495 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2649</ID>
<type>AA_AND2</type>
<position>188,-2048</position>
<input>
<ID>IN_0</ID>1495 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2650</ID>
<type>AE_DFF_LOW</type>
<position>237,-2043</position>
<output>
<ID>OUT_0</ID>1496 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2651</ID>
<type>AA_AND2</type>
<position>246.5,-2050</position>
<input>
<ID>IN_0</ID>1496 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2652</ID>
<type>AE_DFF_LOW</type>
<position>292,-2043</position>
<output>
<ID>OUT_0</ID>1497 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2653</ID>
<type>AA_AND2</type>
<position>300,-2049</position>
<input>
<ID>IN_0</ID>1497 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2654</ID>
<type>AE_DFF_LOW</type>
<position>349,-2043</position>
<output>
<ID>OUT_0</ID>1498 </output>
<input>
<ID>clock</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2655</ID>
<type>AA_AND2</type>
<position>358.5,-2049.5</position>
<input>
<ID>IN_0</ID>1498 </input>
<input>
<ID>IN_1</ID>1492 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2656</ID>
<type>AA_AND2</type>
<position>-47,-2042</position>
<input>
<ID>IN_0</ID>1546 </input>
<output>
<ID>OUT</ID>1492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2657</ID>
<type>AE_DFF_LOW</type>
<position>-16,-2055.5</position>
<output>
<ID>OUT_0</ID>1499 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2658</ID>
<type>AA_AND2</type>
<position>-6,-2061</position>
<input>
<ID>IN_0</ID>1499 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2659</ID>
<type>AE_DFF_LOW</type>
<position>33.5,-2055.5</position>
<output>
<ID>OUT_0</ID>1500 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2660</ID>
<type>AA_AND2</type>
<position>42.5,-2062</position>
<input>
<ID>IN_0</ID>1500 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2661</ID>
<type>AE_DFF_LOW</type>
<position>81.5,-2055.5</position>
<output>
<ID>OUT_0</ID>1502 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2662</ID>
<type>AA_AND2</type>
<position>89,-2061</position>
<input>
<ID>IN_0</ID>1502 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2663</ID>
<type>AE_DFF_LOW</type>
<position>131,-2055.5</position>
<output>
<ID>OUT_0</ID>1503 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2664</ID>
<type>AA_AND2</type>
<position>139.5,-2061</position>
<input>
<ID>IN_0</ID>1503 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2665</ID>
<type>AE_DFF_LOW</type>
<position>179,-2055.5</position>
<output>
<ID>OUT_0</ID>1504 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2666</ID>
<type>AA_AND2</type>
<position>187.5,-2060.5</position>
<input>
<ID>IN_0</ID>1504 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2667</ID>
<type>AE_DFF_LOW</type>
<position>236.5,-2055.5</position>
<output>
<ID>OUT_0</ID>1505 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2668</ID>
<type>AA_AND2</type>
<position>246,-2062.5</position>
<input>
<ID>IN_0</ID>1505 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2669</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-2055.5</position>
<output>
<ID>OUT_0</ID>1506 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2670</ID>
<type>AA_AND2</type>
<position>299.5,-2061.5</position>
<input>
<ID>IN_0</ID>1506 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2671</ID>
<type>AE_DFF_LOW</type>
<position>348.5,-2055.5</position>
<output>
<ID>OUT_0</ID>1507 </output>
<input>
<ID>clock</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2672</ID>
<type>AA_AND2</type>
<position>358,-2062</position>
<input>
<ID>IN_0</ID>1507 </input>
<input>
<ID>IN_1</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2673</ID>
<type>AA_AND2</type>
<position>-47.5,-2054.5</position>
<input>
<ID>IN_0</ID>1547 </input>
<output>
<ID>OUT</ID>1501 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2674</ID>
<type>AE_DFF_LOW</type>
<position>-16.5,-2068.5</position>
<output>
<ID>OUT_0</ID>1508 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2675</ID>
<type>AA_AND2</type>
<position>-6.5,-2074</position>
<input>
<ID>IN_0</ID>1508 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2676</ID>
<type>AE_DFF_LOW</type>
<position>33,-2068.5</position>
<output>
<ID>OUT_0</ID>1509 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2677</ID>
<type>AA_AND2</type>
<position>42,-2075</position>
<input>
<ID>IN_0</ID>1509 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2678</ID>
<type>AE_DFF_LOW</type>
<position>81,-2068.5</position>
<output>
<ID>OUT_0</ID>1511 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2679</ID>
<type>AA_AND2</type>
<position>88.5,-2074</position>
<input>
<ID>IN_0</ID>1511 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2680</ID>
<type>AE_DFF_LOW</type>
<position>130.5,-2068.5</position>
<output>
<ID>OUT_0</ID>1512 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2681</ID>
<type>AA_AND2</type>
<position>139,-2074</position>
<input>
<ID>IN_0</ID>1512 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2682</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-2068.5</position>
<output>
<ID>OUT_0</ID>1513 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2683</ID>
<type>AA_AND2</type>
<position>187,-2073.5</position>
<input>
<ID>IN_0</ID>1513 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2684</ID>
<type>AE_DFF_LOW</type>
<position>236,-2068.5</position>
<output>
<ID>OUT_0</ID>1514 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2685</ID>
<type>AA_AND2</type>
<position>245.5,-2075.5</position>
<input>
<ID>IN_0</ID>1514 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2686</ID>
<type>AE_DFF_LOW</type>
<position>291,-2068.5</position>
<output>
<ID>OUT_0</ID>1515 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2687</ID>
<type>AA_AND2</type>
<position>299,-2074.5</position>
<input>
<ID>IN_0</ID>1515 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2688</ID>
<type>AE_DFF_LOW</type>
<position>348,-2068.5</position>
<output>
<ID>OUT_0</ID>1516 </output>
<input>
<ID>clock</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2689</ID>
<type>AA_AND2</type>
<position>357.5,-2075</position>
<input>
<ID>IN_0</ID>1516 </input>
<input>
<ID>IN_1</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2690</ID>
<type>AA_AND2</type>
<position>-48,-2067.5</position>
<input>
<ID>IN_0</ID>1548 </input>
<output>
<ID>OUT</ID>1510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1152</ID>
<type>AA_TOGGLE</type>
<position>-268,-1329</position>
<output>
<ID>OUT_0</ID>671 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1153</ID>
<type>AA_TOGGLE</type>
<position>-268,-1325.5</position>
<output>
<ID>OUT_0</ID>674 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1154</ID>
<type>AA_TOGGLE</type>
<position>-268,-1322.5</position>
<output>
<ID>OUT_0</ID>673 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1156</ID>
<type>AA_LABEL</type>
<position>-260.5,-1320.5</position>
<gparam>LABEL_TEXT 3rd</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1158</ID>
<type>AA_LABEL</type>
<position>-260.5,-1323.5</position>
<gparam>LABEL_TEXT 2nd</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1160</ID>
<type>AA_LABEL</type>
<position>-261,-1327</position>
<gparam>LABEL_TEXT 1st</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1450</ID>
<type>AE_DFF_LOW</type>
<position>-25.5,-54</position>
<output>
<ID>OUT_0</ID>829 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1451</ID>
<type>AA_AND2</type>
<position>-15.5,-59.5</position>
<input>
<ID>IN_0</ID>829 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1452</ID>
<type>AE_DFF_LOW</type>
<position>24,-54</position>
<output>
<ID>OUT_0</ID>830 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1453</ID>
<type>AA_AND2</type>
<position>33,-60.5</position>
<input>
<ID>IN_0</ID>830 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1454</ID>
<type>AE_DFF_LOW</type>
<position>72,-54</position>
<output>
<ID>OUT_0</ID>832 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1455</ID>
<type>AA_AND2</type>
<position>79.5,-59.5</position>
<input>
<ID>IN_0</ID>832 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1456</ID>
<type>AE_DFF_LOW</type>
<position>121.5,-54</position>
<output>
<ID>OUT_0</ID>833 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1457</ID>
<type>AA_AND2</type>
<position>130,-59.5</position>
<input>
<ID>IN_0</ID>833 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1458</ID>
<type>AE_DFF_LOW</type>
<position>169.5,-54</position>
<output>
<ID>OUT_0</ID>834 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1459</ID>
<type>AA_AND2</type>
<position>178,-59</position>
<input>
<ID>IN_0</ID>834 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1460</ID>
<type>AE_DFF_LOW</type>
<position>227,-54</position>
<output>
<ID>OUT_0</ID>835 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1461</ID>
<type>AA_AND2</type>
<position>236.5,-61</position>
<input>
<ID>IN_0</ID>835 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1462</ID>
<type>AE_DFF_LOW</type>
<position>282,-54</position>
<output>
<ID>OUT_0</ID>836 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1463</ID>
<type>AA_AND2</type>
<position>290,-60</position>
<input>
<ID>IN_0</ID>836 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1464</ID>
<type>AE_DFF_LOW</type>
<position>339,-54</position>
<output>
<ID>OUT_0</ID>837 </output>
<input>
<ID>clock</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1465</ID>
<type>AA_AND2</type>
<position>348.5,-60.5</position>
<input>
<ID>IN_0</ID>837 </input>
<input>
<ID>IN_1</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1466</ID>
<type>AA_AND2</type>
<position>-57,-53</position>
<input>
<ID>IN_0</ID>838 </input>
<output>
<ID>OUT</ID>831 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1467</ID>
<type>AE_DFF_LOW</type>
<position>-25.5,-67</position>
<output>
<ID>OUT_0</ID>839 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1468</ID>
<type>AA_AND2</type>
<position>-15.5,-72.5</position>
<input>
<ID>IN_0</ID>839 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1469</ID>
<type>AE_DFF_LOW</type>
<position>24,-67</position>
<output>
<ID>OUT_0</ID>840 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1470</ID>
<type>AA_AND2</type>
<position>33,-73.5</position>
<input>
<ID>IN_0</ID>840 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1471</ID>
<type>AE_DFF_LOW</type>
<position>72,-67</position>
<output>
<ID>OUT_0</ID>842 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1472</ID>
<type>AA_AND2</type>
<position>79.5,-72.5</position>
<input>
<ID>IN_0</ID>842 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1473</ID>
<type>AE_DFF_LOW</type>
<position>121.5,-67</position>
<output>
<ID>OUT_0</ID>843 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1474</ID>
<type>AA_AND2</type>
<position>130,-72.5</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1475</ID>
<type>AE_DFF_LOW</type>
<position>169.5,-67</position>
<output>
<ID>OUT_0</ID>844 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1476</ID>
<type>AA_AND2</type>
<position>178,-72</position>
<input>
<ID>IN_0</ID>844 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1477</ID>
<type>AE_DFF_LOW</type>
<position>227,-67</position>
<output>
<ID>OUT_0</ID>845 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1478</ID>
<type>AA_AND2</type>
<position>236.5,-74</position>
<input>
<ID>IN_0</ID>845 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1479</ID>
<type>AE_DFF_LOW</type>
<position>282,-67</position>
<output>
<ID>OUT_0</ID>846 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1480</ID>
<type>AA_AND2</type>
<position>290,-73</position>
<input>
<ID>IN_0</ID>846 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1481</ID>
<type>AE_DFF_LOW</type>
<position>339,-67</position>
<output>
<ID>OUT_0</ID>847 </output>
<input>
<ID>clock</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1482</ID>
<type>AA_AND2</type>
<position>348.5,-73.5</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1483</ID>
<type>AA_AND2</type>
<position>-57,-66</position>
<input>
<ID>IN_0</ID>848 </input>
<output>
<ID>OUT</ID>841 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1484</ID>
<type>AE_DFF_LOW</type>
<position>-25.5,-81.5</position>
<output>
<ID>OUT_0</ID>849 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1485</ID>
<type>AA_AND2</type>
<position>-15.5,-87</position>
<input>
<ID>IN_0</ID>849 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1486</ID>
<type>AE_DFF_LOW</type>
<position>24,-81.5</position>
<output>
<ID>OUT_0</ID>850 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1487</ID>
<type>AA_AND2</type>
<position>33,-88</position>
<input>
<ID>IN_0</ID>850 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1488</ID>
<type>AE_DFF_LOW</type>
<position>72,-81.5</position>
<output>
<ID>OUT_0</ID>852 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1489</ID>
<type>AA_AND2</type>
<position>79.5,-87</position>
<input>
<ID>IN_0</ID>852 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1490</ID>
<type>AE_DFF_LOW</type>
<position>121.5,-81.5</position>
<output>
<ID>OUT_0</ID>853 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1491</ID>
<type>AA_AND2</type>
<position>130,-87</position>
<input>
<ID>IN_0</ID>853 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1492</ID>
<type>AE_DFF_LOW</type>
<position>169.5,-81.5</position>
<output>
<ID>OUT_0</ID>854 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1493</ID>
<type>AA_AND2</type>
<position>178,-86.5</position>
<input>
<ID>IN_0</ID>854 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1494</ID>
<type>AE_DFF_LOW</type>
<position>227,-81.5</position>
<output>
<ID>OUT_0</ID>855 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1495</ID>
<type>AA_AND2</type>
<position>236.5,-88.5</position>
<input>
<ID>IN_0</ID>855 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1496</ID>
<type>AE_DFF_LOW</type>
<position>282,-81.5</position>
<output>
<ID>OUT_0</ID>856 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1497</ID>
<type>AA_AND2</type>
<position>290,-87.5</position>
<input>
<ID>IN_0</ID>856 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1498</ID>
<type>AE_DFF_LOW</type>
<position>339,-81.5</position>
<output>
<ID>OUT_0</ID>857 </output>
<input>
<ID>clock</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1499</ID>
<type>AA_AND2</type>
<position>348.5,-88</position>
<input>
<ID>IN_0</ID>857 </input>
<input>
<ID>IN_1</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1500</ID>
<type>AA_AND2</type>
<position>-57,-80.5</position>
<input>
<ID>IN_0</ID>858 </input>
<output>
<ID>OUT</ID>851 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1501</ID>
<type>AE_DFF_LOW</type>
<position>-26,-94</position>
<output>
<ID>OUT_0</ID>859 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1502</ID>
<type>AA_AND2</type>
<position>-16,-99.5</position>
<input>
<ID>IN_0</ID>859 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1503</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-94</position>
<output>
<ID>OUT_0</ID>860 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1504</ID>
<type>AA_AND2</type>
<position>32.5,-100.5</position>
<input>
<ID>IN_0</ID>860 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1505</ID>
<type>AE_DFF_LOW</type>
<position>71.5,-94</position>
<output>
<ID>OUT_0</ID>862 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1506</ID>
<type>AA_AND2</type>
<position>79,-99.5</position>
<input>
<ID>IN_0</ID>862 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1507</ID>
<type>AE_DFF_LOW</type>
<position>121,-94</position>
<output>
<ID>OUT_0</ID>863 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1508</ID>
<type>AA_AND2</type>
<position>129.5,-99.5</position>
<input>
<ID>IN_0</ID>863 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1509</ID>
<type>AE_DFF_LOW</type>
<position>169,-94</position>
<output>
<ID>OUT_0</ID>864 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1510</ID>
<type>AA_AND2</type>
<position>177.5,-99</position>
<input>
<ID>IN_0</ID>864 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1511</ID>
<type>AE_DFF_LOW</type>
<position>226.5,-94</position>
<output>
<ID>OUT_0</ID>865 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1512</ID>
<type>AA_AND2</type>
<position>236,-101</position>
<input>
<ID>IN_0</ID>865 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1513</ID>
<type>AE_DFF_LOW</type>
<position>281.5,-94</position>
<output>
<ID>OUT_0</ID>866 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1514</ID>
<type>AA_AND2</type>
<position>289.5,-100</position>
<input>
<ID>IN_0</ID>866 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1515</ID>
<type>AE_DFF_LOW</type>
<position>338.5,-94</position>
<output>
<ID>OUT_0</ID>867 </output>
<input>
<ID>clock</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1516</ID>
<type>AA_AND2</type>
<position>348,-100.5</position>
<input>
<ID>IN_0</ID>867 </input>
<input>
<ID>IN_1</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1517</ID>
<type>AA_AND2</type>
<position>-57.5,-93</position>
<input>
<ID>IN_0</ID>868 </input>
<output>
<ID>OUT</ID>861 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1518</ID>
<type>AE_DFF_LOW</type>
<position>-26.5,-107</position>
<output>
<ID>OUT_0</ID>869 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1519</ID>
<type>AA_AND2</type>
<position>-16.5,-112.5</position>
<input>
<ID>IN_0</ID>869 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1520</ID>
<type>AE_DFF_LOW</type>
<position>23,-107</position>
<output>
<ID>OUT_0</ID>870 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1521</ID>
<type>AA_AND2</type>
<position>32,-113.5</position>
<input>
<ID>IN_0</ID>870 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1522</ID>
<type>AE_DFF_LOW</type>
<position>71,-107</position>
<output>
<ID>OUT_0</ID>872 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1523</ID>
<type>AA_AND2</type>
<position>78.5,-112.5</position>
<input>
<ID>IN_0</ID>872 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1524</ID>
<type>AE_DFF_LOW</type>
<position>120.5,-107</position>
<output>
<ID>OUT_0</ID>873 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1525</ID>
<type>AA_AND2</type>
<position>129,-112.5</position>
<input>
<ID>IN_0</ID>873 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1526</ID>
<type>AE_DFF_LOW</type>
<position>168.5,-107</position>
<output>
<ID>OUT_0</ID>874 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1527</ID>
<type>AA_AND2</type>
<position>177,-112</position>
<input>
<ID>IN_0</ID>874 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1528</ID>
<type>AE_DFF_LOW</type>
<position>226,-107</position>
<output>
<ID>OUT_0</ID>875 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1529</ID>
<type>AA_AND2</type>
<position>235.5,-114</position>
<input>
<ID>IN_0</ID>875 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1530</ID>
<type>AE_DFF_LOW</type>
<position>281,-107</position>
<output>
<ID>OUT_0</ID>876 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1531</ID>
<type>AA_AND2</type>
<position>289,-113</position>
<input>
<ID>IN_0</ID>876 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1532</ID>
<type>AE_DFF_LOW</type>
<position>338,-107</position>
<output>
<ID>OUT_0</ID>877 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1533</ID>
<type>AA_AND2</type>
<position>347.5,-113.5</position>
<input>
<ID>IN_0</ID>877 </input>
<input>
<ID>IN_1</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1534</ID>
<type>AA_AND2</type>
<position>-58,-106</position>
<input>
<ID>IN_0</ID>878 </input>
<output>
<ID>OUT</ID>871 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-2119.5,85,-2113</points>
<connection>
<GID>2594</GID>
<name>IN_0</name></connection>
<intersection>-2113 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83.5,-2113,85,-2113</points>
<connection>
<GID>2593</GID>
<name>OUT_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>1539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-2119.5,134.5,-2113</points>
<intersection>-2119.5 1</intersection>
<intersection>-2113 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,-2119.5,135.5,-2119.5</points>
<connection>
<GID>2596</GID>
<name>IN_0</name></connection>
<intersection>134.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133,-2113,134.5,-2113</points>
<connection>
<GID>2595</GID>
<name>OUT_0</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-170,-1333.5,-170,-79</points>
<intersection>-1333.5 1</intersection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1333.5,-170,-1333.5</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<intersection>-170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-170,-79,-88,-79</points>
<intersection>-170 0</intersection>
<intersection>-88 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-88,-84.5,-88,-79</points>
<connection>
<GID>57</GID>
<name>ENABLE</name></connection>
<intersection>-79 2</intersection></vsegment></shape></wire>
<wire>
<ID>1540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-2119,183,-2113</points>
<intersection>-2119 5</intersection>
<intersection>-2113 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>181,-2113,183,-2113</points>
<connection>
<GID>2597</GID>
<name>OUT_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>183,-2119,183.5,-2119</points>
<connection>
<GID>2598</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-169,-1334.5,-169,-323</points>
<intersection>-1334.5 1</intersection>
<intersection>-323 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1334.5,-169,-1334.5</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>-169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-169,-323,-84.5,-323</points>
<connection>
<GID>195</GID>
<name>ENABLE</name></connection>
<intersection>-169 0</intersection></hsegment></shape></wire>
<wire>
<ID>1541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-2121,241.5,-2113</points>
<intersection>-2121 1</intersection>
<intersection>-2113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241.5,-2121,242,-2121</points>
<connection>
<GID>2600</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-2113,241.5,-2113</points>
<connection>
<GID>2599</GID>
<name>OUT_0</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-168,-1335.5,-168,-618</points>
<intersection>-1335.5 1</intersection>
<intersection>-618 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1335.5,-168,-1335.5</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>-168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-168,-618,-92,-618</points>
<connection>
<GID>332</GID>
<name>ENABLE</name></connection>
<intersection>-168 0</intersection></hsegment></shape></wire>
<wire>
<ID>1542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-2120,295,-2113</points>
<intersection>-2120 4</intersection>
<intersection>-2113 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293.5,-2113,295,-2113</points>
<connection>
<GID>2601</GID>
<name>OUT_0</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>295,-2120,295.5,-2120</points>
<connection>
<GID>2602</GID>
<name>IN_0</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-1336.5,-167,-917</points>
<intersection>-1336.5 1</intersection>
<intersection>-917 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1336.5,-167,-1336.5</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>-167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-167,-917,-85,-917</points>
<connection>
<GID>469</GID>
<name>ENABLE</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>1543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353.5,-2120.5,353.5,-2113</points>
<intersection>-2120.5 1</intersection>
<intersection>-2113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353.5,-2120.5,354,-2120.5</points>
<connection>
<GID>2604</GID>
<name>IN_0</name></connection>
<intersection>353.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350.5,-2113,353.5,-2113</points>
<connection>
<GID>2603</GID>
<name>OUT_0</name></connection>
<intersection>353.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-166,-1337.5,-166,-1234.5</points>
<intersection>-1337.5 1</intersection>
<intersection>-1234.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1337.5,-166,-1337.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>-166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-166,-1234.5,-92,-1234.5</points>
<connection>
<GID>606</GID>
<name>ENABLE</name></connection>
<intersection>-166 0</intersection></hsegment></shape></wire>
<wire>
<ID>1544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-2063.5,-69.5,-2013.5</points>
<intersection>-2063.5 2</intersection>
<intersection>-2013.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-2013.5,-50,-2013.5</points>
<connection>
<GID>2622</GID>
<name>IN_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2063.5,-69.5,-2063.5</points>
<connection>
<GID>1017</GID>
<name>OUT_7</name></connection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-2064.5,-68.5,-2026.5</points>
<intersection>-2064.5 2</intersection>
<intersection>-2026.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,-2026.5,-50,-2026.5</points>
<connection>
<GID>2639</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2064.5,-68.5,-2064.5</points>
<connection>
<GID>1017</GID>
<name>OUT_6</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-2065.5,-67.5,-2041</points>
<intersection>-2065.5 2</intersection>
<intersection>-2041 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-2041,-50,-2041</points>
<connection>
<GID>2656</GID>
<name>IN_0</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2065.5,-67.5,-2065.5</points>
<connection>
<GID>1017</GID>
<name>OUT_5</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-2066.5,-66.5,-2053.5</points>
<intersection>-2066.5 2</intersection>
<intersection>-2053.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,-2053.5,-50.5,-2053.5</points>
<connection>
<GID>2673</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2066.5,-66.5,-2066.5</points>
<connection>
<GID>1017</GID>
<name>OUT_4</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83.5,-2067.5,-66,-2067.5</points>
<connection>
<GID>1017</GID>
<name>OUT_3</name></connection>
<intersection>-66 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-66,-2067.5,-66,-2066.5</points>
<intersection>-2067.5 1</intersection>
<intersection>-2066.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-66,-2066.5,-51,-2066.5</points>
<connection>
<GID>2690</GID>
<name>IN_0</name></connection>
<intersection>-66 5</intersection></hsegment></shape></wire>
<wire>
<ID>1549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-2081.5,-67,-2068.5</points>
<intersection>-2081.5 1</intersection>
<intersection>-2068.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,-2081.5,-51,-2081.5</points>
<connection>
<GID>2571</GID>
<name>IN_0</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2068.5,-67,-2068.5</points>
<connection>
<GID>1017</GID>
<name>OUT_2</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>1550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,-2095.5,-68,-2069.5</points>
<intersection>-2095.5 1</intersection>
<intersection>-2069.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-2095.5,-51,-2095.5</points>
<connection>
<GID>2588</GID>
<name>IN_0</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2069.5,-68,-2069.5</points>
<connection>
<GID>1017</GID>
<name>OUT_1</name></connection>
<intersection>-68 0</intersection></hsegment></shape></wire>
<wire>
<ID>1551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-2113,-69,-2070.5</points>
<intersection>-2113 1</intersection>
<intersection>-2070.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-2113,-51.5,-2113</points>
<connection>
<GID>2605</GID>
<name>IN_0</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-2070.5,-69,-2070.5</points>
<connection>
<GID>1017</GID>
<name>OUT_0</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>1553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-166,-1471,-166,-1338.5</points>
<intersection>-1471 2</intersection>
<intersection>-1338.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1338.5,-166,-1338.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>-166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-166,-1471,-88.5,-1471</points>
<connection>
<GID>743</GID>
<name>ENABLE</name></connection>
<intersection>-166 0</intersection></hsegment></shape></wire>
<wire>
<ID>1554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-1765.5,-167,-1339.5</points>
<intersection>-1765.5 2</intersection>
<intersection>-1339.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1339.5,-167,-1339.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>-167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-167,-1765.5,-92.5,-1765.5</points>
<connection>
<GID>880</GID>
<name>ENABLE</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>1555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-168,-2063.5,-168,-1340.5</points>
<intersection>-2063.5 2</intersection>
<intersection>-1340.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-263.5,-1340.5,-168,-1340.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-168,-2063.5,-89.5,-2063.5</points>
<connection>
<GID>1017</GID>
<name>ENABLE</name></connection>
<intersection>-168 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,-975.5,-54,-961.5</points>
<intersection>-975.5 2</intersection>
<intersection>-961.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-961.5,-49,-961.5</points>
<connection>
<GID>1925</GID>
<name>IN_1</name></connection>
<intersection>-54 0</intersection>
<intersection>-49 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-58.5,-975.5,-54,-975.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-54 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-49,-961.5,-49,-944</points>
<connection>
<GID>1908</GID>
<name>IN_1</name></connection>
<intersection>-961.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-58.5,-21,-52</points>
<intersection>-58.5 1</intersection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-58.5,-18.5,-58.5</points>
<connection>
<GID>1451</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-22.5,-52,-21,-52</points>
<connection>
<GID>1450</GID>
<name>OUT_0</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-59.5,28,-52</points>
<intersection>-59.5 1</intersection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-59.5,30,-59.5</points>
<connection>
<GID>1453</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-52,28,-52</points>
<connection>
<GID>1452</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-53,345.5,-53</points>
<connection>
<GID>1466</GID>
<name>OUT</name></connection>
<intersection>-28.5 107</intersection>
<intersection>-20 4</intersection>
<intersection>21 108</intersection>
<intersection>28.5 16</intersection>
<intersection>69 109</intersection>
<intersection>76 23</intersection>
<intersection>118.5 110</intersection>
<intersection>126.5 31</intersection>
<intersection>166.5 111</intersection>
<intersection>175 55</intersection>
<intersection>224 112</intersection>
<intersection>233.5 56</intersection>
<intersection>279 113</intersection>
<intersection>287.5 66</intersection>
<intersection>336 114</intersection>
<intersection>345.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-20,-60.5,-20,-53</points>
<intersection>-60.5 5</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-20,-60.5,-18.5,-60.5</points>
<connection>
<GID>1451</GID>
<name>IN_1</name></connection>
<intersection>-20 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>28.5,-61.5,28.5,-53</points>
<intersection>-61.5 21</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>28.5,-61.5,30,-61.5</points>
<connection>
<GID>1453</GID>
<name>IN_1</name></connection>
<intersection>28.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>76,-60.5,76,-53</points>
<intersection>-60.5 53</intersection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>126.5,-60.5,126.5,-53</points>
<intersection>-60.5 115</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>76,-60.5,76.5,-60.5</points>
<connection>
<GID>1455</GID>
<name>IN_1</name></connection>
<intersection>76 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>175,-60,175,-53</points>
<connection>
<GID>1459</GID>
<name>IN_1</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>233.5,-62,233.5,-53</points>
<connection>
<GID>1461</GID>
<name>IN_1</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>287.5,-61,287.5,-53</points>
<intersection>-61 118</intersection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>345.5,-61.5,345.5,-53</points>
<connection>
<GID>1465</GID>
<name>IN_1</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-28.5,-55,-28.5,-53</points>
<connection>
<GID>1450</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>21,-55,21,-53</points>
<connection>
<GID>1452</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>69,-55,69,-53</points>
<connection>
<GID>1454</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>118.5,-55,118.5,-53</points>
<connection>
<GID>1456</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>166.5,-55,166.5,-53</points>
<connection>
<GID>1458</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>224,-55,224,-53</points>
<connection>
<GID>1460</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>279,-55,279,-53</points>
<connection>
<GID>1462</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>336,-55,336,-53</points>
<connection>
<GID>1464</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>126.5,-60.5,127,-60.5</points>
<connection>
<GID>1457</GID>
<name>IN_1</name></connection>
<intersection>126.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>287,-61,287.5,-61</points>
<connection>
<GID>1463</GID>
<name>IN_1</name></connection>
<intersection>287.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-58.5,76.5,-52</points>
<connection>
<GID>1455</GID>
<name>IN_0</name></connection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-52,76.5,-52</points>
<connection>
<GID>1454</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>833</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-58.5,126,-52</points>
<intersection>-58.5 1</intersection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-58.5,127,-58.5</points>
<connection>
<GID>1457</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>124.5,-52,126,-52</points>
<connection>
<GID>1456</GID>
<name>OUT_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>834</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-58,174.5,-52</points>
<intersection>-58 5</intersection>
<intersection>-52 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172.5,-52,174.5,-52</points>
<connection>
<GID>1458</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>174.5,-58,175,-58</points>
<connection>
<GID>1459</GID>
<name>IN_0</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-60,233,-52</points>
<intersection>-60 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,-60,233.5,-60</points>
<connection>
<GID>1461</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230,-52,233,-52</points>
<connection>
<GID>1460</GID>
<name>OUT_0</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>836</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-59,286.5,-52</points>
<intersection>-59 4</intersection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>285,-52,286.5,-52</points>
<connection>
<GID>1462</GID>
<name>OUT_0</name></connection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>286.5,-59,287,-59</points>
<connection>
<GID>1463</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345,-59.5,345,-52</points>
<intersection>-59.5 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345,-59.5,345.5,-59.5</points>
<connection>
<GID>1465</GID>
<name>IN_0</name></connection>
<intersection>345 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,-52,345,-52</points>
<connection>
<GID>1464</GID>
<name>OUT_0</name></connection>
<intersection>345 0</intersection></hsegment></shape></wire>
<wire>
<ID>838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-84.5,-65,-52</points>
<intersection>-84.5 2</intersection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-52,-60,-52</points>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-84.5,-65,-84.5</points>
<connection>
<GID>57</GID>
<name>OUT_7</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-71.5,-21,-65</points>
<intersection>-71.5 1</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-71.5,-18.5,-71.5</points>
<connection>
<GID>1468</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-22.5,-65,-21,-65</points>
<connection>
<GID>1467</GID>
<name>OUT_0</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-72.5,28,-65</points>
<intersection>-72.5 1</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-72.5,30,-72.5</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-65,28,-65</points>
<connection>
<GID>1469</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>841</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-66,345.5,-66</points>
<connection>
<GID>1483</GID>
<name>OUT</name></connection>
<intersection>-28.5 107</intersection>
<intersection>-20 4</intersection>
<intersection>21 108</intersection>
<intersection>28.5 16</intersection>
<intersection>69 109</intersection>
<intersection>76 23</intersection>
<intersection>118.5 110</intersection>
<intersection>126.5 31</intersection>
<intersection>166.5 111</intersection>
<intersection>175 55</intersection>
<intersection>224 112</intersection>
<intersection>233.5 56</intersection>
<intersection>279 113</intersection>
<intersection>287.5 66</intersection>
<intersection>336 114</intersection>
<intersection>345.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-20,-73.5,-20,-66</points>
<intersection>-73.5 5</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-20,-73.5,-18.5,-73.5</points>
<connection>
<GID>1468</GID>
<name>IN_1</name></connection>
<intersection>-20 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>28.5,-74.5,28.5,-66</points>
<intersection>-74.5 21</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>28.5,-74.5,30,-74.5</points>
<connection>
<GID>1470</GID>
<name>IN_1</name></connection>
<intersection>28.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>76,-73.5,76,-66</points>
<intersection>-73.5 53</intersection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>126.5,-73.5,126.5,-66</points>
<intersection>-73.5 115</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>76,-73.5,76.5,-73.5</points>
<connection>
<GID>1472</GID>
<name>IN_1</name></connection>
<intersection>76 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>175,-73,175,-66</points>
<connection>
<GID>1476</GID>
<name>IN_1</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>233.5,-75,233.5,-66</points>
<connection>
<GID>1478</GID>
<name>IN_1</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>287.5,-74,287.5,-66</points>
<intersection>-74 118</intersection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>345.5,-74.5,345.5,-66</points>
<connection>
<GID>1482</GID>
<name>IN_1</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-28.5,-68,-28.5,-66</points>
<connection>
<GID>1467</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>21,-68,21,-66</points>
<connection>
<GID>1469</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>69,-68,69,-66</points>
<connection>
<GID>1471</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>118.5,-68,118.5,-66</points>
<connection>
<GID>1473</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>166.5,-68,166.5,-66</points>
<connection>
<GID>1475</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>224,-68,224,-66</points>
<connection>
<GID>1477</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>279,-68,279,-66</points>
<connection>
<GID>1479</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>336,-68,336,-66</points>
<connection>
<GID>1481</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>126.5,-73.5,127,-73.5</points>
<connection>
<GID>1474</GID>
<name>IN_1</name></connection>
<intersection>126.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>287,-74,287.5,-74</points>
<connection>
<GID>1480</GID>
<name>IN_1</name></connection>
<intersection>287.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-71.5,76.5,-65</points>
<connection>
<GID>1472</GID>
<name>IN_0</name></connection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-65,76.5,-65</points>
<connection>
<GID>1471</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>843</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-71.5,126,-65</points>
<intersection>-71.5 1</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-71.5,127,-71.5</points>
<connection>
<GID>1474</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>124.5,-65,126,-65</points>
<connection>
<GID>1473</GID>
<name>OUT_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-71,174.5,-65</points>
<intersection>-71 5</intersection>
<intersection>-65 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172.5,-65,174.5,-65</points>
<connection>
<GID>1475</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>174.5,-71,175,-71</points>
<connection>
<GID>1476</GID>
<name>IN_0</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-73,233,-65</points>
<intersection>-73 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,-73,233.5,-73</points>
<connection>
<GID>1478</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230,-65,233,-65</points>
<connection>
<GID>1477</GID>
<name>OUT_0</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>846</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-72,286.5,-65</points>
<intersection>-72 4</intersection>
<intersection>-65 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>285,-65,286.5,-65</points>
<connection>
<GID>1479</GID>
<name>OUT_0</name></connection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>286.5,-72,287,-72</points>
<connection>
<GID>1480</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345,-72.5,345,-65</points>
<intersection>-72.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345,-72.5,345.5,-72.5</points>
<connection>
<GID>1482</GID>
<name>IN_0</name></connection>
<intersection>345 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,-65,345,-65</points>
<connection>
<GID>1481</GID>
<name>OUT_0</name></connection>
<intersection>345 0</intersection></hsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,-85.5,-64,-65</points>
<intersection>-85.5 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-65,-60,-65</points>
<connection>
<GID>1483</GID>
<name>IN_0</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-85.5,-64,-85.5</points>
<connection>
<GID>57</GID>
<name>OUT_6</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-86,-21,-79.5</points>
<intersection>-86 1</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-86,-18.5,-86</points>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-22.5,-79.5,-21,-79.5</points>
<connection>
<GID>1484</GID>
<name>OUT_0</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>850</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-87,28,-79.5</points>
<intersection>-87 1</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-87,30,-87</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-79.5,28,-79.5</points>
<connection>
<GID>1486</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-80.5,345.5,-80.5</points>
<connection>
<GID>1500</GID>
<name>OUT</name></connection>
<intersection>-28.5 107</intersection>
<intersection>-20 4</intersection>
<intersection>21 108</intersection>
<intersection>28.5 16</intersection>
<intersection>69 109</intersection>
<intersection>76 23</intersection>
<intersection>118.5 110</intersection>
<intersection>126.5 31</intersection>
<intersection>166.5 111</intersection>
<intersection>175 55</intersection>
<intersection>224 112</intersection>
<intersection>233.5 56</intersection>
<intersection>279 113</intersection>
<intersection>287.5 66</intersection>
<intersection>336 114</intersection>
<intersection>345.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-20,-88,-20,-80.5</points>
<intersection>-88 5</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-20,-88,-18.5,-88</points>
<connection>
<GID>1485</GID>
<name>IN_1</name></connection>
<intersection>-20 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>28.5,-89,28.5,-80.5</points>
<intersection>-89 21</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>28.5,-89,30,-89</points>
<connection>
<GID>1487</GID>
<name>IN_1</name></connection>
<intersection>28.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>76,-88,76,-80.5</points>
<intersection>-88 53</intersection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>126.5,-88,126.5,-80.5</points>
<intersection>-88 115</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>76,-88,76.5,-88</points>
<connection>
<GID>1489</GID>
<name>IN_1</name></connection>
<intersection>76 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>175,-87.5,175,-80.5</points>
<connection>
<GID>1493</GID>
<name>IN_1</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>233.5,-89.5,233.5,-80.5</points>
<connection>
<GID>1495</GID>
<name>IN_1</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>287.5,-88.5,287.5,-80.5</points>
<intersection>-88.5 118</intersection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>345.5,-89,345.5,-80.5</points>
<connection>
<GID>1499</GID>
<name>IN_1</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-28.5,-82.5,-28.5,-80.5</points>
<connection>
<GID>1484</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>21,-82.5,21,-80.5</points>
<connection>
<GID>1486</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>69,-82.5,69,-80.5</points>
<connection>
<GID>1488</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>118.5,-82.5,118.5,-80.5</points>
<connection>
<GID>1490</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>166.5,-82.5,166.5,-80.5</points>
<connection>
<GID>1492</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>224,-82.5,224,-80.5</points>
<connection>
<GID>1494</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>279,-82.5,279,-80.5</points>
<connection>
<GID>1496</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>336,-82.5,336,-80.5</points>
<connection>
<GID>1498</GID>
<name>clock</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>126.5,-88,127,-88</points>
<connection>
<GID>1491</GID>
<name>IN_1</name></connection>
<intersection>126.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>287,-88.5,287.5,-88.5</points>
<connection>
<GID>1497</GID>
<name>IN_1</name></connection>
<intersection>287.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-86,76.5,-79.5</points>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-79.5,76.5,-79.5</points>
<connection>
<GID>1488</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>853</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-86,126,-79.5</points>
<intersection>-86 1</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-86,127,-86</points>
<connection>
<GID>1491</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>124.5,-79.5,126,-79.5</points>
<connection>
<GID>1490</GID>
<name>OUT_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-85.5,174.5,-79.5</points>
<intersection>-85.5 5</intersection>
<intersection>-79.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172.5,-79.5,174.5,-79.5</points>
<connection>
<GID>1492</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>174.5,-85.5,175,-85.5</points>
<connection>
<GID>1493</GID>
<name>IN_0</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>855</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-87.5,233,-79.5</points>
<intersection>-87.5 1</intersection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233,-87.5,233.5,-87.5</points>
<connection>
<GID>1495</GID>
<name>IN_0</name></connection>
<intersection>233 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230,-79.5,233,-79.5</points>
<connection>
<GID>1494</GID>
<name>OUT_0</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-86.5,286.5,-79.5</points>
<intersection>-86.5 4</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>285,-79.5,286.5,-79.5</points>
<connection>
<GID>1496</GID>
<name>OUT_0</name></connection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>286.5,-86.5,287,-86.5</points>
<connection>
<GID>1497</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345,-87,345,-79.5</points>
<intersection>-87 1</intersection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345,-87,345.5,-87</points>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<intersection>345 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,-79.5,345,-79.5</points>
<connection>
<GID>1498</GID>
<name>OUT_0</name></connection>
<intersection>345 0</intersection></hsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-86.5,-63,-79.5</points>
<intersection>-86.5 2</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-79.5,-60,-79.5</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-86.5,-63,-86.5</points>
<connection>
<GID>57</GID>
<name>OUT_5</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21.5,-98.5,-21.5,-92</points>
<intersection>-98.5 1</intersection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21.5,-98.5,-19,-98.5</points>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<intersection>-21.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-23,-92,-21.5,-92</points>
<connection>
<GID>1501</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-99.5,27.5,-92</points>
<intersection>-99.5 1</intersection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-99.5,29.5,-99.5</points>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-92,27.5,-92</points>
<connection>
<GID>1503</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54.5,-93,345,-93</points>
<connection>
<GID>1517</GID>
<name>OUT</name></connection>
<intersection>-29 107</intersection>
<intersection>-20.5 4</intersection>
<intersection>20.5 108</intersection>
<intersection>28 16</intersection>
<intersection>68.5 109</intersection>
<intersection>75.5 23</intersection>
<intersection>118 110</intersection>
<intersection>126 31</intersection>
<intersection>166 111</intersection>
<intersection>174.5 55</intersection>
<intersection>223.5 112</intersection>
<intersection>233 56</intersection>
<intersection>278.5 113</intersection>
<intersection>287 66</intersection>
<intersection>335.5 114</intersection>
<intersection>345 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-20.5,-100.5,-20.5,-93</points>
<intersection>-100.5 5</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-20.5,-100.5,-19,-100.5</points>
<connection>
<GID>1502</GID>
<name>IN_1</name></connection>
<intersection>-20.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>28,-101.5,28,-93</points>
<intersection>-101.5 21</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>28,-101.5,29.5,-101.5</points>
<connection>
<GID>1504</GID>
<name>IN_1</name></connection>
<intersection>28 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>75.5,-100.5,75.5,-93</points>
<intersection>-100.5 53</intersection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>126,-100.5,126,-93</points>
<intersection>-100.5 115</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>75.5,-100.5,76,-100.5</points>
<connection>
<GID>1506</GID>
<name>IN_1</name></connection>
<intersection>75.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>174.5,-100,174.5,-93</points>
<connection>
<GID>1510</GID>
<name>IN_1</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>233,-102,233,-93</points>
<connection>
<GID>1512</GID>
<name>IN_1</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>287,-101,287,-93</points>
<intersection>-101 118</intersection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>345,-101.5,345,-93</points>
<connection>
<GID>1516</GID>
<name>IN_1</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-29,-95,-29,-93</points>
<connection>
<GID>1501</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>20.5,-95,20.5,-93</points>
<connection>
<GID>1503</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>68.5,-95,68.5,-93</points>
<connection>
<GID>1505</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>118,-95,118,-93</points>
<connection>
<GID>1507</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>166,-95,166,-93</points>
<connection>
<GID>1509</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>223.5,-95,223.5,-93</points>
<connection>
<GID>1511</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>278.5,-95,278.5,-93</points>
<connection>
<GID>1513</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>335.5,-95,335.5,-93</points>
<connection>
<GID>1515</GID>
<name>clock</name></connection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>126,-100.5,126.5,-100.5</points>
<connection>
<GID>1508</GID>
<name>IN_1</name></connection>
<intersection>126 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>286.5,-101,287,-101</points>
<connection>
<GID>1514</GID>
<name>IN_1</name></connection>
<intersection>287 66</intersection></hsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-98.5,76,-92</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-92,76,-92</points>
<connection>
<GID>1505</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>863</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-98.5,125.5,-92</points>
<intersection>-98.5 1</intersection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-98.5,126.5,-98.5</points>
<connection>
<GID>1508</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>124,-92,125.5,-92</points>
<connection>
<GID>1507</GID>
<name>OUT_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>864</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-98,174,-92</points>
<intersection>-98 5</intersection>
<intersection>-92 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172,-92,174,-92</points>
<connection>
<GID>1509</GID>
<name>OUT_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>174,-98,174.5,-98</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>865</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-100,232.5,-92</points>
<intersection>-100 1</intersection>
<intersection>-92 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,-100,233,-100</points>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229.5,-92,232.5,-92</points>
<connection>
<GID>1511</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>866</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-99,286,-92</points>
<intersection>-99 4</intersection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>284.5,-92,286,-92</points>
<connection>
<GID>1513</GID>
<name>OUT_0</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>286,-99,286.5,-99</points>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>286 0</intersection></hsegment></shape></wire>
<wire>
<ID>867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,-99.5,344.5,-92</points>
<intersection>-99.5 1</intersection>
<intersection>-92 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,-99.5,345,-99.5</points>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-92,344.5,-92</points>
<connection>
<GID>1515</GID>
<name>OUT_0</name></connection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-92,-63,-87.5</points>
<intersection>-92 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-92,-60.5,-92</points>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-87.5,-63,-87.5</points>
<connection>
<GID>57</GID>
<name>OUT_4</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>869</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-111.5,-22,-105</points>
<intersection>-111.5 1</intersection>
<intersection>-105 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-111.5,-19.5,-111.5</points>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-23.5,-105,-22,-105</points>
<connection>
<GID>1518</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-112.5,27,-105</points>
<intersection>-112.5 1</intersection>
<intersection>-105 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-112.5,29,-112.5</points>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-105,27,-105</points>
<connection>
<GID>1520</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,-106,344.5,-106</points>
<connection>
<GID>1534</GID>
<name>OUT</name></connection>
<intersection>-29.5 107</intersection>
<intersection>-21 4</intersection>
<intersection>20 108</intersection>
<intersection>27.5 16</intersection>
<intersection>68 109</intersection>
<intersection>75 23</intersection>
<intersection>117.5 110</intersection>
<intersection>125.5 31</intersection>
<intersection>165.5 111</intersection>
<intersection>174 55</intersection>
<intersection>223 112</intersection>
<intersection>232.5 56</intersection>
<intersection>278 113</intersection>
<intersection>286.5 66</intersection>
<intersection>335 114</intersection>
<intersection>344.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-21,-113.5,-21,-106</points>
<intersection>-113.5 5</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-21,-113.5,-19.5,-113.5</points>
<connection>
<GID>1519</GID>
<name>IN_1</name></connection>
<intersection>-21 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>27.5,-114.5,27.5,-106</points>
<intersection>-114.5 21</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>27.5,-114.5,29,-114.5</points>
<connection>
<GID>1521</GID>
<name>IN_1</name></connection>
<intersection>27.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>75,-113.5,75,-106</points>
<intersection>-113.5 53</intersection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>125.5,-113.5,125.5,-106</points>
<intersection>-113.5 115</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>75,-113.5,75.5,-113.5</points>
<connection>
<GID>1523</GID>
<name>IN_1</name></connection>
<intersection>75 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>174,-113,174,-106</points>
<connection>
<GID>1527</GID>
<name>IN_1</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>232.5,-115,232.5,-106</points>
<connection>
<GID>1529</GID>
<name>IN_1</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>286.5,-114,286.5,-106</points>
<intersection>-114 118</intersection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>344.5,-114.5,344.5,-106</points>
<connection>
<GID>1533</GID>
<name>IN_1</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-29.5,-108,-29.5,-106</points>
<connection>
<GID>1518</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>20,-108,20,-106</points>
<connection>
<GID>1520</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>68,-108,68,-106</points>
<connection>
<GID>1522</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>117.5,-108,117.5,-106</points>
<connection>
<GID>1524</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>165.5,-108,165.5,-106</points>
<connection>
<GID>1526</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>223,-108,223,-106</points>
<connection>
<GID>1528</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>278,-108,278,-106</points>
<connection>
<GID>1530</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>335,-108,335,-106</points>
<connection>
<GID>1532</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>125.5,-113.5,126,-113.5</points>
<connection>
<GID>1525</GID>
<name>IN_1</name></connection>
<intersection>125.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>286,-114,286.5,-114</points>
<connection>
<GID>1531</GID>
<name>IN_1</name></connection>
<intersection>286.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-111.5,75.5,-105</points>
<connection>
<GID>1523</GID>
<name>IN_0</name></connection>
<intersection>-105 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-105,75.5,-105</points>
<connection>
<GID>1522</GID>
<name>OUT_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-111.5,125,-105</points>
<intersection>-111.5 1</intersection>
<intersection>-105 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-111.5,126,-111.5</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123.5,-105,125,-105</points>
<connection>
<GID>1524</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-111,173.5,-105</points>
<intersection>-111 5</intersection>
<intersection>-105 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>171.5,-105,173.5,-105</points>
<connection>
<GID>1526</GID>
<name>OUT_0</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>173.5,-111,174,-111</points>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-113,232,-105</points>
<intersection>-113 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232,-113,232.5,-113</points>
<connection>
<GID>1529</GID>
<name>IN_0</name></connection>
<intersection>232 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,-105,232,-105</points>
<connection>
<GID>1528</GID>
<name>OUT_0</name></connection>
<intersection>232 0</intersection></hsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-112,285.5,-105</points>
<intersection>-112 4</intersection>
<intersection>-105 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>284,-105,285.5,-105</points>
<connection>
<GID>1530</GID>
<name>OUT_0</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>285.5,-112,286,-112</points>
<connection>
<GID>1531</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,-112.5,344,-105</points>
<intersection>-112.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,-112.5,344.5,-112.5</points>
<connection>
<GID>1533</GID>
<name>IN_0</name></connection>
<intersection>344 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341,-105,344,-105</points>
<connection>
<GID>1532</GID>
<name>OUT_0</name></connection>
<intersection>344 0</intersection></hsegment></shape></wire>
<wire>
<ID>878</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-105,-64.5,-88.5</points>
<intersection>-105 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-105,-61,-105</points>
<connection>
<GID>1534</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-88.5,-64.5,-88.5</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>888</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-126.5,-22,-120</points>
<intersection>-126.5 1</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-126.5,-19.5,-126.5</points>
<connection>
<GID>1553</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-23.5,-120,-22,-120</points>
<connection>
<GID>1552</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>889</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-127.5,27,-120</points>
<intersection>-127.5 1</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-127.5,29,-127.5</points>
<connection>
<GID>1555</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-120,27,-120</points>
<connection>
<GID>1554</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>890</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,-121,344.5,-121</points>
<connection>
<GID>1568</GID>
<name>OUT</name></connection>
<intersection>-29.5 107</intersection>
<intersection>-21 4</intersection>
<intersection>20 108</intersection>
<intersection>27.5 16</intersection>
<intersection>68 109</intersection>
<intersection>75 23</intersection>
<intersection>117.5 110</intersection>
<intersection>125.5 31</intersection>
<intersection>165.5 111</intersection>
<intersection>174 55</intersection>
<intersection>223 112</intersection>
<intersection>232.5 56</intersection>
<intersection>278 113</intersection>
<intersection>286.5 66</intersection>
<intersection>335 114</intersection>
<intersection>344.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-21,-128.5,-21,-121</points>
<intersection>-128.5 5</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-21,-128.5,-19.5,-128.5</points>
<connection>
<GID>1553</GID>
<name>IN_1</name></connection>
<intersection>-21 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>27.5,-129.5,27.5,-121</points>
<intersection>-129.5 21</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>27.5,-129.5,29,-129.5</points>
<connection>
<GID>1555</GID>
<name>IN_1</name></connection>
<intersection>27.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>75,-128.5,75,-121</points>
<intersection>-128.5 53</intersection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>125.5,-128.5,125.5,-121</points>
<intersection>-128.5 115</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>75,-128.5,75.5,-128.5</points>
<connection>
<GID>1557</GID>
<name>IN_1</name></connection>
<intersection>75 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>174,-128,174,-121</points>
<connection>
<GID>1561</GID>
<name>IN_1</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>232.5,-130,232.5,-121</points>
<connection>
<GID>1563</GID>
<name>IN_1</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>286.5,-129,286.5,-121</points>
<intersection>-129 118</intersection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>344.5,-129.5,344.5,-121</points>
<connection>
<GID>1567</GID>
<name>IN_1</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-29.5,-123,-29.5,-121</points>
<connection>
<GID>1552</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>20,-123,20,-121</points>
<connection>
<GID>1554</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>68,-123,68,-121</points>
<connection>
<GID>1556</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>117.5,-123,117.5,-121</points>
<connection>
<GID>1558</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>165.5,-123,165.5,-121</points>
<connection>
<GID>1560</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>223,-123,223,-121</points>
<connection>
<GID>1562</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>278,-123,278,-121</points>
<connection>
<GID>1564</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>335,-123,335,-121</points>
<connection>
<GID>1566</GID>
<name>clock</name></connection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>125.5,-128.5,126,-128.5</points>
<connection>
<GID>1559</GID>
<name>IN_1</name></connection>
<intersection>125.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>286,-129,286.5,-129</points>
<connection>
<GID>1565</GID>
<name>IN_1</name></connection>
<intersection>286.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-126.5,75.5,-120</points>
<connection>
<GID>1557</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-120,75.5,-120</points>
<connection>
<GID>1556</GID>
<name>OUT_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>892</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-126.5,125,-120</points>
<intersection>-126.5 1</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-126.5,126,-126.5</points>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123.5,-120,125,-120</points>
<connection>
<GID>1558</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>893</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-126,173.5,-120</points>
<intersection>-126 5</intersection>
<intersection>-120 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>171.5,-120,173.5,-120</points>
<connection>
<GID>1560</GID>
<name>OUT_0</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>173.5,-126,174,-126</points>
<connection>
<GID>1561</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>894</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-128,232,-120</points>
<intersection>-128 1</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232,-128,232.5,-128</points>
<connection>
<GID>1563</GID>
<name>IN_0</name></connection>
<intersection>232 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,-120,232,-120</points>
<connection>
<GID>1562</GID>
<name>OUT_0</name></connection>
<intersection>232 0</intersection></hsegment></shape></wire>
<wire>
<ID>895</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-127,285.5,-120</points>
<intersection>-127 4</intersection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>284,-120,285.5,-120</points>
<connection>
<GID>1564</GID>
<name>OUT_0</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>285.5,-127,286,-127</points>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>896</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,-127.5,344,-120</points>
<intersection>-127.5 1</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,-127.5,344.5,-127.5</points>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection>
<intersection>344 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341,-120,344,-120</points>
<connection>
<GID>1566</GID>
<name>OUT_0</name></connection>
<intersection>344 0</intersection></hsegment></shape></wire>
<wire>
<ID>897</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,-120,-65.5,-89.5</points>
<intersection>-120 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,-120,-61,-120</points>
<connection>
<GID>1568</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-89.5,-65.5,-89.5</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>898</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-140.5,-22,-134</points>
<intersection>-140.5 1</intersection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-140.5,-19.5,-140.5</points>
<connection>
<GID>1570</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-23.5,-134,-22,-134</points>
<connection>
<GID>1569</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>899</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-141.5,27,-134</points>
<intersection>-141.5 1</intersection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-141.5,29,-141.5</points>
<connection>
<GID>1572</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-134,27,-134</points>
<connection>
<GID>1571</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>900</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,-135,344.5,-135</points>
<connection>
<GID>1585</GID>
<name>OUT</name></connection>
<intersection>-29.5 107</intersection>
<intersection>-21 4</intersection>
<intersection>20 108</intersection>
<intersection>27.5 16</intersection>
<intersection>68 109</intersection>
<intersection>75 23</intersection>
<intersection>117.5 110</intersection>
<intersection>125.5 31</intersection>
<intersection>165.5 111</intersection>
<intersection>174 55</intersection>
<intersection>223 112</intersection>
<intersection>232.5 56</intersection>
<intersection>278 113</intersection>
<intersection>286.5 66</intersection>
<intersection>335 114</intersection>
<intersection>344.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-21,-142.5,-21,-135</points>
<intersection>-142.5 5</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-21,-142.5,-19.5,-142.5</points>
<connection>
<GID>1570</GID>
<name>IN_1</name></connection>
<intersection>-21 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>27.5,-143.5,27.5,-135</points>
<intersection>-143.5 21</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>27.5,-143.5,29,-143.5</points>
<connection>
<GID>1572</GID>
<name>IN_1</name></connection>
<intersection>27.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>75,-142.5,75,-135</points>
<intersection>-142.5 53</intersection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>125.5,-142.5,125.5,-135</points>
<intersection>-142.5 115</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>75,-142.5,75.5,-142.5</points>
<connection>
<GID>1574</GID>
<name>IN_1</name></connection>
<intersection>75 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>174,-142,174,-135</points>
<connection>
<GID>1578</GID>
<name>IN_1</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>232.5,-144,232.5,-135</points>
<connection>
<GID>1580</GID>
<name>IN_1</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>286.5,-143,286.5,-135</points>
<intersection>-143 118</intersection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>344.5,-143.5,344.5,-135</points>
<connection>
<GID>1584</GID>
<name>IN_1</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-29.5,-137,-29.5,-135</points>
<connection>
<GID>1569</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>20,-137,20,-135</points>
<connection>
<GID>1571</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>68,-137,68,-135</points>
<connection>
<GID>1573</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>117.5,-137,117.5,-135</points>
<connection>
<GID>1575</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>165.5,-137,165.5,-135</points>
<connection>
<GID>1577</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>223,-137,223,-135</points>
<connection>
<GID>1579</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>278,-137,278,-135</points>
<connection>
<GID>1581</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>335,-137,335,-135</points>
<connection>
<GID>1583</GID>
<name>clock</name></connection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>125.5,-142.5,126,-142.5</points>
<connection>
<GID>1576</GID>
<name>IN_1</name></connection>
<intersection>125.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>286,-143,286.5,-143</points>
<connection>
<GID>1582</GID>
<name>IN_1</name></connection>
<intersection>286.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>901</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-140.5,75.5,-134</points>
<connection>
<GID>1574</GID>
<name>IN_0</name></connection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>74,-134,75.5,-134</points>
<connection>
<GID>1573</GID>
<name>OUT_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>902</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-140.5,125,-134</points>
<intersection>-140.5 1</intersection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-140.5,126,-140.5</points>
<connection>
<GID>1576</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123.5,-134,125,-134</points>
<connection>
<GID>1575</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>903</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-140,173.5,-134</points>
<intersection>-140 5</intersection>
<intersection>-134 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>171.5,-134,173.5,-134</points>
<connection>
<GID>1577</GID>
<name>OUT_0</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>173.5,-140,174,-140</points>
<connection>
<GID>1578</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>904</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-142,232,-134</points>
<intersection>-142 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232,-142,232.5,-142</points>
<connection>
<GID>1580</GID>
<name>IN_0</name></connection>
<intersection>232 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,-134,232,-134</points>
<connection>
<GID>1579</GID>
<name>OUT_0</name></connection>
<intersection>232 0</intersection></hsegment></shape></wire>
<wire>
<ID>905</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-141,285.5,-134</points>
<intersection>-141 4</intersection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>284,-134,285.5,-134</points>
<connection>
<GID>1581</GID>
<name>OUT_0</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>285.5,-141,286,-141</points>
<connection>
<GID>1582</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>906</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,-141.5,344,-134</points>
<intersection>-141.5 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,-141.5,344.5,-141.5</points>
<connection>
<GID>1584</GID>
<name>IN_0</name></connection>
<intersection>344 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341,-134,344,-134</points>
<connection>
<GID>1583</GID>
<name>OUT_0</name></connection>
<intersection>344 0</intersection></hsegment></shape></wire>
<wire>
<ID>907</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-134,-66.5,-90.5</points>
<intersection>-134 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,-134,-61,-134</points>
<connection>
<GID>1585</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-90.5,-66.5,-90.5</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-158,-22.5,-151.5</points>
<intersection>-158 1</intersection>
<intersection>-151.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22.5,-158,-20,-158</points>
<connection>
<GID>1587</GID>
<name>IN_0</name></connection>
<intersection>-22.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-24,-151.5,-22.5,-151.5</points>
<connection>
<GID>1586</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>909</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-159,26.5,-151.5</points>
<intersection>-159 1</intersection>
<intersection>-151.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-159,28.5,-159</points>
<connection>
<GID>1589</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-151.5,26.5,-151.5</points>
<connection>
<GID>1588</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>910</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55.5,-152.5,344,-152.5</points>
<connection>
<GID>1602</GID>
<name>OUT</name></connection>
<intersection>-30 107</intersection>
<intersection>-21.5 4</intersection>
<intersection>19.5 108</intersection>
<intersection>27 16</intersection>
<intersection>67.5 109</intersection>
<intersection>74.5 23</intersection>
<intersection>117 110</intersection>
<intersection>125 31</intersection>
<intersection>165 111</intersection>
<intersection>173.5 55</intersection>
<intersection>222.5 112</intersection>
<intersection>232 56</intersection>
<intersection>277.5 113</intersection>
<intersection>286 66</intersection>
<intersection>334.5 114</intersection>
<intersection>344 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-21.5,-160,-21.5,-152.5</points>
<intersection>-160 5</intersection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-21.5,-160,-20,-160</points>
<connection>
<GID>1587</GID>
<name>IN_1</name></connection>
<intersection>-21.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>27,-161,27,-152.5</points>
<intersection>-161 21</intersection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>27,-161,28.5,-161</points>
<connection>
<GID>1589</GID>
<name>IN_1</name></connection>
<intersection>27 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>74.5,-160,74.5,-152.5</points>
<intersection>-160 53</intersection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>125,-160,125,-152.5</points>
<intersection>-160 115</intersection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>74.5,-160,75,-160</points>
<connection>
<GID>1591</GID>
<name>IN_1</name></connection>
<intersection>74.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>173.5,-159.5,173.5,-152.5</points>
<connection>
<GID>1595</GID>
<name>IN_1</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>232,-161.5,232,-152.5</points>
<connection>
<GID>1597</GID>
<name>IN_1</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>286,-160.5,286,-152.5</points>
<intersection>-160.5 118</intersection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>344,-161,344,-152.5</points>
<connection>
<GID>1601</GID>
<name>IN_1</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-30,-154.5,-30,-152.5</points>
<connection>
<GID>1586</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>19.5,-154.5,19.5,-152.5</points>
<connection>
<GID>1588</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>67.5,-154.5,67.5,-152.5</points>
<connection>
<GID>1590</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>117,-154.5,117,-152.5</points>
<connection>
<GID>1592</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>165,-154.5,165,-152.5</points>
<connection>
<GID>1594</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>222.5,-154.5,222.5,-152.5</points>
<connection>
<GID>1596</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>277.5,-154.5,277.5,-152.5</points>
<connection>
<GID>1598</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>334.5,-154.5,334.5,-152.5</points>
<connection>
<GID>1600</GID>
<name>clock</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>125,-160,125.5,-160</points>
<connection>
<GID>1593</GID>
<name>IN_1</name></connection>
<intersection>125 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>285.5,-160.5,286,-160.5</points>
<connection>
<GID>1599</GID>
<name>IN_1</name></connection>
<intersection>286 66</intersection></hsegment></shape></wire>
<wire>
<ID>911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-158,75,-151.5</points>
<connection>
<GID>1591</GID>
<name>IN_0</name></connection>
<intersection>-151.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73.5,-151.5,75,-151.5</points>
<connection>
<GID>1590</GID>
<name>OUT_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-158,124.5,-151.5</points>
<intersection>-158 1</intersection>
<intersection>-151.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-158,125.5,-158</points>
<connection>
<GID>1593</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123,-151.5,124.5,-151.5</points>
<connection>
<GID>1592</GID>
<name>OUT_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>913</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-157.5,173,-151.5</points>
<intersection>-157.5 5</intersection>
<intersection>-151.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>171,-151.5,173,-151.5</points>
<connection>
<GID>1594</GID>
<name>OUT_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>173,-157.5,173.5,-157.5</points>
<connection>
<GID>1595</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>914</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-159.5,231.5,-151.5</points>
<intersection>-159.5 1</intersection>
<intersection>-151.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231.5,-159.5,232,-159.5</points>
<connection>
<GID>1597</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-151.5,231.5,-151.5</points>
<connection>
<GID>1596</GID>
<name>OUT_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285,-158.5,285,-151.5</points>
<intersection>-158.5 4</intersection>
<intersection>-151.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>283.5,-151.5,285,-151.5</points>
<connection>
<GID>1598</GID>
<name>OUT_0</name></connection>
<intersection>285 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>285,-158.5,285.5,-158.5</points>
<connection>
<GID>1599</GID>
<name>IN_0</name></connection>
<intersection>285 0</intersection></hsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343.5,-159,343.5,-151.5</points>
<intersection>-159 1</intersection>
<intersection>-151.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>343.5,-159,344,-159</points>
<connection>
<GID>1601</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>340.5,-151.5,343.5,-151.5</points>
<connection>
<GID>1600</GID>
<name>OUT_0</name></connection>
<intersection>343.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-151.5,-67.5,-91.5</points>
<intersection>-151.5 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-151.5,-61.5,-151.5</points>
<connection>
<GID>1602</GID>
<name>IN_0</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,-91.5,-67.5,-91.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-291.5,4,-285</points>
<intersection>-291.5 1</intersection>
<intersection>-285 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-291.5,6.5,-291.5</points>
<connection>
<GID>1655</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-285,4,-285</points>
<connection>
<GID>1654</GID>
<name>OUT_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-292.5,53,-285</points>
<intersection>-292.5 1</intersection>
<intersection>-285 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-292.5,55,-292.5</points>
<connection>
<GID>1657</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-285,53,-285</points>
<connection>
<GID>1656</GID>
<name>OUT_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>920</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29,-286,370.5,-286</points>
<connection>
<GID>1670</GID>
<name>OUT</name></connection>
<intersection>-3.5 107</intersection>
<intersection>5 4</intersection>
<intersection>46 108</intersection>
<intersection>53.5 16</intersection>
<intersection>94 109</intersection>
<intersection>101 23</intersection>
<intersection>143.5 110</intersection>
<intersection>151.5 31</intersection>
<intersection>191.5 111</intersection>
<intersection>200 55</intersection>
<intersection>249 112</intersection>
<intersection>258.5 56</intersection>
<intersection>304 113</intersection>
<intersection>312.5 66</intersection>
<intersection>361 114</intersection>
<intersection>370.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5,-293.5,5,-286</points>
<intersection>-293.5 5</intersection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>5,-293.5,6.5,-293.5</points>
<connection>
<GID>1655</GID>
<name>IN_1</name></connection>
<intersection>5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>53.5,-294.5,53.5,-286</points>
<intersection>-294.5 21</intersection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>53.5,-294.5,55,-294.5</points>
<connection>
<GID>1657</GID>
<name>IN_1</name></connection>
<intersection>53.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>101,-293.5,101,-286</points>
<intersection>-293.5 53</intersection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>151.5,-293.5,151.5,-286</points>
<intersection>-293.5 115</intersection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>101,-293.5,101.5,-293.5</points>
<connection>
<GID>1659</GID>
<name>IN_1</name></connection>
<intersection>101 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>200,-293,200,-286</points>
<connection>
<GID>1663</GID>
<name>IN_1</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>258.5,-295,258.5,-286</points>
<connection>
<GID>1665</GID>
<name>IN_1</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>312.5,-294,312.5,-286</points>
<intersection>-294 118</intersection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>370.5,-294.5,370.5,-286</points>
<connection>
<GID>1669</GID>
<name>IN_1</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-3.5,-288,-3.5,-286</points>
<connection>
<GID>1654</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>46,-288,46,-286</points>
<connection>
<GID>1656</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>94,-288,94,-286</points>
<connection>
<GID>1658</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>143.5,-288,143.5,-286</points>
<connection>
<GID>1660</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>191.5,-288,191.5,-286</points>
<connection>
<GID>1662</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>249,-288,249,-286</points>
<connection>
<GID>1664</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>304,-288,304,-286</points>
<connection>
<GID>1666</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>361,-288,361,-286</points>
<connection>
<GID>1668</GID>
<name>clock</name></connection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>151.5,-293.5,152,-293.5</points>
<connection>
<GID>1661</GID>
<name>IN_1</name></connection>
<intersection>151.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>312,-294,312.5,-294</points>
<connection>
<GID>1667</GID>
<name>IN_1</name></connection>
<intersection>312.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-291.5,101.5,-285</points>
<connection>
<GID>1659</GID>
<name>IN_0</name></connection>
<intersection>-285 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-285,101.5,-285</points>
<connection>
<GID>1658</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-291.5,151,-285</points>
<intersection>-291.5 1</intersection>
<intersection>-285 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-291.5,152,-291.5</points>
<connection>
<GID>1661</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149.5,-285,151,-285</points>
<connection>
<GID>1660</GID>
<name>OUT_0</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>923</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-291,199.5,-285</points>
<intersection>-291 5</intersection>
<intersection>-285 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197.5,-285,199.5,-285</points>
<connection>
<GID>1662</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>199.5,-291,200,-291</points>
<connection>
<GID>1663</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>924</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-293,258,-285</points>
<intersection>-293 1</intersection>
<intersection>-285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-293,258.5,-293</points>
<connection>
<GID>1665</GID>
<name>IN_0</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255,-285,258,-285</points>
<connection>
<GID>1664</GID>
<name>OUT_0</name></connection>
<intersection>258 0</intersection></hsegment></shape></wire>
<wire>
<ID>925</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-292,311.5,-285</points>
<intersection>-292 4</intersection>
<intersection>-285 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>310,-285,311.5,-285</points>
<connection>
<GID>1666</GID>
<name>OUT_0</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>311.5,-292,312,-292</points>
<connection>
<GID>1667</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>926</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,-292.5,370,-285</points>
<intersection>-292.5 1</intersection>
<intersection>-285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>370,-292.5,370.5,-292.5</points>
<connection>
<GID>1669</GID>
<name>IN_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>367,-285,370,-285</points>
<connection>
<GID>1668</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment></shape></wire>
<wire>
<ID>927</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-304.5,4,-298</points>
<intersection>-304.5 1</intersection>
<intersection>-298 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-304.5,6.5,-304.5</points>
<connection>
<GID>1672</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-298,4,-298</points>
<connection>
<GID>1671</GID>
<name>OUT_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>928</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-305.5,53,-298</points>
<intersection>-305.5 1</intersection>
<intersection>-298 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-305.5,55,-305.5</points>
<connection>
<GID>1674</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-298,53,-298</points>
<connection>
<GID>1673</GID>
<name>OUT_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>929</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29,-299,370.5,-299</points>
<connection>
<GID>1687</GID>
<name>OUT</name></connection>
<intersection>-3.5 107</intersection>
<intersection>5 4</intersection>
<intersection>46 108</intersection>
<intersection>53.5 16</intersection>
<intersection>94 109</intersection>
<intersection>101 23</intersection>
<intersection>143.5 110</intersection>
<intersection>151.5 31</intersection>
<intersection>191.5 111</intersection>
<intersection>200 55</intersection>
<intersection>249 112</intersection>
<intersection>258.5 56</intersection>
<intersection>304 113</intersection>
<intersection>312.5 66</intersection>
<intersection>361 114</intersection>
<intersection>370.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5,-306.5,5,-299</points>
<intersection>-306.5 5</intersection>
<intersection>-299 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>5,-306.5,6.5,-306.5</points>
<connection>
<GID>1672</GID>
<name>IN_1</name></connection>
<intersection>5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>53.5,-307.5,53.5,-299</points>
<intersection>-307.5 21</intersection>
<intersection>-299 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>53.5,-307.5,55,-307.5</points>
<connection>
<GID>1674</GID>
<name>IN_1</name></connection>
<intersection>53.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>101,-306.5,101,-299</points>
<intersection>-306.5 53</intersection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>151.5,-306.5,151.5,-299</points>
<intersection>-306.5 115</intersection>
<intersection>-299 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>101,-306.5,101.5,-306.5</points>
<connection>
<GID>1676</GID>
<name>IN_1</name></connection>
<intersection>101 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>200,-306,200,-299</points>
<connection>
<GID>1680</GID>
<name>IN_1</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>258.5,-308,258.5,-299</points>
<connection>
<GID>1682</GID>
<name>IN_1</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>312.5,-307,312.5,-299</points>
<intersection>-307 118</intersection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>370.5,-307.5,370.5,-299</points>
<connection>
<GID>1686</GID>
<name>IN_1</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-3.5,-301,-3.5,-299</points>
<connection>
<GID>1671</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>46,-301,46,-299</points>
<connection>
<GID>1673</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>94,-301,94,-299</points>
<connection>
<GID>1675</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>143.5,-301,143.5,-299</points>
<connection>
<GID>1677</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>191.5,-301,191.5,-299</points>
<connection>
<GID>1679</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>249,-301,249,-299</points>
<connection>
<GID>1681</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>304,-301,304,-299</points>
<connection>
<GID>1683</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>361,-301,361,-299</points>
<connection>
<GID>1685</GID>
<name>clock</name></connection>
<intersection>-299 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>151.5,-306.5,152,-306.5</points>
<connection>
<GID>1678</GID>
<name>IN_1</name></connection>
<intersection>151.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>312,-307,312.5,-307</points>
<connection>
<GID>1684</GID>
<name>IN_1</name></connection>
<intersection>312.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-304.5,101.5,-298</points>
<connection>
<GID>1676</GID>
<name>IN_0</name></connection>
<intersection>-298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-298,101.5,-298</points>
<connection>
<GID>1675</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-304.5,151,-298</points>
<intersection>-304.5 1</intersection>
<intersection>-298 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-304.5,152,-304.5</points>
<connection>
<GID>1678</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149.5,-298,151,-298</points>
<connection>
<GID>1677</GID>
<name>OUT_0</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-304,199.5,-298</points>
<intersection>-304 5</intersection>
<intersection>-298 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197.5,-298,199.5,-298</points>
<connection>
<GID>1679</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>199.5,-304,200,-304</points>
<connection>
<GID>1680</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-306,258,-298</points>
<intersection>-306 1</intersection>
<intersection>-298 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-306,258.5,-306</points>
<connection>
<GID>1682</GID>
<name>IN_0</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255,-298,258,-298</points>
<connection>
<GID>1681</GID>
<name>OUT_0</name></connection>
<intersection>258 0</intersection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-305,311.5,-298</points>
<intersection>-305 4</intersection>
<intersection>-298 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>310,-298,311.5,-298</points>
<connection>
<GID>1683</GID>
<name>OUT_0</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>311.5,-305,312,-305</points>
<connection>
<GID>1684</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,-305.5,370,-298</points>
<intersection>-305.5 1</intersection>
<intersection>-298 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>370,-305.5,370.5,-305.5</points>
<connection>
<GID>1686</GID>
<name>IN_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>367,-298,370,-298</points>
<connection>
<GID>1685</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-319,4,-312.5</points>
<intersection>-319 1</intersection>
<intersection>-312.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-319,6.5,-319</points>
<connection>
<GID>1689</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-312.5,4,-312.5</points>
<connection>
<GID>1688</GID>
<name>OUT_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-320,53,-312.5</points>
<intersection>-320 1</intersection>
<intersection>-312.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-320,55,-320</points>
<connection>
<GID>1691</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-312.5,53,-312.5</points>
<connection>
<GID>1690</GID>
<name>OUT_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29,-313.5,370.5,-313.5</points>
<connection>
<GID>1704</GID>
<name>OUT</name></connection>
<intersection>-3.5 107</intersection>
<intersection>5 4</intersection>
<intersection>46 108</intersection>
<intersection>53.5 16</intersection>
<intersection>94 109</intersection>
<intersection>101 23</intersection>
<intersection>143.5 110</intersection>
<intersection>151.5 31</intersection>
<intersection>191.5 111</intersection>
<intersection>200 55</intersection>
<intersection>249 112</intersection>
<intersection>258.5 56</intersection>
<intersection>304 113</intersection>
<intersection>312.5 66</intersection>
<intersection>361 114</intersection>
<intersection>370.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5,-321,5,-313.5</points>
<intersection>-321 5</intersection>
<intersection>-313.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>5,-321,6.5,-321</points>
<connection>
<GID>1689</GID>
<name>IN_1</name></connection>
<intersection>5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>53.5,-322,53.5,-313.5</points>
<intersection>-322 21</intersection>
<intersection>-313.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>53.5,-322,55,-322</points>
<connection>
<GID>1691</GID>
<name>IN_1</name></connection>
<intersection>53.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>101,-321,101,-313.5</points>
<intersection>-321 53</intersection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>151.5,-321,151.5,-313.5</points>
<intersection>-321 115</intersection>
<intersection>-313.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>101,-321,101.5,-321</points>
<connection>
<GID>1693</GID>
<name>IN_1</name></connection>
<intersection>101 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>200,-320.5,200,-313.5</points>
<connection>
<GID>1697</GID>
<name>IN_1</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>258.5,-322.5,258.5,-313.5</points>
<connection>
<GID>1699</GID>
<name>IN_1</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>312.5,-321.5,312.5,-313.5</points>
<intersection>-321.5 118</intersection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>370.5,-322,370.5,-313.5</points>
<connection>
<GID>1703</GID>
<name>IN_1</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-3.5,-315.5,-3.5,-313.5</points>
<connection>
<GID>1688</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>46,-315.5,46,-313.5</points>
<connection>
<GID>1690</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>94,-315.5,94,-313.5</points>
<connection>
<GID>1692</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>143.5,-315.5,143.5,-313.5</points>
<connection>
<GID>1694</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>191.5,-315.5,191.5,-313.5</points>
<connection>
<GID>1696</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>249,-315.5,249,-313.5</points>
<connection>
<GID>1698</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>304,-315.5,304,-313.5</points>
<connection>
<GID>1700</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>361,-315.5,361,-313.5</points>
<connection>
<GID>1702</GID>
<name>clock</name></connection>
<intersection>-313.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>151.5,-321,152,-321</points>
<connection>
<GID>1695</GID>
<name>IN_1</name></connection>
<intersection>151.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>312,-321.5,312.5,-321.5</points>
<connection>
<GID>1701</GID>
<name>IN_1</name></connection>
<intersection>312.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-319,101.5,-312.5</points>
<connection>
<GID>1693</GID>
<name>IN_0</name></connection>
<intersection>-312.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>100,-312.5,101.5,-312.5</points>
<connection>
<GID>1692</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-319,151,-312.5</points>
<intersection>-319 1</intersection>
<intersection>-312.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-319,152,-319</points>
<connection>
<GID>1695</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149.5,-312.5,151,-312.5</points>
<connection>
<GID>1694</GID>
<name>OUT_0</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-318.5,199.5,-312.5</points>
<intersection>-318.5 5</intersection>
<intersection>-312.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197.5,-312.5,199.5,-312.5</points>
<connection>
<GID>1696</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>199.5,-318.5,200,-318.5</points>
<connection>
<GID>1697</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-320.5,258,-312.5</points>
<intersection>-320.5 1</intersection>
<intersection>-312.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-320.5,258.5,-320.5</points>
<connection>
<GID>1699</GID>
<name>IN_0</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255,-312.5,258,-312.5</points>
<connection>
<GID>1698</GID>
<name>OUT_0</name></connection>
<intersection>258 0</intersection></hsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-319.5,311.5,-312.5</points>
<intersection>-319.5 4</intersection>
<intersection>-312.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>310,-312.5,311.5,-312.5</points>
<connection>
<GID>1700</GID>
<name>OUT_0</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>311.5,-319.5,312,-319.5</points>
<connection>
<GID>1701</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,-320,370,-312.5</points>
<intersection>-320 1</intersection>
<intersection>-312.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>370,-320,370.5,-320</points>
<connection>
<GID>1703</GID>
<name>IN_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>367,-312.5,370,-312.5</points>
<connection>
<GID>1702</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-331.5,3.5,-325</points>
<intersection>-331.5 1</intersection>
<intersection>-325 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-331.5,6,-331.5</points>
<connection>
<GID>1706</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2,-325,3.5,-325</points>
<connection>
<GID>1705</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-332.5,52.5,-325</points>
<intersection>-332.5 1</intersection>
<intersection>-325 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-332.5,54.5,-332.5</points>
<connection>
<GID>1708</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,-325,52.5,-325</points>
<connection>
<GID>1707</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>947</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,-326,370,-326</points>
<connection>
<GID>1721</GID>
<name>OUT</name></connection>
<intersection>-4 107</intersection>
<intersection>4.5 4</intersection>
<intersection>45.5 108</intersection>
<intersection>53 16</intersection>
<intersection>93.5 109</intersection>
<intersection>100.5 23</intersection>
<intersection>143 110</intersection>
<intersection>151 31</intersection>
<intersection>191 111</intersection>
<intersection>199.5 55</intersection>
<intersection>248.5 112</intersection>
<intersection>258 56</intersection>
<intersection>303.5 113</intersection>
<intersection>312 66</intersection>
<intersection>360.5 114</intersection>
<intersection>370 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>4.5,-333.5,4.5,-326</points>
<intersection>-333.5 5</intersection>
<intersection>-326 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4.5,-333.5,6,-333.5</points>
<connection>
<GID>1706</GID>
<name>IN_1</name></connection>
<intersection>4.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>53,-334.5,53,-326</points>
<intersection>-334.5 21</intersection>
<intersection>-326 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>53,-334.5,54.5,-334.5</points>
<connection>
<GID>1708</GID>
<name>IN_1</name></connection>
<intersection>53 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>100.5,-333.5,100.5,-326</points>
<intersection>-333.5 53</intersection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>151,-333.5,151,-326</points>
<intersection>-333.5 115</intersection>
<intersection>-326 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>100.5,-333.5,101,-333.5</points>
<connection>
<GID>1710</GID>
<name>IN_1</name></connection>
<intersection>100.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>199.5,-333,199.5,-326</points>
<connection>
<GID>1714</GID>
<name>IN_1</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>258,-335,258,-326</points>
<connection>
<GID>1716</GID>
<name>IN_1</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>312,-334,312,-326</points>
<intersection>-334 118</intersection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>370,-334.5,370,-326</points>
<connection>
<GID>1720</GID>
<name>IN_1</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-4,-328,-4,-326</points>
<connection>
<GID>1705</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>45.5,-328,45.5,-326</points>
<connection>
<GID>1707</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>93.5,-328,93.5,-326</points>
<connection>
<GID>1709</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>143,-328,143,-326</points>
<connection>
<GID>1711</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>191,-328,191,-326</points>
<connection>
<GID>1713</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>248.5,-328,248.5,-326</points>
<connection>
<GID>1715</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>303.5,-328,303.5,-326</points>
<connection>
<GID>1717</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>360.5,-328,360.5,-326</points>
<connection>
<GID>1719</GID>
<name>clock</name></connection>
<intersection>-326 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>151,-333.5,151.5,-333.5</points>
<connection>
<GID>1712</GID>
<name>IN_1</name></connection>
<intersection>151 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>311.5,-334,312,-334</points>
<connection>
<GID>1718</GID>
<name>IN_1</name></connection>
<intersection>312 66</intersection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-331.5,101,-325</points>
<connection>
<GID>1710</GID>
<name>IN_0</name></connection>
<intersection>-325 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-325,101,-325</points>
<connection>
<GID>1709</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-331.5,150.5,-325</points>
<intersection>-331.5 1</intersection>
<intersection>-325 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-331.5,151.5,-331.5</points>
<connection>
<GID>1712</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-325,150.5,-325</points>
<connection>
<GID>1711</GID>
<name>OUT_0</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-331,199,-325</points>
<intersection>-331 5</intersection>
<intersection>-325 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197,-325,199,-325</points>
<connection>
<GID>1713</GID>
<name>OUT_0</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>199,-331,199.5,-331</points>
<connection>
<GID>1714</GID>
<name>IN_0</name></connection>
<intersection>199 0</intersection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-333,257.5,-325</points>
<intersection>-333 1</intersection>
<intersection>-325 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-333,258,-333</points>
<connection>
<GID>1716</GID>
<name>IN_0</name></connection>
<intersection>257.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>254.5,-325,257.5,-325</points>
<connection>
<GID>1715</GID>
<name>OUT_0</name></connection>
<intersection>257.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-332,311,-325</points>
<intersection>-332 4</intersection>
<intersection>-325 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309.5,-325,311,-325</points>
<connection>
<GID>1717</GID>
<name>OUT_0</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>311,-332,311.5,-332</points>
<connection>
<GID>1718</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369.5,-332.5,369.5,-325</points>
<intersection>-332.5 1</intersection>
<intersection>-325 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369.5,-332.5,370,-332.5</points>
<connection>
<GID>1720</GID>
<name>IN_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366.5,-325,369.5,-325</points>
<connection>
<GID>1719</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-344.5,3,-338</points>
<intersection>-344.5 1</intersection>
<intersection>-338 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-344.5,5.5,-344.5</points>
<connection>
<GID>1723</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-338,3,-338</points>
<connection>
<GID>1722</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-345.5,52,-338</points>
<intersection>-345.5 1</intersection>
<intersection>-338 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-345.5,54,-345.5</points>
<connection>
<GID>1725</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51,-338,52,-338</points>
<connection>
<GID>1724</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-339,369.5,-339</points>
<connection>
<GID>1738</GID>
<name>OUT</name></connection>
<intersection>-4.5 107</intersection>
<intersection>4 4</intersection>
<intersection>45 108</intersection>
<intersection>52.5 16</intersection>
<intersection>93 109</intersection>
<intersection>100 23</intersection>
<intersection>142.5 110</intersection>
<intersection>150.5 31</intersection>
<intersection>190.5 111</intersection>
<intersection>199 55</intersection>
<intersection>248 112</intersection>
<intersection>257.5 56</intersection>
<intersection>303 113</intersection>
<intersection>311.5 66</intersection>
<intersection>360 114</intersection>
<intersection>369.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>4,-346.5,4,-339</points>
<intersection>-346.5 5</intersection>
<intersection>-339 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4,-346.5,5.5,-346.5</points>
<connection>
<GID>1723</GID>
<name>IN_1</name></connection>
<intersection>4 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>52.5,-347.5,52.5,-339</points>
<intersection>-347.5 21</intersection>
<intersection>-339 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>52.5,-347.5,54,-347.5</points>
<connection>
<GID>1725</GID>
<name>IN_1</name></connection>
<intersection>52.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>100,-346.5,100,-339</points>
<intersection>-346.5 53</intersection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>150.5,-346.5,150.5,-339</points>
<intersection>-346.5 115</intersection>
<intersection>-339 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>100,-346.5,100.5,-346.5</points>
<connection>
<GID>1727</GID>
<name>IN_1</name></connection>
<intersection>100 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>199,-346,199,-339</points>
<connection>
<GID>1731</GID>
<name>IN_1</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>257.5,-348,257.5,-339</points>
<connection>
<GID>1733</GID>
<name>IN_1</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>311.5,-347,311.5,-339</points>
<intersection>-347 118</intersection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>369.5,-347.5,369.5,-339</points>
<connection>
<GID>1737</GID>
<name>IN_1</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-4.5,-341,-4.5,-339</points>
<connection>
<GID>1722</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>45,-341,45,-339</points>
<connection>
<GID>1724</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>93,-341,93,-339</points>
<connection>
<GID>1726</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>142.5,-341,142.5,-339</points>
<connection>
<GID>1728</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>190.5,-341,190.5,-339</points>
<connection>
<GID>1730</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>248,-341,248,-339</points>
<connection>
<GID>1732</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>303,-341,303,-339</points>
<connection>
<GID>1734</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>360,-341,360,-339</points>
<connection>
<GID>1736</GID>
<name>clock</name></connection>
<intersection>-339 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>150.5,-346.5,151,-346.5</points>
<connection>
<GID>1729</GID>
<name>IN_1</name></connection>
<intersection>150.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>311,-347,311.5,-347</points>
<connection>
<GID>1735</GID>
<name>IN_1</name></connection>
<intersection>311.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-344.5,100.5,-338</points>
<connection>
<GID>1727</GID>
<name>IN_0</name></connection>
<intersection>-338 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>99,-338,100.5,-338</points>
<connection>
<GID>1726</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-344.5,150,-338</points>
<intersection>-344.5 1</intersection>
<intersection>-338 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-344.5,151,-344.5</points>
<connection>
<GID>1729</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148.5,-338,150,-338</points>
<connection>
<GID>1728</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-344,198.5,-338</points>
<intersection>-344 5</intersection>
<intersection>-338 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196.5,-338,198.5,-338</points>
<connection>
<GID>1730</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>198.5,-344,199,-344</points>
<connection>
<GID>1731</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-346,257,-338</points>
<intersection>-346 1</intersection>
<intersection>-338 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-346,257.5,-346</points>
<connection>
<GID>1733</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>254,-338,257,-338</points>
<connection>
<GID>1732</GID>
<name>OUT_0</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-345,310.5,-338</points>
<intersection>-345 4</intersection>
<intersection>-338 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,-338,310.5,-338</points>
<connection>
<GID>1734</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>310.5,-345,311,-345</points>
<connection>
<GID>1735</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-345.5,369,-338</points>
<intersection>-345.5 1</intersection>
<intersection>-338 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369,-345.5,369.5,-345.5</points>
<connection>
<GID>1737</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366,-338,369,-338</points>
<connection>
<GID>1736</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-359.5,3,-353</points>
<intersection>-359.5 1</intersection>
<intersection>-353 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-359.5,5.5,-359.5</points>
<connection>
<GID>1604</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-353,3,-353</points>
<connection>
<GID>1603</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-360.5,52,-353</points>
<intersection>-360.5 1</intersection>
<intersection>-353 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-360.5,54,-360.5</points>
<connection>
<GID>1606</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51,-353,52,-353</points>
<connection>
<GID>1605</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>965</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-354,369.5,-354</points>
<connection>
<GID>1619</GID>
<name>OUT</name></connection>
<intersection>-4.5 107</intersection>
<intersection>4 4</intersection>
<intersection>45 108</intersection>
<intersection>52.5 16</intersection>
<intersection>93 109</intersection>
<intersection>100 23</intersection>
<intersection>142.5 110</intersection>
<intersection>150.5 31</intersection>
<intersection>190.5 111</intersection>
<intersection>199 55</intersection>
<intersection>248 112</intersection>
<intersection>257.5 56</intersection>
<intersection>303 113</intersection>
<intersection>311.5 66</intersection>
<intersection>360 114</intersection>
<intersection>369.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>4,-361.5,4,-354</points>
<intersection>-361.5 5</intersection>
<intersection>-354 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4,-361.5,5.5,-361.5</points>
<connection>
<GID>1604</GID>
<name>IN_1</name></connection>
<intersection>4 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>52.5,-362.5,52.5,-354</points>
<intersection>-362.5 21</intersection>
<intersection>-354 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>52.5,-362.5,54,-362.5</points>
<connection>
<GID>1606</GID>
<name>IN_1</name></connection>
<intersection>52.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>100,-361.5,100,-354</points>
<intersection>-361.5 53</intersection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>150.5,-361.5,150.5,-354</points>
<intersection>-361.5 115</intersection>
<intersection>-354 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>100,-361.5,100.5,-361.5</points>
<connection>
<GID>1608</GID>
<name>IN_1</name></connection>
<intersection>100 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>199,-361,199,-354</points>
<connection>
<GID>1612</GID>
<name>IN_1</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>257.5,-363,257.5,-354</points>
<connection>
<GID>1614</GID>
<name>IN_1</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>311.5,-362,311.5,-354</points>
<intersection>-362 118</intersection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>369.5,-362.5,369.5,-354</points>
<connection>
<GID>1618</GID>
<name>IN_1</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-4.5,-356,-4.5,-354</points>
<connection>
<GID>1603</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>45,-356,45,-354</points>
<connection>
<GID>1605</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>93,-356,93,-354</points>
<connection>
<GID>1607</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>142.5,-356,142.5,-354</points>
<connection>
<GID>1609</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>190.5,-356,190.5,-354</points>
<connection>
<GID>1611</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>248,-356,248,-354</points>
<connection>
<GID>1613</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>303,-356,303,-354</points>
<connection>
<GID>1615</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>360,-356,360,-354</points>
<connection>
<GID>1617</GID>
<name>clock</name></connection>
<intersection>-354 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>150.5,-361.5,151,-361.5</points>
<connection>
<GID>1610</GID>
<name>IN_1</name></connection>
<intersection>150.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>311,-362,311.5,-362</points>
<connection>
<GID>1616</GID>
<name>IN_1</name></connection>
<intersection>311.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-359.5,100.5,-353</points>
<connection>
<GID>1608</GID>
<name>IN_0</name></connection>
<intersection>-353 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>99,-353,100.5,-353</points>
<connection>
<GID>1607</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-359.5,150,-353</points>
<intersection>-359.5 1</intersection>
<intersection>-353 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-359.5,151,-359.5</points>
<connection>
<GID>1610</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148.5,-353,150,-353</points>
<connection>
<GID>1609</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-359,198.5,-353</points>
<intersection>-359 5</intersection>
<intersection>-353 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196.5,-353,198.5,-353</points>
<connection>
<GID>1611</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>198.5,-359,199,-359</points>
<connection>
<GID>1612</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-361,257,-353</points>
<intersection>-361 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-361,257.5,-361</points>
<connection>
<GID>1614</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>254,-353,257,-353</points>
<connection>
<GID>1613</GID>
<name>OUT_0</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-360,310.5,-353</points>
<intersection>-360 4</intersection>
<intersection>-353 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,-353,310.5,-353</points>
<connection>
<GID>1615</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>310.5,-360,311,-360</points>
<connection>
<GID>1616</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-360.5,369,-353</points>
<intersection>-360.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369,-360.5,369.5,-360.5</points>
<connection>
<GID>1618</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366,-353,369,-353</points>
<connection>
<GID>1617</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-373.5,3,-367</points>
<intersection>-373.5 1</intersection>
<intersection>-367 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-373.5,5.5,-373.5</points>
<connection>
<GID>1621</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-367,3,-367</points>
<connection>
<GID>1620</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-374.5,52,-367</points>
<intersection>-374.5 1</intersection>
<intersection>-367 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-374.5,54,-374.5</points>
<connection>
<GID>1623</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51,-367,52,-367</points>
<connection>
<GID>1622</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-368,369.5,-368</points>
<connection>
<GID>1636</GID>
<name>OUT</name></connection>
<intersection>-4.5 107</intersection>
<intersection>4 4</intersection>
<intersection>45 108</intersection>
<intersection>52.5 16</intersection>
<intersection>93 109</intersection>
<intersection>100 23</intersection>
<intersection>142.5 110</intersection>
<intersection>150.5 31</intersection>
<intersection>190.5 111</intersection>
<intersection>199 55</intersection>
<intersection>248 112</intersection>
<intersection>257.5 56</intersection>
<intersection>303 113</intersection>
<intersection>311.5 66</intersection>
<intersection>360 114</intersection>
<intersection>369.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>4,-375.5,4,-368</points>
<intersection>-375.5 5</intersection>
<intersection>-368 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4,-375.5,5.5,-375.5</points>
<connection>
<GID>1621</GID>
<name>IN_1</name></connection>
<intersection>4 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>52.5,-376.5,52.5,-368</points>
<intersection>-376.5 21</intersection>
<intersection>-368 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>52.5,-376.5,54,-376.5</points>
<connection>
<GID>1623</GID>
<name>IN_1</name></connection>
<intersection>52.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>100,-375.5,100,-368</points>
<intersection>-375.5 53</intersection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>150.5,-375.5,150.5,-368</points>
<intersection>-375.5 115</intersection>
<intersection>-368 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>100,-375.5,100.5,-375.5</points>
<connection>
<GID>1625</GID>
<name>IN_1</name></connection>
<intersection>100 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>199,-375,199,-368</points>
<connection>
<GID>1629</GID>
<name>IN_1</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>257.5,-377,257.5,-368</points>
<connection>
<GID>1631</GID>
<name>IN_1</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>311.5,-376,311.5,-368</points>
<intersection>-376 118</intersection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>369.5,-376.5,369.5,-368</points>
<connection>
<GID>1635</GID>
<name>IN_1</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-4.5,-370,-4.5,-368</points>
<connection>
<GID>1620</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>45,-370,45,-368</points>
<connection>
<GID>1622</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>93,-370,93,-368</points>
<connection>
<GID>1624</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>142.5,-370,142.5,-368</points>
<connection>
<GID>1626</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>190.5,-370,190.5,-368</points>
<connection>
<GID>1628</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>248,-370,248,-368</points>
<connection>
<GID>1630</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>303,-370,303,-368</points>
<connection>
<GID>1632</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>360,-370,360,-368</points>
<connection>
<GID>1634</GID>
<name>clock</name></connection>
<intersection>-368 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>150.5,-375.5,151,-375.5</points>
<connection>
<GID>1627</GID>
<name>IN_1</name></connection>
<intersection>150.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>311,-376,311.5,-376</points>
<connection>
<GID>1633</GID>
<name>IN_1</name></connection>
<intersection>311.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-373.5,100.5,-367</points>
<connection>
<GID>1625</GID>
<name>IN_0</name></connection>
<intersection>-367 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>99,-367,100.5,-367</points>
<connection>
<GID>1624</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-373.5,150,-367</points>
<intersection>-373.5 1</intersection>
<intersection>-367 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-373.5,151,-373.5</points>
<connection>
<GID>1627</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148.5,-367,150,-367</points>
<connection>
<GID>1626</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-373,198.5,-367</points>
<intersection>-373 5</intersection>
<intersection>-367 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196.5,-367,198.5,-367</points>
<connection>
<GID>1628</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>198.5,-373,199,-373</points>
<connection>
<GID>1629</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-375,257,-367</points>
<intersection>-375 1</intersection>
<intersection>-367 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-375,257.5,-375</points>
<connection>
<GID>1631</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>254,-367,257,-367</points>
<connection>
<GID>1630</GID>
<name>OUT_0</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-374,310.5,-367</points>
<intersection>-374 4</intersection>
<intersection>-367 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,-367,310.5,-367</points>
<connection>
<GID>1632</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>310.5,-374,311,-374</points>
<connection>
<GID>1633</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-374.5,369,-367</points>
<intersection>-374.5 1</intersection>
<intersection>-367 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369,-374.5,369.5,-374.5</points>
<connection>
<GID>1635</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366,-367,369,-367</points>
<connection>
<GID>1634</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-391,2.5,-384.5</points>
<intersection>-391 1</intersection>
<intersection>-384.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-391,5,-391</points>
<connection>
<GID>1638</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1,-384.5,2.5,-384.5</points>
<connection>
<GID>1637</GID>
<name>OUT_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-392,51.5,-384.5</points>
<intersection>-392 1</intersection>
<intersection>-384.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-392,53.5,-392</points>
<connection>
<GID>1640</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-384.5,51.5,-384.5</points>
<connection>
<GID>1639</GID>
<name>OUT_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30.5,-385.5,369,-385.5</points>
<connection>
<GID>1653</GID>
<name>OUT</name></connection>
<intersection>-5 107</intersection>
<intersection>3.5 4</intersection>
<intersection>44.5 108</intersection>
<intersection>52 16</intersection>
<intersection>92.5 109</intersection>
<intersection>99.5 23</intersection>
<intersection>142 110</intersection>
<intersection>150 31</intersection>
<intersection>190 111</intersection>
<intersection>198.5 55</intersection>
<intersection>247.5 112</intersection>
<intersection>257 56</intersection>
<intersection>302.5 113</intersection>
<intersection>311 66</intersection>
<intersection>359.5 114</intersection>
<intersection>369 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>3.5,-393,3.5,-385.5</points>
<intersection>-393 5</intersection>
<intersection>-385.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>3.5,-393,5,-393</points>
<connection>
<GID>1638</GID>
<name>IN_1</name></connection>
<intersection>3.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>52,-394,52,-385.5</points>
<intersection>-394 21</intersection>
<intersection>-385.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>52,-394,53.5,-394</points>
<connection>
<GID>1640</GID>
<name>IN_1</name></connection>
<intersection>52 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>99.5,-393,99.5,-385.5</points>
<intersection>-393 53</intersection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>150,-393,150,-385.5</points>
<intersection>-393 115</intersection>
<intersection>-385.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>99.5,-393,100,-393</points>
<connection>
<GID>1642</GID>
<name>IN_1</name></connection>
<intersection>99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>198.5,-392.5,198.5,-385.5</points>
<connection>
<GID>1646</GID>
<name>IN_1</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>257,-394.5,257,-385.5</points>
<connection>
<GID>1648</GID>
<name>IN_1</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>311,-393.5,311,-385.5</points>
<intersection>-393.5 118</intersection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>369,-394,369,-385.5</points>
<connection>
<GID>1652</GID>
<name>IN_1</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-5,-387.5,-5,-385.5</points>
<connection>
<GID>1637</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>44.5,-387.5,44.5,-385.5</points>
<connection>
<GID>1639</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>92.5,-387.5,92.5,-385.5</points>
<connection>
<GID>1641</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>142,-387.5,142,-385.5</points>
<connection>
<GID>1643</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>190,-387.5,190,-385.5</points>
<connection>
<GID>1645</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>247.5,-387.5,247.5,-385.5</points>
<connection>
<GID>1647</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>302.5,-387.5,302.5,-385.5</points>
<connection>
<GID>1649</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>359.5,-387.5,359.5,-385.5</points>
<connection>
<GID>1651</GID>
<name>clock</name></connection>
<intersection>-385.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>150,-393,150.5,-393</points>
<connection>
<GID>1644</GID>
<name>IN_1</name></connection>
<intersection>150 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>310.5,-393.5,311,-393.5</points>
<connection>
<GID>1650</GID>
<name>IN_1</name></connection>
<intersection>311 66</intersection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-391,100,-384.5</points>
<connection>
<GID>1642</GID>
<name>IN_0</name></connection>
<intersection>-384.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>98.5,-384.5,100,-384.5</points>
<connection>
<GID>1641</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-391,149.5,-384.5</points>
<intersection>-391 1</intersection>
<intersection>-384.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-391,150.5,-391</points>
<connection>
<GID>1644</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148,-384.5,149.5,-384.5</points>
<connection>
<GID>1643</GID>
<name>OUT_0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-390.5,198,-384.5</points>
<intersection>-390.5 5</intersection>
<intersection>-384.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196,-384.5,198,-384.5</points>
<connection>
<GID>1645</GID>
<name>OUT_0</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>198,-390.5,198.5,-390.5</points>
<connection>
<GID>1646</GID>
<name>IN_0</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-392.5,256.5,-384.5</points>
<intersection>-392.5 1</intersection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,-392.5,257,-392.5</points>
<connection>
<GID>1648</GID>
<name>IN_0</name></connection>
<intersection>256.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>253.5,-384.5,256.5,-384.5</points>
<connection>
<GID>1647</GID>
<name>OUT_0</name></connection>
<intersection>256.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-391.5,310,-384.5</points>
<intersection>-391.5 4</intersection>
<intersection>-384.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>308.5,-384.5,310,-384.5</points>
<connection>
<GID>1649</GID>
<name>OUT_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>310,-391.5,310.5,-391.5</points>
<connection>
<GID>1650</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368.5,-392,368.5,-384.5</points>
<intersection>-392 1</intersection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>368.5,-392,369,-392</points>
<connection>
<GID>1652</GID>
<name>IN_0</name></connection>
<intersection>368.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>365.5,-384.5,368.5,-384.5</points>
<connection>
<GID>1651</GID>
<name>OUT_0</name></connection>
<intersection>368.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-323,-53,-285</points>
<intersection>-323 2</intersection>
<intersection>-285 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53,-285,-35,-285</points>
<connection>
<GID>1670</GID>
<name>IN_0</name></connection>
<intersection>-53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-323,-53,-323</points>
<connection>
<GID>195</GID>
<name>OUT_7</name></connection>
<intersection>-53 0</intersection></hsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-324,-51.5,-298</points>
<intersection>-324 2</intersection>
<intersection>-298 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-298,-35,-298</points>
<connection>
<GID>1687</GID>
<name>IN_0</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-324,-51.5,-324</points>
<connection>
<GID>195</GID>
<name>OUT_6</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,-325,-50,-312.5</points>
<intersection>-325 2</intersection>
<intersection>-312.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,-312.5,-35,-312.5</points>
<connection>
<GID>1704</GID>
<name>IN_0</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-325,-50,-325</points>
<connection>
<GID>195</GID>
<name>OUT_5</name></connection>
<intersection>-50 0</intersection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-78.5,-326,-36,-326</points>
<connection>
<GID>195</GID>
<name>OUT_4</name></connection>
<intersection>-36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-36,-326,-36,-325</points>
<intersection>-326 1</intersection>
<intersection>-325 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-36,-325,-35.5,-325</points>
<connection>
<GID>1721</GID>
<name>IN_0</name></connection>
<intersection>-36 3</intersection></hsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50.5,-338,-50.5,-327</points>
<intersection>-338 1</intersection>
<intersection>-327 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50.5,-338,-36,-338</points>
<connection>
<GID>1738</GID>
<name>IN_0</name></connection>
<intersection>-50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-327,-50.5,-327</points>
<connection>
<GID>195</GID>
<name>OUT_3</name></connection>
<intersection>-50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-353,-52,-328</points>
<intersection>-353 1</intersection>
<intersection>-328 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-353,-36,-353</points>
<connection>
<GID>1619</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-328,-52,-328</points>
<connection>
<GID>195</GID>
<name>OUT_2</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-367,-53.5,-329</points>
<intersection>-367 1</intersection>
<intersection>-329 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53.5,-367,-36,-367</points>
<connection>
<GID>1636</GID>
<name>IN_0</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-329,-53.5,-329</points>
<connection>
<GID>195</GID>
<name>OUT_1</name></connection>
<intersection>-53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-384.5,-55.5,-330</points>
<intersection>-384.5 1</intersection>
<intersection>-330 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,-384.5,-36.5,-384.5</points>
<connection>
<GID>1653</GID>
<name>IN_0</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,-330,-55.5,-330</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>-55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-578,-13,-571.5</points>
<intersection>-578 1</intersection>
<intersection>-571.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-578,-10.5,-578</points>
<connection>
<GID>1791</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14.5,-571.5,-13,-571.5</points>
<connection>
<GID>1790</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-579,36,-571.5</points>
<intersection>-579 1</intersection>
<intersection>-571.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-579,38,-579</points>
<connection>
<GID>1793</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-571.5,36,-571.5</points>
<connection>
<GID>1792</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-572.5,353.5,-572.5</points>
<connection>
<GID>1806</GID>
<name>OUT</name></connection>
<intersection>-20.5 107</intersection>
<intersection>-12 4</intersection>
<intersection>29 108</intersection>
<intersection>36.5 16</intersection>
<intersection>77 109</intersection>
<intersection>84 23</intersection>
<intersection>126.5 110</intersection>
<intersection>134.5 31</intersection>
<intersection>174.5 111</intersection>
<intersection>183 55</intersection>
<intersection>232 112</intersection>
<intersection>241.5 56</intersection>
<intersection>287 113</intersection>
<intersection>295.5 66</intersection>
<intersection>344 114</intersection>
<intersection>353.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-580,-12,-572.5</points>
<intersection>-580 5</intersection>
<intersection>-572.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-580,-10.5,-580</points>
<connection>
<GID>1791</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36.5,-581,36.5,-572.5</points>
<intersection>-581 21</intersection>
<intersection>-572.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36.5,-581,38,-581</points>
<connection>
<GID>1793</GID>
<name>IN_1</name></connection>
<intersection>36.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84,-580,84,-572.5</points>
<intersection>-580 53</intersection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134.5,-580,134.5,-572.5</points>
<intersection>-580 115</intersection>
<intersection>-572.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84,-580,84.5,-580</points>
<connection>
<GID>1795</GID>
<name>IN_1</name></connection>
<intersection>84 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183,-579.5,183,-572.5</points>
<connection>
<GID>1799</GID>
<name>IN_1</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241.5,-581.5,241.5,-572.5</points>
<connection>
<GID>1801</GID>
<name>IN_1</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295.5,-580.5,295.5,-572.5</points>
<intersection>-580.5 118</intersection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353.5,-581,353.5,-572.5</points>
<connection>
<GID>1805</GID>
<name>IN_1</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20.5,-574.5,-20.5,-572.5</points>
<connection>
<GID>1790</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29,-574.5,29,-572.5</points>
<connection>
<GID>1792</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77,-574.5,77,-572.5</points>
<connection>
<GID>1794</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126.5,-574.5,126.5,-572.5</points>
<connection>
<GID>1796</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174.5,-574.5,174.5,-572.5</points>
<connection>
<GID>1798</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232,-574.5,232,-572.5</points>
<connection>
<GID>1800</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287,-574.5,287,-572.5</points>
<connection>
<GID>1802</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344,-574.5,344,-572.5</points>
<connection>
<GID>1804</GID>
<name>clock</name></connection>
<intersection>-572.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134.5,-580,135,-580</points>
<connection>
<GID>1797</GID>
<name>IN_1</name></connection>
<intersection>134.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295,-580.5,295.5,-580.5</points>
<connection>
<GID>1803</GID>
<name>IN_1</name></connection>
<intersection>295.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1001</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-578,84.5,-571.5</points>
<connection>
<GID>1795</GID>
<name>IN_0</name></connection>
<intersection>-571.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83,-571.5,84.5,-571.5</points>
<connection>
<GID>1794</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-578,134,-571.5</points>
<intersection>-578 1</intersection>
<intersection>-571.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-578,135,-578</points>
<connection>
<GID>1797</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-571.5,134,-571.5</points>
<connection>
<GID>1796</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1003</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-577.5,182.5,-571.5</points>
<intersection>-577.5 5</intersection>
<intersection>-571.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180.5,-571.5,182.5,-571.5</points>
<connection>
<GID>1798</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-577.5,183,-577.5</points>
<connection>
<GID>1799</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-579.5,241,-571.5</points>
<intersection>-579.5 1</intersection>
<intersection>-571.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-579.5,241.5,-579.5</points>
<connection>
<GID>1801</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-571.5,241,-571.5</points>
<connection>
<GID>1800</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-578.5,294.5,-571.5</points>
<intersection>-578.5 4</intersection>
<intersection>-571.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-571.5,294.5,-571.5</points>
<connection>
<GID>1802</GID>
<name>OUT_0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-578.5,295,-578.5</points>
<connection>
<GID>1803</GID>
<name>IN_0</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-579,353,-571.5</points>
<intersection>-579 1</intersection>
<intersection>-571.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-579,353.5,-579</points>
<connection>
<GID>1805</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-571.5,353,-571.5</points>
<connection>
<GID>1804</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-591,-13,-584.5</points>
<intersection>-591 1</intersection>
<intersection>-584.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-591,-10.5,-591</points>
<connection>
<GID>1808</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14.5,-584.5,-13,-584.5</points>
<connection>
<GID>1807</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-592,36,-584.5</points>
<intersection>-592 1</intersection>
<intersection>-584.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-592,38,-592</points>
<connection>
<GID>1810</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-584.5,36,-584.5</points>
<connection>
<GID>1809</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-585.5,353.5,-585.5</points>
<connection>
<GID>1823</GID>
<name>OUT</name></connection>
<intersection>-20.5 107</intersection>
<intersection>-12 4</intersection>
<intersection>29 108</intersection>
<intersection>36.5 16</intersection>
<intersection>77 109</intersection>
<intersection>84 23</intersection>
<intersection>126.5 110</intersection>
<intersection>134.5 31</intersection>
<intersection>174.5 111</intersection>
<intersection>183 55</intersection>
<intersection>232 112</intersection>
<intersection>241.5 56</intersection>
<intersection>287 113</intersection>
<intersection>295.5 66</intersection>
<intersection>344 114</intersection>
<intersection>353.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-593,-12,-585.5</points>
<intersection>-593 5</intersection>
<intersection>-585.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-593,-10.5,-593</points>
<connection>
<GID>1808</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36.5,-594,36.5,-585.5</points>
<intersection>-594 21</intersection>
<intersection>-585.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36.5,-594,38,-594</points>
<connection>
<GID>1810</GID>
<name>IN_1</name></connection>
<intersection>36.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84,-593,84,-585.5</points>
<intersection>-593 53</intersection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134.5,-593,134.5,-585.5</points>
<intersection>-593 115</intersection>
<intersection>-585.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84,-593,84.5,-593</points>
<connection>
<GID>1812</GID>
<name>IN_1</name></connection>
<intersection>84 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183,-592.5,183,-585.5</points>
<connection>
<GID>1816</GID>
<name>IN_1</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241.5,-594.5,241.5,-585.5</points>
<connection>
<GID>1818</GID>
<name>IN_1</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295.5,-593.5,295.5,-585.5</points>
<intersection>-593.5 118</intersection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353.5,-594,353.5,-585.5</points>
<connection>
<GID>1822</GID>
<name>IN_1</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20.5,-587.5,-20.5,-585.5</points>
<connection>
<GID>1807</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29,-587.5,29,-585.5</points>
<connection>
<GID>1809</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77,-587.5,77,-585.5</points>
<connection>
<GID>1811</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126.5,-587.5,126.5,-585.5</points>
<connection>
<GID>1813</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174.5,-587.5,174.5,-585.5</points>
<connection>
<GID>1815</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232,-587.5,232,-585.5</points>
<connection>
<GID>1817</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287,-587.5,287,-585.5</points>
<connection>
<GID>1819</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344,-587.5,344,-585.5</points>
<connection>
<GID>1821</GID>
<name>clock</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134.5,-593,135,-593</points>
<connection>
<GID>1814</GID>
<name>IN_1</name></connection>
<intersection>134.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295,-593.5,295.5,-593.5</points>
<connection>
<GID>1820</GID>
<name>IN_1</name></connection>
<intersection>295.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-591,84.5,-584.5</points>
<connection>
<GID>1812</GID>
<name>IN_0</name></connection>
<intersection>-584.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83,-584.5,84.5,-584.5</points>
<connection>
<GID>1811</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-591,134,-584.5</points>
<intersection>-591 1</intersection>
<intersection>-584.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-591,135,-591</points>
<connection>
<GID>1814</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-584.5,134,-584.5</points>
<connection>
<GID>1813</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-590.5,182.5,-584.5</points>
<intersection>-590.5 5</intersection>
<intersection>-584.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180.5,-584.5,182.5,-584.5</points>
<connection>
<GID>1815</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-590.5,183,-590.5</points>
<connection>
<GID>1816</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-592.5,241,-584.5</points>
<intersection>-592.5 1</intersection>
<intersection>-584.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-592.5,241.5,-592.5</points>
<connection>
<GID>1818</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-584.5,241,-584.5</points>
<connection>
<GID>1817</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-591.5,294.5,-584.5</points>
<intersection>-591.5 4</intersection>
<intersection>-584.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-584.5,294.5,-584.5</points>
<connection>
<GID>1819</GID>
<name>OUT_0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-591.5,295,-591.5</points>
<connection>
<GID>1820</GID>
<name>IN_0</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-592,353,-584.5</points>
<intersection>-592 1</intersection>
<intersection>-584.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-592,353.5,-592</points>
<connection>
<GID>1822</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-584.5,353,-584.5</points>
<connection>
<GID>1821</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-605.5,-13,-599</points>
<intersection>-605.5 1</intersection>
<intersection>-599 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-605.5,-10.5,-605.5</points>
<connection>
<GID>1825</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14.5,-599,-13,-599</points>
<connection>
<GID>1824</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-606.5,36,-599</points>
<intersection>-606.5 1</intersection>
<intersection>-599 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-606.5,38,-606.5</points>
<connection>
<GID>1827</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-599,36,-599</points>
<connection>
<GID>1826</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-600,353.5,-600</points>
<connection>
<GID>1840</GID>
<name>OUT</name></connection>
<intersection>-20.5 107</intersection>
<intersection>-12 4</intersection>
<intersection>29 108</intersection>
<intersection>36.5 16</intersection>
<intersection>77 109</intersection>
<intersection>84 23</intersection>
<intersection>126.5 110</intersection>
<intersection>134.5 31</intersection>
<intersection>174.5 111</intersection>
<intersection>183 55</intersection>
<intersection>232 112</intersection>
<intersection>241.5 56</intersection>
<intersection>287 113</intersection>
<intersection>295.5 66</intersection>
<intersection>344 114</intersection>
<intersection>353.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-607.5,-12,-600</points>
<intersection>-607.5 5</intersection>
<intersection>-600 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-607.5,-10.5,-607.5</points>
<connection>
<GID>1825</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36.5,-608.5,36.5,-600</points>
<intersection>-608.5 21</intersection>
<intersection>-600 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36.5,-608.5,38,-608.5</points>
<connection>
<GID>1827</GID>
<name>IN_1</name></connection>
<intersection>36.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84,-607.5,84,-600</points>
<intersection>-607.5 53</intersection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134.5,-607.5,134.5,-600</points>
<intersection>-607.5 115</intersection>
<intersection>-600 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84,-607.5,84.5,-607.5</points>
<connection>
<GID>1829</GID>
<name>IN_1</name></connection>
<intersection>84 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183,-607,183,-600</points>
<connection>
<GID>1833</GID>
<name>IN_1</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241.5,-609,241.5,-600</points>
<connection>
<GID>1835</GID>
<name>IN_1</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295.5,-608,295.5,-600</points>
<intersection>-608 118</intersection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353.5,-608.5,353.5,-600</points>
<connection>
<GID>1839</GID>
<name>IN_1</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20.5,-602,-20.5,-600</points>
<connection>
<GID>1824</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29,-602,29,-600</points>
<connection>
<GID>1826</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77,-602,77,-600</points>
<connection>
<GID>1828</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126.5,-602,126.5,-600</points>
<connection>
<GID>1830</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174.5,-602,174.5,-600</points>
<connection>
<GID>1832</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232,-602,232,-600</points>
<connection>
<GID>1834</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287,-602,287,-600</points>
<connection>
<GID>1836</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344,-602,344,-600</points>
<connection>
<GID>1838</GID>
<name>clock</name></connection>
<intersection>-600 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134.5,-607.5,135,-607.5</points>
<connection>
<GID>1831</GID>
<name>IN_1</name></connection>
<intersection>134.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295,-608,295.5,-608</points>
<connection>
<GID>1837</GID>
<name>IN_1</name></connection>
<intersection>295.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-605.5,84.5,-599</points>
<connection>
<GID>1829</GID>
<name>IN_0</name></connection>
<intersection>-599 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83,-599,84.5,-599</points>
<connection>
<GID>1828</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-605.5,134,-599</points>
<intersection>-605.5 1</intersection>
<intersection>-599 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-605.5,135,-605.5</points>
<connection>
<GID>1831</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-599,134,-599</points>
<connection>
<GID>1830</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-605,182.5,-599</points>
<intersection>-605 5</intersection>
<intersection>-599 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180.5,-599,182.5,-599</points>
<connection>
<GID>1832</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-605,183,-605</points>
<connection>
<GID>1833</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-607,241,-599</points>
<intersection>-607 1</intersection>
<intersection>-599 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-607,241.5,-607</points>
<connection>
<GID>1835</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-599,241,-599</points>
<connection>
<GID>1834</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-606,294.5,-599</points>
<intersection>-606 4</intersection>
<intersection>-599 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-599,294.5,-599</points>
<connection>
<GID>1836</GID>
<name>OUT_0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-606,295,-606</points>
<connection>
<GID>1837</GID>
<name>IN_0</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-606.5,353,-599</points>
<intersection>-606.5 1</intersection>
<intersection>-599 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-606.5,353.5,-606.5</points>
<connection>
<GID>1839</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-599,353,-599</points>
<connection>
<GID>1838</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-618,-13.5,-611.5</points>
<intersection>-618 1</intersection>
<intersection>-611.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-618,-11,-618</points>
<connection>
<GID>1842</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15,-611.5,-13.5,-611.5</points>
<connection>
<GID>1841</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-619,35.5,-611.5</points>
<intersection>-619 1</intersection>
<intersection>-611.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-619,37.5,-619</points>
<connection>
<GID>1844</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34.5,-611.5,35.5,-611.5</points>
<connection>
<GID>1843</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46.5,-612.5,353,-612.5</points>
<connection>
<GID>1857</GID>
<name>OUT</name></connection>
<intersection>-21 107</intersection>
<intersection>-12.5 4</intersection>
<intersection>28.5 108</intersection>
<intersection>36 16</intersection>
<intersection>76.5 109</intersection>
<intersection>83.5 23</intersection>
<intersection>126 110</intersection>
<intersection>134 31</intersection>
<intersection>174 111</intersection>
<intersection>182.5 55</intersection>
<intersection>231.5 112</intersection>
<intersection>241 56</intersection>
<intersection>286.5 113</intersection>
<intersection>295 66</intersection>
<intersection>343.5 114</intersection>
<intersection>353 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12.5,-620,-12.5,-612.5</points>
<intersection>-620 5</intersection>
<intersection>-612.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,-620,-11,-620</points>
<connection>
<GID>1842</GID>
<name>IN_1</name></connection>
<intersection>-12.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36,-621,36,-612.5</points>
<intersection>-621 21</intersection>
<intersection>-612.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36,-621,37.5,-621</points>
<connection>
<GID>1844</GID>
<name>IN_1</name></connection>
<intersection>36 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83.5,-620,83.5,-612.5</points>
<intersection>-620 53</intersection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134,-620,134,-612.5</points>
<intersection>-620 115</intersection>
<intersection>-612.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83.5,-620,84,-620</points>
<connection>
<GID>1846</GID>
<name>IN_1</name></connection>
<intersection>83.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182.5,-619.5,182.5,-612.5</points>
<connection>
<GID>1850</GID>
<name>IN_1</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241,-621.5,241,-612.5</points>
<connection>
<GID>1852</GID>
<name>IN_1</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295,-620.5,295,-612.5</points>
<intersection>-620.5 118</intersection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353,-621,353,-612.5</points>
<connection>
<GID>1856</GID>
<name>IN_1</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21,-614.5,-21,-612.5</points>
<connection>
<GID>1841</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28.5,-614.5,28.5,-612.5</points>
<connection>
<GID>1843</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76.5,-614.5,76.5,-612.5</points>
<connection>
<GID>1845</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126,-614.5,126,-612.5</points>
<connection>
<GID>1847</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174,-614.5,174,-612.5</points>
<connection>
<GID>1849</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231.5,-614.5,231.5,-612.5</points>
<connection>
<GID>1851</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286.5,-614.5,286.5,-612.5</points>
<connection>
<GID>1853</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343.5,-614.5,343.5,-612.5</points>
<connection>
<GID>1855</GID>
<name>clock</name></connection>
<intersection>-612.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134,-620,134.5,-620</points>
<connection>
<GID>1848</GID>
<name>IN_1</name></connection>
<intersection>134 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294.5,-620.5,295,-620.5</points>
<connection>
<GID>1854</GID>
<name>IN_1</name></connection>
<intersection>295 66</intersection></hsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-618,84,-611.5</points>
<connection>
<GID>1846</GID>
<name>IN_0</name></connection>
<intersection>-611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82.5,-611.5,84,-611.5</points>
<connection>
<GID>1845</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-618,133.5,-611.5</points>
<intersection>-618 1</intersection>
<intersection>-611.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-618,134.5,-618</points>
<connection>
<GID>1848</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,-611.5,133.5,-611.5</points>
<connection>
<GID>1847</GID>
<name>OUT_0</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-617.5,182,-611.5</points>
<intersection>-617.5 5</intersection>
<intersection>-611.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180,-611.5,182,-611.5</points>
<connection>
<GID>1849</GID>
<name>OUT_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182,-617.5,182.5,-617.5</points>
<connection>
<GID>1850</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-619.5,240.5,-611.5</points>
<intersection>-619.5 1</intersection>
<intersection>-611.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240.5,-619.5,241,-619.5</points>
<connection>
<GID>1852</GID>
<name>IN_0</name></connection>
<intersection>240.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237.5,-611.5,240.5,-611.5</points>
<connection>
<GID>1851</GID>
<name>OUT_0</name></connection>
<intersection>240.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-618.5,294,-611.5</points>
<intersection>-618.5 4</intersection>
<intersection>-611.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292.5,-611.5,294,-611.5</points>
<connection>
<GID>1853</GID>
<name>OUT_0</name></connection>
<intersection>294 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294,-618.5,294.5,-618.5</points>
<connection>
<GID>1854</GID>
<name>IN_0</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352.5,-619,352.5,-611.5</points>
<intersection>-619 1</intersection>
<intersection>-611.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352.5,-619,353,-619</points>
<connection>
<GID>1856</GID>
<name>IN_0</name></connection>
<intersection>352.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-611.5,352.5,-611.5</points>
<connection>
<GID>1855</GID>
<name>OUT_0</name></connection>
<intersection>352.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-631,-14,-624.5</points>
<intersection>-631 1</intersection>
<intersection>-624.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-631,-11.5,-631</points>
<connection>
<GID>1859</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-624.5,-14,-624.5</points>
<connection>
<GID>1858</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-632,35,-624.5</points>
<intersection>-632 1</intersection>
<intersection>-624.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-632,37,-632</points>
<connection>
<GID>1861</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-624.5,35,-624.5</points>
<connection>
<GID>1860</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-625.5,352.5,-625.5</points>
<connection>
<GID>1874</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-633,-13,-625.5</points>
<intersection>-633 5</intersection>
<intersection>-625.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-633,-11.5,-633</points>
<connection>
<GID>1859</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-634,35.5,-625.5</points>
<intersection>-634 21</intersection>
<intersection>-625.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-634,37,-634</points>
<connection>
<GID>1861</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-633,83,-625.5</points>
<intersection>-633 53</intersection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-633,133.5,-625.5</points>
<intersection>-633 115</intersection>
<intersection>-625.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-633,83.5,-633</points>
<connection>
<GID>1863</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-632.5,182,-625.5</points>
<connection>
<GID>1867</GID>
<name>IN_1</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-634.5,240.5,-625.5</points>
<connection>
<GID>1869</GID>
<name>IN_1</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-633.5,294.5,-625.5</points>
<intersection>-633.5 118</intersection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-634,352.5,-625.5</points>
<connection>
<GID>1873</GID>
<name>IN_1</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-627.5,-21.5,-625.5</points>
<connection>
<GID>1858</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-627.5,28,-625.5</points>
<connection>
<GID>1860</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-627.5,76,-625.5</points>
<connection>
<GID>1862</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-627.5,125.5,-625.5</points>
<connection>
<GID>1864</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-627.5,173.5,-625.5</points>
<connection>
<GID>1866</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-627.5,231,-625.5</points>
<connection>
<GID>1868</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-627.5,286,-625.5</points>
<connection>
<GID>1870</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-627.5,343,-625.5</points>
<connection>
<GID>1872</GID>
<name>clock</name></connection>
<intersection>-625.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-633,134,-633</points>
<connection>
<GID>1865</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-633.5,294.5,-633.5</points>
<connection>
<GID>1871</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-631,83.5,-624.5</points>
<connection>
<GID>1863</GID>
<name>IN_0</name></connection>
<intersection>-624.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-624.5,83.5,-624.5</points>
<connection>
<GID>1862</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-631,133,-624.5</points>
<intersection>-631 1</intersection>
<intersection>-624.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-631,134,-631</points>
<connection>
<GID>1865</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-624.5,133,-624.5</points>
<connection>
<GID>1864</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-630.5,181.5,-624.5</points>
<intersection>-630.5 5</intersection>
<intersection>-624.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-624.5,181.5,-624.5</points>
<connection>
<GID>1866</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-630.5,182,-630.5</points>
<connection>
<GID>1867</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-632.5,240,-624.5</points>
<intersection>-632.5 1</intersection>
<intersection>-624.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-632.5,240.5,-632.5</points>
<connection>
<GID>1869</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-624.5,240,-624.5</points>
<connection>
<GID>1868</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-631.5,293.5,-624.5</points>
<intersection>-631.5 4</intersection>
<intersection>-624.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-624.5,293.5,-624.5</points>
<connection>
<GID>1870</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-631.5,294,-631.5</points>
<connection>
<GID>1871</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-632,352,-624.5</points>
<intersection>-632 1</intersection>
<intersection>-624.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-632,352.5,-632</points>
<connection>
<GID>1873</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-624.5,352,-624.5</points>
<connection>
<GID>1872</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-646,-14,-639.5</points>
<intersection>-646 1</intersection>
<intersection>-639.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-646,-11.5,-646</points>
<connection>
<GID>1740</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-639.5,-14,-639.5</points>
<connection>
<GID>1739</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-647,35,-639.5</points>
<intersection>-647 1</intersection>
<intersection>-639.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-647,37,-647</points>
<connection>
<GID>1742</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-639.5,35,-639.5</points>
<connection>
<GID>1741</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-640.5,352.5,-640.5</points>
<connection>
<GID>1755</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-648,-13,-640.5</points>
<intersection>-648 5</intersection>
<intersection>-640.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-648,-11.5,-648</points>
<connection>
<GID>1740</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-649,35.5,-640.5</points>
<intersection>-649 21</intersection>
<intersection>-640.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-649,37,-649</points>
<connection>
<GID>1742</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-648,83,-640.5</points>
<intersection>-648 53</intersection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-648,133.5,-640.5</points>
<intersection>-648 115</intersection>
<intersection>-640.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-648,83.5,-648</points>
<connection>
<GID>1744</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-647.5,182,-640.5</points>
<connection>
<GID>1748</GID>
<name>IN_1</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-649.5,240.5,-640.5</points>
<connection>
<GID>1750</GID>
<name>IN_1</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-648.5,294.5,-640.5</points>
<intersection>-648.5 118</intersection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-649,352.5,-640.5</points>
<connection>
<GID>1754</GID>
<name>IN_1</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-642.5,-21.5,-640.5</points>
<connection>
<GID>1739</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-642.5,28,-640.5</points>
<connection>
<GID>1741</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-642.5,76,-640.5</points>
<connection>
<GID>1743</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-642.5,125.5,-640.5</points>
<connection>
<GID>1745</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-642.5,173.5,-640.5</points>
<connection>
<GID>1747</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-642.5,231,-640.5</points>
<connection>
<GID>1749</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-642.5,286,-640.5</points>
<connection>
<GID>1751</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-642.5,343,-640.5</points>
<connection>
<GID>1753</GID>
<name>clock</name></connection>
<intersection>-640.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-648,134,-648</points>
<connection>
<GID>1746</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-648.5,294.5,-648.5</points>
<connection>
<GID>1752</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-646,83.5,-639.5</points>
<connection>
<GID>1744</GID>
<name>IN_0</name></connection>
<intersection>-639.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-639.5,83.5,-639.5</points>
<connection>
<GID>1743</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-646,133,-639.5</points>
<intersection>-646 1</intersection>
<intersection>-639.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-646,134,-646</points>
<connection>
<GID>1746</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-639.5,133,-639.5</points>
<connection>
<GID>1745</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-645.5,181.5,-639.5</points>
<intersection>-645.5 5</intersection>
<intersection>-639.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-639.5,181.5,-639.5</points>
<connection>
<GID>1747</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-645.5,182,-645.5</points>
<connection>
<GID>1748</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-647.5,240,-639.5</points>
<intersection>-647.5 1</intersection>
<intersection>-639.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-647.5,240.5,-647.5</points>
<connection>
<GID>1750</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-639.5,240,-639.5</points>
<connection>
<GID>1749</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-646.5,293.5,-639.5</points>
<intersection>-646.5 4</intersection>
<intersection>-639.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-639.5,293.5,-639.5</points>
<connection>
<GID>1751</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-646.5,294,-646.5</points>
<connection>
<GID>1752</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-647,352,-639.5</points>
<intersection>-647 1</intersection>
<intersection>-639.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-647,352.5,-647</points>
<connection>
<GID>1754</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-639.5,352,-639.5</points>
<connection>
<GID>1753</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-660,-14,-653.5</points>
<intersection>-660 1</intersection>
<intersection>-653.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-660,-11.5,-660</points>
<connection>
<GID>1757</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-653.5,-14,-653.5</points>
<connection>
<GID>1756</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-661,35,-653.5</points>
<intersection>-661 1</intersection>
<intersection>-653.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-661,37,-661</points>
<connection>
<GID>1759</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-653.5,35,-653.5</points>
<connection>
<GID>1758</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-654.5,352.5,-654.5</points>
<connection>
<GID>1772</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-662,-13,-654.5</points>
<intersection>-662 5</intersection>
<intersection>-654.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-662,-11.5,-662</points>
<connection>
<GID>1757</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-663,35.5,-654.5</points>
<intersection>-663 21</intersection>
<intersection>-654.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-663,37,-663</points>
<connection>
<GID>1759</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-662,83,-654.5</points>
<intersection>-662 53</intersection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-662,133.5,-654.5</points>
<intersection>-662 115</intersection>
<intersection>-654.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-662,83.5,-662</points>
<connection>
<GID>1761</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-661.5,182,-654.5</points>
<connection>
<GID>1765</GID>
<name>IN_1</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-663.5,240.5,-654.5</points>
<connection>
<GID>1767</GID>
<name>IN_1</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-662.5,294.5,-654.5</points>
<intersection>-662.5 118</intersection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-663,352.5,-654.5</points>
<connection>
<GID>1771</GID>
<name>IN_1</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-656.5,-21.5,-654.5</points>
<connection>
<GID>1756</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-656.5,28,-654.5</points>
<connection>
<GID>1758</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-656.5,76,-654.5</points>
<connection>
<GID>1760</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-656.5,125.5,-654.5</points>
<connection>
<GID>1762</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-656.5,173.5,-654.5</points>
<connection>
<GID>1764</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-656.5,231,-654.5</points>
<connection>
<GID>1766</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-656.5,286,-654.5</points>
<connection>
<GID>1768</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-656.5,343,-654.5</points>
<connection>
<GID>1770</GID>
<name>clock</name></connection>
<intersection>-654.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-662,134,-662</points>
<connection>
<GID>1763</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-662.5,294.5,-662.5</points>
<connection>
<GID>1769</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-660,83.5,-653.5</points>
<connection>
<GID>1761</GID>
<name>IN_0</name></connection>
<intersection>-653.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-653.5,83.5,-653.5</points>
<connection>
<GID>1760</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-660,133,-653.5</points>
<intersection>-660 1</intersection>
<intersection>-653.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-660,134,-660</points>
<connection>
<GID>1763</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-653.5,133,-653.5</points>
<connection>
<GID>1762</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-659.5,181.5,-653.5</points>
<intersection>-659.5 5</intersection>
<intersection>-653.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-653.5,181.5,-653.5</points>
<connection>
<GID>1764</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-659.5,182,-659.5</points>
<connection>
<GID>1765</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-661.5,240,-653.5</points>
<intersection>-661.5 1</intersection>
<intersection>-653.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-661.5,240.5,-661.5</points>
<connection>
<GID>1767</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-653.5,240,-653.5</points>
<connection>
<GID>1766</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-660.5,293.5,-653.5</points>
<intersection>-660.5 4</intersection>
<intersection>-653.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-653.5,293.5,-653.5</points>
<connection>
<GID>1768</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-660.5,294,-660.5</points>
<connection>
<GID>1769</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-661,352,-653.5</points>
<intersection>-661 1</intersection>
<intersection>-653.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-661,352.5,-661</points>
<connection>
<GID>1771</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-653.5,352,-653.5</points>
<connection>
<GID>1770</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-677.5,-14.5,-671</points>
<intersection>-677.5 1</intersection>
<intersection>-671 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-677.5,-12,-677.5</points>
<connection>
<GID>1774</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-671,-14.5,-671</points>
<connection>
<GID>1773</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-678.5,34.5,-671</points>
<intersection>-678.5 1</intersection>
<intersection>-671 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-678.5,36.5,-678.5</points>
<connection>
<GID>1776</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-671,34.5,-671</points>
<connection>
<GID>1775</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47.5,-672,352,-672</points>
<connection>
<GID>1789</GID>
<name>OUT</name></connection>
<intersection>-22 107</intersection>
<intersection>-13.5 4</intersection>
<intersection>27.5 108</intersection>
<intersection>35 16</intersection>
<intersection>75.5 109</intersection>
<intersection>82.5 23</intersection>
<intersection>125 110</intersection>
<intersection>133 31</intersection>
<intersection>173 111</intersection>
<intersection>181.5 55</intersection>
<intersection>230.5 112</intersection>
<intersection>240 56</intersection>
<intersection>285.5 113</intersection>
<intersection>294 66</intersection>
<intersection>342.5 114</intersection>
<intersection>352 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13.5,-679.5,-13.5,-672</points>
<intersection>-679.5 5</intersection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13.5,-679.5,-12,-679.5</points>
<connection>
<GID>1774</GID>
<name>IN_1</name></connection>
<intersection>-13.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35,-680.5,35,-672</points>
<intersection>-680.5 21</intersection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35,-680.5,36.5,-680.5</points>
<connection>
<GID>1776</GID>
<name>IN_1</name></connection>
<intersection>35 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>82.5,-679.5,82.5,-672</points>
<intersection>-679.5 53</intersection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133,-679.5,133,-672</points>
<intersection>-679.5 115</intersection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>82.5,-679.5,83,-679.5</points>
<connection>
<GID>1778</GID>
<name>IN_1</name></connection>
<intersection>82.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>181.5,-679,181.5,-672</points>
<connection>
<GID>1782</GID>
<name>IN_1</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240,-681,240,-672</points>
<connection>
<GID>1784</GID>
<name>IN_1</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294,-680,294,-672</points>
<intersection>-680 118</intersection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352,-680.5,352,-672</points>
<connection>
<GID>1788</GID>
<name>IN_1</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-22,-674,-22,-672</points>
<connection>
<GID>1773</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>27.5,-674,27.5,-672</points>
<connection>
<GID>1775</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>75.5,-674,75.5,-672</points>
<connection>
<GID>1777</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125,-674,125,-672</points>
<connection>
<GID>1779</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173,-674,173,-672</points>
<connection>
<GID>1781</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>230.5,-674,230.5,-672</points>
<connection>
<GID>1783</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>285.5,-674,285.5,-672</points>
<connection>
<GID>1785</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>342.5,-674,342.5,-672</points>
<connection>
<GID>1787</GID>
<name>clock</name></connection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133,-679.5,133.5,-679.5</points>
<connection>
<GID>1780</GID>
<name>IN_1</name></connection>
<intersection>133 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>293.5,-680,294,-680</points>
<connection>
<GID>1786</GID>
<name>IN_1</name></connection>
<intersection>294 66</intersection></hsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-677.5,83,-671</points>
<connection>
<GID>1778</GID>
<name>IN_0</name></connection>
<intersection>-671 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-671,83,-671</points>
<connection>
<GID>1777</GID>
<name>OUT_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-677.5,132.5,-671</points>
<intersection>-677.5 1</intersection>
<intersection>-671 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-677.5,133.5,-677.5</points>
<connection>
<GID>1780</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-671,132.5,-671</points>
<connection>
<GID>1779</GID>
<name>OUT_0</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-677,181,-671</points>
<intersection>-677 5</intersection>
<intersection>-671 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179,-671,181,-671</points>
<connection>
<GID>1781</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181,-677,181.5,-677</points>
<connection>
<GID>1782</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-679,239.5,-671</points>
<intersection>-679 1</intersection>
<intersection>-671 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-679,240,-679</points>
<connection>
<GID>1784</GID>
<name>IN_0</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-671,239.5,-671</points>
<connection>
<GID>1783</GID>
<name>OUT_0</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-678,293,-671</points>
<intersection>-678 4</intersection>
<intersection>-671 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-671,293,-671</points>
<connection>
<GID>1785</GID>
<name>OUT_0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-678,293.5,-678</points>
<connection>
<GID>1786</GID>
<name>IN_0</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,-678.5,351.5,-671</points>
<intersection>-678.5 1</intersection>
<intersection>-671 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,-678.5,352,-678.5</points>
<connection>
<GID>1788</GID>
<name>IN_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,-671,351.5,-671</points>
<connection>
<GID>1787</GID>
<name>OUT_0</name></connection>
<intersection>351.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-618,-63.5,-571.5</points>
<intersection>-618 2</intersection>
<intersection>-571.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-571.5,-52,-571.5</points>
<connection>
<GID>1806</GID>
<name>IN_0</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-618,-63.5,-618</points>
<connection>
<GID>332</GID>
<name>OUT_7</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-619,-62,-584.5</points>
<intersection>-619 2</intersection>
<intersection>-584.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-584.5,-52,-584.5</points>
<connection>
<GID>1823</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-619,-62,-619</points>
<connection>
<GID>332</GID>
<name>OUT_6</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-620,-60.5,-599</points>
<intersection>-620 2</intersection>
<intersection>-599 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60.5,-599,-52,-599</points>
<connection>
<GID>1840</GID>
<name>IN_0</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-620,-60.5,-620</points>
<connection>
<GID>332</GID>
<name>OUT_5</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-621,-59.5,-611.5</points>
<intersection>-621 2</intersection>
<intersection>-611.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-611.5,-52.5,-611.5</points>
<connection>
<GID>1857</GID>
<name>IN_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-621,-59.5,-621</points>
<connection>
<GID>332</GID>
<name>OUT_4</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-624.5,-60.5,-622</points>
<intersection>-624.5 1</intersection>
<intersection>-622 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60.5,-624.5,-53,-624.5</points>
<connection>
<GID>1874</GID>
<name>IN_0</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-622,-60.5,-622</points>
<connection>
<GID>332</GID>
<name>OUT_3</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-639.5,-62,-623</points>
<intersection>-639.5 1</intersection>
<intersection>-623 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-639.5,-53,-639.5</points>
<connection>
<GID>1755</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-623,-62,-623</points>
<connection>
<GID>332</GID>
<name>OUT_2</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-653.5,-63.5,-624</points>
<intersection>-653.5 2</intersection>
<intersection>-624 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-86,-624,-63.5,-624</points>
<connection>
<GID>332</GID>
<name>OUT_1</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63.5,-653.5,-53,-653.5</points>
<connection>
<GID>1772</GID>
<name>IN_0</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-671,-64.5,-625</points>
<intersection>-671 2</intersection>
<intersection>-625 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-86,-625,-64.5,-625</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-64.5,-671,-53.5,-671</points>
<connection>
<GID>1789</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-866.5,-9,-860</points>
<intersection>-866.5 1</intersection>
<intersection>-860 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-866.5,-6.5,-866.5</points>
<connection>
<GID>1927</GID>
<name>IN_0</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10.5,-860,-9,-860</points>
<connection>
<GID>1926</GID>
<name>OUT_0</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-867.5,40,-860</points>
<intersection>-867.5 1</intersection>
<intersection>-860 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-867.5,42,-867.5</points>
<connection>
<GID>1929</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,-860,40,-860</points>
<connection>
<GID>1928</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-861,357.5,-861</points>
<connection>
<GID>1942</GID>
<name>OUT</name></connection>
<intersection>-16.5 107</intersection>
<intersection>-8 4</intersection>
<intersection>33 108</intersection>
<intersection>40.5 16</intersection>
<intersection>81 109</intersection>
<intersection>88 23</intersection>
<intersection>130.5 110</intersection>
<intersection>138.5 31</intersection>
<intersection>178.5 111</intersection>
<intersection>187 55</intersection>
<intersection>236 112</intersection>
<intersection>245.5 56</intersection>
<intersection>291 113</intersection>
<intersection>299.5 66</intersection>
<intersection>348 114</intersection>
<intersection>357.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-8,-868.5,-8,-861</points>
<intersection>-868.5 5</intersection>
<intersection>-861 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-8,-868.5,-6.5,-868.5</points>
<connection>
<GID>1927</GID>
<name>IN_1</name></connection>
<intersection>-8 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>40.5,-869.5,40.5,-861</points>
<intersection>-869.5 21</intersection>
<intersection>-861 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>40.5,-869.5,42,-869.5</points>
<connection>
<GID>1929</GID>
<name>IN_1</name></connection>
<intersection>40.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>88,-868.5,88,-861</points>
<intersection>-868.5 53</intersection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>138.5,-868.5,138.5,-861</points>
<intersection>-868.5 115</intersection>
<intersection>-861 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>88,-868.5,88.5,-868.5</points>
<connection>
<GID>1931</GID>
<name>IN_1</name></connection>
<intersection>88 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>187,-868,187,-861</points>
<connection>
<GID>1935</GID>
<name>IN_1</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>245.5,-870,245.5,-861</points>
<connection>
<GID>1937</GID>
<name>IN_1</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>299.5,-869,299.5,-861</points>
<intersection>-869 118</intersection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>357.5,-869.5,357.5,-861</points>
<connection>
<GID>1941</GID>
<name>IN_1</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-16.5,-863,-16.5,-861</points>
<connection>
<GID>1926</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>33,-863,33,-861</points>
<connection>
<GID>1928</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>81,-863,81,-861</points>
<connection>
<GID>1930</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>130.5,-863,130.5,-861</points>
<connection>
<GID>1932</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>178.5,-863,178.5,-861</points>
<connection>
<GID>1934</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>236,-863,236,-861</points>
<connection>
<GID>1936</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>291,-863,291,-861</points>
<connection>
<GID>1938</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>348,-863,348,-861</points>
<connection>
<GID>1940</GID>
<name>clock</name></connection>
<intersection>-861 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>138.5,-868.5,139,-868.5</points>
<connection>
<GID>1933</GID>
<name>IN_1</name></connection>
<intersection>138.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>299,-869,299.5,-869</points>
<connection>
<GID>1939</GID>
<name>IN_1</name></connection>
<intersection>299.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-866.5,88.5,-860</points>
<connection>
<GID>1931</GID>
<name>IN_0</name></connection>
<intersection>-860 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>87,-860,88.5,-860</points>
<connection>
<GID>1930</GID>
<name>OUT_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-866.5,138,-860</points>
<intersection>-866.5 1</intersection>
<intersection>-860 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-866.5,139,-866.5</points>
<connection>
<GID>1933</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136.5,-860,138,-860</points>
<connection>
<GID>1932</GID>
<name>OUT_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-866,186.5,-860</points>
<intersection>-866 5</intersection>
<intersection>-860 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>184.5,-860,186.5,-860</points>
<connection>
<GID>1934</GID>
<name>OUT_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>186.5,-866,187,-866</points>
<connection>
<GID>1935</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-868,245,-860</points>
<intersection>-868 1</intersection>
<intersection>-860 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-868,245.5,-868</points>
<connection>
<GID>1937</GID>
<name>IN_0</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-860,245,-860</points>
<connection>
<GID>1936</GID>
<name>OUT_0</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-867,298.5,-860</points>
<intersection>-867 4</intersection>
<intersection>-860 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>297,-860,298.5,-860</points>
<connection>
<GID>1938</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>298.5,-867,299,-867</points>
<connection>
<GID>1939</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-867.5,357,-860</points>
<intersection>-867.5 1</intersection>
<intersection>-860 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-867.5,357.5,-867.5</points>
<connection>
<GID>1941</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-860,357,-860</points>
<connection>
<GID>1940</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-879.5,-9,-873</points>
<intersection>-879.5 1</intersection>
<intersection>-873 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-879.5,-6.5,-879.5</points>
<connection>
<GID>1944</GID>
<name>IN_0</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10.5,-873,-9,-873</points>
<connection>
<GID>1943</GID>
<name>OUT_0</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-880.5,40,-873</points>
<intersection>-880.5 1</intersection>
<intersection>-873 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-880.5,42,-880.5</points>
<connection>
<GID>1946</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,-873,40,-873</points>
<connection>
<GID>1945</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-874,357.5,-874</points>
<connection>
<GID>1959</GID>
<name>OUT</name></connection>
<intersection>-16.5 107</intersection>
<intersection>-8 4</intersection>
<intersection>33 108</intersection>
<intersection>40.5 16</intersection>
<intersection>81 109</intersection>
<intersection>88 23</intersection>
<intersection>130.5 110</intersection>
<intersection>138.5 31</intersection>
<intersection>178.5 111</intersection>
<intersection>187 55</intersection>
<intersection>236 112</intersection>
<intersection>245.5 56</intersection>
<intersection>291 113</intersection>
<intersection>299.5 66</intersection>
<intersection>348 114</intersection>
<intersection>357.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-8,-881.5,-8,-874</points>
<intersection>-881.5 5</intersection>
<intersection>-874 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-8,-881.5,-6.5,-881.5</points>
<connection>
<GID>1944</GID>
<name>IN_1</name></connection>
<intersection>-8 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>40.5,-882.5,40.5,-874</points>
<intersection>-882.5 21</intersection>
<intersection>-874 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>40.5,-882.5,42,-882.5</points>
<connection>
<GID>1946</GID>
<name>IN_1</name></connection>
<intersection>40.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>88,-881.5,88,-874</points>
<intersection>-881.5 53</intersection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>138.5,-881.5,138.5,-874</points>
<intersection>-881.5 115</intersection>
<intersection>-874 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>88,-881.5,88.5,-881.5</points>
<connection>
<GID>1948</GID>
<name>IN_1</name></connection>
<intersection>88 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>187,-881,187,-874</points>
<connection>
<GID>1952</GID>
<name>IN_1</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>245.5,-883,245.5,-874</points>
<connection>
<GID>1954</GID>
<name>IN_1</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>299.5,-882,299.5,-874</points>
<intersection>-882 118</intersection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>357.5,-882.5,357.5,-874</points>
<connection>
<GID>1958</GID>
<name>IN_1</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-16.5,-876,-16.5,-874</points>
<connection>
<GID>1943</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>33,-876,33,-874</points>
<connection>
<GID>1945</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>81,-876,81,-874</points>
<connection>
<GID>1947</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>130.5,-876,130.5,-874</points>
<connection>
<GID>1949</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>178.5,-876,178.5,-874</points>
<connection>
<GID>1951</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>236,-876,236,-874</points>
<connection>
<GID>1953</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>291,-876,291,-874</points>
<connection>
<GID>1955</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>348,-876,348,-874</points>
<connection>
<GID>1957</GID>
<name>clock</name></connection>
<intersection>-874 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>138.5,-881.5,139,-881.5</points>
<connection>
<GID>1950</GID>
<name>IN_1</name></connection>
<intersection>138.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>299,-882,299.5,-882</points>
<connection>
<GID>1956</GID>
<name>IN_1</name></connection>
<intersection>299.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-879.5,88.5,-873</points>
<connection>
<GID>1948</GID>
<name>IN_0</name></connection>
<intersection>-873 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>87,-873,88.5,-873</points>
<connection>
<GID>1947</GID>
<name>OUT_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-879.5,138,-873</points>
<intersection>-879.5 1</intersection>
<intersection>-873 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-879.5,139,-879.5</points>
<connection>
<GID>1950</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136.5,-873,138,-873</points>
<connection>
<GID>1949</GID>
<name>OUT_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-879,186.5,-873</points>
<intersection>-879 5</intersection>
<intersection>-873 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>184.5,-873,186.5,-873</points>
<connection>
<GID>1951</GID>
<name>OUT_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>186.5,-879,187,-879</points>
<connection>
<GID>1952</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-881,245,-873</points>
<intersection>-881 1</intersection>
<intersection>-873 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-881,245.5,-881</points>
<connection>
<GID>1954</GID>
<name>IN_0</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-873,245,-873</points>
<connection>
<GID>1953</GID>
<name>OUT_0</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-880,298.5,-873</points>
<intersection>-880 4</intersection>
<intersection>-873 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>297,-873,298.5,-873</points>
<connection>
<GID>1955</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>298.5,-880,299,-880</points>
<connection>
<GID>1956</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-880.5,357,-873</points>
<intersection>-880.5 1</intersection>
<intersection>-873 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-880.5,357.5,-880.5</points>
<connection>
<GID>1958</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-873,357,-873</points>
<connection>
<GID>1957</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-894,-9,-887.5</points>
<intersection>-894 1</intersection>
<intersection>-887.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-894,-6.5,-894</points>
<connection>
<GID>1961</GID>
<name>IN_0</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10.5,-887.5,-9,-887.5</points>
<connection>
<GID>1960</GID>
<name>OUT_0</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-895,40,-887.5</points>
<intersection>-895 1</intersection>
<intersection>-887.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-895,42,-895</points>
<connection>
<GID>1963</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,-887.5,40,-887.5</points>
<connection>
<GID>1962</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-888.5,357.5,-888.5</points>
<connection>
<GID>1976</GID>
<name>OUT</name></connection>
<intersection>-16.5 107</intersection>
<intersection>-8 4</intersection>
<intersection>33 108</intersection>
<intersection>40.5 16</intersection>
<intersection>81 109</intersection>
<intersection>88 23</intersection>
<intersection>130.5 110</intersection>
<intersection>138.5 31</intersection>
<intersection>178.5 111</intersection>
<intersection>187 55</intersection>
<intersection>236 112</intersection>
<intersection>245.5 56</intersection>
<intersection>291 113</intersection>
<intersection>299.5 66</intersection>
<intersection>348 114</intersection>
<intersection>357.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-8,-896,-8,-888.5</points>
<intersection>-896 5</intersection>
<intersection>-888.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-8,-896,-6.5,-896</points>
<connection>
<GID>1961</GID>
<name>IN_1</name></connection>
<intersection>-8 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>40.5,-897,40.5,-888.5</points>
<intersection>-897 21</intersection>
<intersection>-888.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>40.5,-897,42,-897</points>
<connection>
<GID>1963</GID>
<name>IN_1</name></connection>
<intersection>40.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>88,-896,88,-888.5</points>
<intersection>-896 53</intersection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>138.5,-896,138.5,-888.5</points>
<intersection>-896 115</intersection>
<intersection>-888.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>88,-896,88.5,-896</points>
<connection>
<GID>1965</GID>
<name>IN_1</name></connection>
<intersection>88 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>187,-895.5,187,-888.5</points>
<connection>
<GID>1969</GID>
<name>IN_1</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>245.5,-897.5,245.5,-888.5</points>
<connection>
<GID>1971</GID>
<name>IN_1</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>299.5,-896.5,299.5,-888.5</points>
<intersection>-896.5 118</intersection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>357.5,-897,357.5,-888.5</points>
<connection>
<GID>1975</GID>
<name>IN_1</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-16.5,-890.5,-16.5,-888.5</points>
<connection>
<GID>1960</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>33,-890.5,33,-888.5</points>
<connection>
<GID>1962</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>81,-890.5,81,-888.5</points>
<connection>
<GID>1964</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>130.5,-890.5,130.5,-888.5</points>
<connection>
<GID>1966</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>178.5,-890.5,178.5,-888.5</points>
<connection>
<GID>1968</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>236,-890.5,236,-888.5</points>
<connection>
<GID>1970</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>291,-890.5,291,-888.5</points>
<connection>
<GID>1972</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>348,-890.5,348,-888.5</points>
<connection>
<GID>1974</GID>
<name>clock</name></connection>
<intersection>-888.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>138.5,-896,139,-896</points>
<connection>
<GID>1967</GID>
<name>IN_1</name></connection>
<intersection>138.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>299,-896.5,299.5,-896.5</points>
<connection>
<GID>1973</GID>
<name>IN_1</name></connection>
<intersection>299.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-894,88.5,-887.5</points>
<connection>
<GID>1965</GID>
<name>IN_0</name></connection>
<intersection>-887.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>87,-887.5,88.5,-887.5</points>
<connection>
<GID>1964</GID>
<name>OUT_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-894,138,-887.5</points>
<intersection>-894 1</intersection>
<intersection>-887.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-894,139,-894</points>
<connection>
<GID>1967</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136.5,-887.5,138,-887.5</points>
<connection>
<GID>1966</GID>
<name>OUT_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-893.5,186.5,-887.5</points>
<intersection>-893.5 5</intersection>
<intersection>-887.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>184.5,-887.5,186.5,-887.5</points>
<connection>
<GID>1968</GID>
<name>OUT_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>186.5,-893.5,187,-893.5</points>
<connection>
<GID>1969</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-895.5,245,-887.5</points>
<intersection>-895.5 1</intersection>
<intersection>-887.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-895.5,245.5,-895.5</points>
<connection>
<GID>1971</GID>
<name>IN_0</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-887.5,245,-887.5</points>
<connection>
<GID>1970</GID>
<name>OUT_0</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-894.5,298.5,-887.5</points>
<intersection>-894.5 4</intersection>
<intersection>-887.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>297,-887.5,298.5,-887.5</points>
<connection>
<GID>1972</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>298.5,-894.5,299,-894.5</points>
<connection>
<GID>1973</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-895,357,-887.5</points>
<intersection>-895 1</intersection>
<intersection>-887.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-895,357.5,-895</points>
<connection>
<GID>1975</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-887.5,357,-887.5</points>
<connection>
<GID>1974</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-906.5,-9.5,-900</points>
<intersection>-906.5 1</intersection>
<intersection>-900 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-906.5,-7,-906.5</points>
<connection>
<GID>1978</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11,-900,-9.5,-900</points>
<connection>
<GID>1977</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-907.5,39.5,-900</points>
<intersection>-907.5 1</intersection>
<intersection>-900 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-907.5,41.5,-907.5</points>
<connection>
<GID>1980</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38.5,-900,39.5,-900</points>
<connection>
<GID>1979</GID>
<name>OUT_0</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42.5,-901,357,-901</points>
<connection>
<GID>1993</GID>
<name>OUT</name></connection>
<intersection>-17 107</intersection>
<intersection>-8.5 4</intersection>
<intersection>32.5 108</intersection>
<intersection>40 16</intersection>
<intersection>80.5 109</intersection>
<intersection>87.5 23</intersection>
<intersection>130 110</intersection>
<intersection>138 31</intersection>
<intersection>178 111</intersection>
<intersection>186.5 55</intersection>
<intersection>235.5 112</intersection>
<intersection>245 56</intersection>
<intersection>290.5 113</intersection>
<intersection>299 66</intersection>
<intersection>347.5 114</intersection>
<intersection>357 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-8.5,-908.5,-8.5,-901</points>
<intersection>-908.5 5</intersection>
<intersection>-901 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-8.5,-908.5,-7,-908.5</points>
<connection>
<GID>1978</GID>
<name>IN_1</name></connection>
<intersection>-8.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>40,-909.5,40,-901</points>
<intersection>-909.5 21</intersection>
<intersection>-901 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>40,-909.5,41.5,-909.5</points>
<connection>
<GID>1980</GID>
<name>IN_1</name></connection>
<intersection>40 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>87.5,-908.5,87.5,-901</points>
<intersection>-908.5 53</intersection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>138,-908.5,138,-901</points>
<intersection>-908.5 115</intersection>
<intersection>-901 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>87.5,-908.5,88,-908.5</points>
<connection>
<GID>1982</GID>
<name>IN_1</name></connection>
<intersection>87.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>186.5,-908,186.5,-901</points>
<connection>
<GID>1986</GID>
<name>IN_1</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>245,-910,245,-901</points>
<connection>
<GID>1988</GID>
<name>IN_1</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>299,-909,299,-901</points>
<intersection>-909 118</intersection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>357,-909.5,357,-901</points>
<connection>
<GID>1992</GID>
<name>IN_1</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-17,-903,-17,-901</points>
<connection>
<GID>1977</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>32.5,-903,32.5,-901</points>
<connection>
<GID>1979</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>80.5,-903,80.5,-901</points>
<connection>
<GID>1981</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>130,-903,130,-901</points>
<connection>
<GID>1983</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>178,-903,178,-901</points>
<connection>
<GID>1985</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>235.5,-903,235.5,-901</points>
<connection>
<GID>1987</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>290.5,-903,290.5,-901</points>
<connection>
<GID>1989</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>347.5,-903,347.5,-901</points>
<connection>
<GID>1991</GID>
<name>clock</name></connection>
<intersection>-901 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>138,-908.5,138.5,-908.5</points>
<connection>
<GID>1984</GID>
<name>IN_1</name></connection>
<intersection>138 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>298.5,-909,299,-909</points>
<connection>
<GID>1990</GID>
<name>IN_1</name></connection>
<intersection>299 66</intersection></hsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-906.5,88,-900</points>
<connection>
<GID>1982</GID>
<name>IN_0</name></connection>
<intersection>-900 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-900,88,-900</points>
<connection>
<GID>1981</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-906.5,137.5,-900</points>
<intersection>-906.5 1</intersection>
<intersection>-900 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-906.5,138.5,-906.5</points>
<connection>
<GID>1984</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136,-900,137.5,-900</points>
<connection>
<GID>1983</GID>
<name>OUT_0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-906,186,-900</points>
<intersection>-906 5</intersection>
<intersection>-900 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>184,-900,186,-900</points>
<connection>
<GID>1985</GID>
<name>OUT_0</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>186,-906,186.5,-906</points>
<connection>
<GID>1986</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-908,244.5,-900</points>
<intersection>-908 1</intersection>
<intersection>-900 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,-908,245,-908</points>
<connection>
<GID>1988</GID>
<name>IN_0</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241.5,-900,244.5,-900</points>
<connection>
<GID>1987</GID>
<name>OUT_0</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-907,298,-900</points>
<intersection>-907 4</intersection>
<intersection>-900 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>296.5,-900,298,-900</points>
<connection>
<GID>1989</GID>
<name>OUT_0</name></connection>
<intersection>298 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>298,-907,298.5,-907</points>
<connection>
<GID>1990</GID>
<name>IN_0</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,-907.5,356.5,-900</points>
<intersection>-907.5 1</intersection>
<intersection>-900 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356.5,-907.5,357,-907.5</points>
<connection>
<GID>1992</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353.5,-900,356.5,-900</points>
<connection>
<GID>1991</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-919.5,-10,-913</points>
<intersection>-919.5 1</intersection>
<intersection>-913 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-919.5,-7.5,-919.5</points>
<connection>
<GID>1995</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-913,-10,-913</points>
<connection>
<GID>1994</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-920.5,39,-913</points>
<intersection>-920.5 1</intersection>
<intersection>-913 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-920.5,41,-920.5</points>
<connection>
<GID>1997</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-913,39,-913</points>
<connection>
<GID>1996</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-914,356.5,-914</points>
<connection>
<GID>2010</GID>
<name>OUT</name></connection>
<intersection>-17.5 107</intersection>
<intersection>-9 4</intersection>
<intersection>32 108</intersection>
<intersection>39.5 16</intersection>
<intersection>80 109</intersection>
<intersection>87 23</intersection>
<intersection>129.5 110</intersection>
<intersection>137.5 31</intersection>
<intersection>177.5 111</intersection>
<intersection>186 55</intersection>
<intersection>235 112</intersection>
<intersection>244.5 56</intersection>
<intersection>290 113</intersection>
<intersection>298.5 66</intersection>
<intersection>347 114</intersection>
<intersection>356.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-9,-921.5,-9,-914</points>
<intersection>-921.5 5</intersection>
<intersection>-914 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-9,-921.5,-7.5,-921.5</points>
<connection>
<GID>1995</GID>
<name>IN_1</name></connection>
<intersection>-9 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>39.5,-922.5,39.5,-914</points>
<intersection>-922.5 21</intersection>
<intersection>-914 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>39.5,-922.5,41,-922.5</points>
<connection>
<GID>1997</GID>
<name>IN_1</name></connection>
<intersection>39.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>87,-921.5,87,-914</points>
<intersection>-921.5 53</intersection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>137.5,-921.5,137.5,-914</points>
<intersection>-921.5 115</intersection>
<intersection>-914 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>87,-921.5,87.5,-921.5</points>
<connection>
<GID>1999</GID>
<name>IN_1</name></connection>
<intersection>87 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>186,-921,186,-914</points>
<connection>
<GID>2003</GID>
<name>IN_1</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>244.5,-923,244.5,-914</points>
<connection>
<GID>2005</GID>
<name>IN_1</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>298.5,-922,298.5,-914</points>
<intersection>-922 118</intersection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>356.5,-922.5,356.5,-914</points>
<connection>
<GID>2009</GID>
<name>IN_1</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-17.5,-916,-17.5,-914</points>
<connection>
<GID>1994</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>32,-916,32,-914</points>
<connection>
<GID>1996</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>80,-916,80,-914</points>
<connection>
<GID>1998</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>129.5,-916,129.5,-914</points>
<connection>
<GID>2000</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>177.5,-916,177.5,-914</points>
<connection>
<GID>2002</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>235,-916,235,-914</points>
<connection>
<GID>2004</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>290,-916,290,-914</points>
<connection>
<GID>2006</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>347,-916,347,-914</points>
<connection>
<GID>2008</GID>
<name>clock</name></connection>
<intersection>-914 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>137.5,-921.5,138,-921.5</points>
<connection>
<GID>2001</GID>
<name>IN_1</name></connection>
<intersection>137.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>298,-922,298.5,-922</points>
<connection>
<GID>2007</GID>
<name>IN_1</name></connection>
<intersection>298.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-919.5,87.5,-913</points>
<connection>
<GID>1999</GID>
<name>IN_0</name></connection>
<intersection>-913 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86,-913,87.5,-913</points>
<connection>
<GID>1998</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-919.5,137,-913</points>
<intersection>-919.5 1</intersection>
<intersection>-913 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-919.5,138,-919.5</points>
<connection>
<GID>2001</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>135.5,-913,137,-913</points>
<connection>
<GID>2000</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-919,185.5,-913</points>
<intersection>-919 5</intersection>
<intersection>-913 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>183.5,-913,185.5,-913</points>
<connection>
<GID>2002</GID>
<name>OUT_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>185.5,-919,186,-919</points>
<connection>
<GID>2003</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-921,244,-913</points>
<intersection>-921 1</intersection>
<intersection>-913 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-921,244.5,-921</points>
<connection>
<GID>2005</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241,-913,244,-913</points>
<connection>
<GID>2004</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-920,297.5,-913</points>
<intersection>-920 4</intersection>
<intersection>-913 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>296,-913,297.5,-913</points>
<connection>
<GID>2006</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>297.5,-920,298,-920</points>
<connection>
<GID>2007</GID>
<name>IN_0</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-920.5,356,-913</points>
<intersection>-920.5 1</intersection>
<intersection>-913 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-920.5,356.5,-920.5</points>
<connection>
<GID>2009</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-913,356,-913</points>
<connection>
<GID>2008</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-934.5,-10,-928</points>
<intersection>-934.5 1</intersection>
<intersection>-928 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-934.5,-7.5,-934.5</points>
<connection>
<GID>1876</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-928,-10,-928</points>
<connection>
<GID>1875</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-935.5,39,-928</points>
<intersection>-935.5 1</intersection>
<intersection>-928 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-935.5,41,-935.5</points>
<connection>
<GID>1878</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-928,39,-928</points>
<connection>
<GID>1877</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-929,356.5,-929</points>
<connection>
<GID>1891</GID>
<name>OUT</name></connection>
<intersection>-17.5 107</intersection>
<intersection>-9 4</intersection>
<intersection>32 108</intersection>
<intersection>39.5 16</intersection>
<intersection>80 109</intersection>
<intersection>87 23</intersection>
<intersection>129.5 110</intersection>
<intersection>137.5 31</intersection>
<intersection>177.5 111</intersection>
<intersection>186 55</intersection>
<intersection>235 112</intersection>
<intersection>244.5 56</intersection>
<intersection>290 113</intersection>
<intersection>298.5 66</intersection>
<intersection>347 114</intersection>
<intersection>356.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-9,-936.5,-9,-929</points>
<intersection>-936.5 5</intersection>
<intersection>-929 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-9,-936.5,-7.5,-936.5</points>
<connection>
<GID>1876</GID>
<name>IN_1</name></connection>
<intersection>-9 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>39.5,-937.5,39.5,-929</points>
<intersection>-937.5 21</intersection>
<intersection>-929 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>39.5,-937.5,41,-937.5</points>
<connection>
<GID>1878</GID>
<name>IN_1</name></connection>
<intersection>39.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>87,-936.5,87,-929</points>
<intersection>-936.5 53</intersection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>137.5,-936.5,137.5,-929</points>
<intersection>-936.5 115</intersection>
<intersection>-929 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>87,-936.5,87.5,-936.5</points>
<connection>
<GID>1880</GID>
<name>IN_1</name></connection>
<intersection>87 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>186,-936,186,-929</points>
<connection>
<GID>1884</GID>
<name>IN_1</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>244.5,-938,244.5,-929</points>
<connection>
<GID>1886</GID>
<name>IN_1</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>298.5,-937,298.5,-929</points>
<intersection>-937 118</intersection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>356.5,-937.5,356.5,-929</points>
<connection>
<GID>1890</GID>
<name>IN_1</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-17.5,-931,-17.5,-929</points>
<connection>
<GID>1875</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>32,-931,32,-929</points>
<connection>
<GID>1877</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>80,-931,80,-929</points>
<connection>
<GID>1879</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>129.5,-931,129.5,-929</points>
<connection>
<GID>1881</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>177.5,-931,177.5,-929</points>
<connection>
<GID>1883</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>235,-931,235,-929</points>
<connection>
<GID>1885</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>290,-931,290,-929</points>
<connection>
<GID>1887</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>347,-931,347,-929</points>
<connection>
<GID>1889</GID>
<name>clock</name></connection>
<intersection>-929 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>137.5,-936.5,138,-936.5</points>
<connection>
<GID>1882</GID>
<name>IN_1</name></connection>
<intersection>137.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>298,-937,298.5,-937</points>
<connection>
<GID>1888</GID>
<name>IN_1</name></connection>
<intersection>298.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-934.5,87.5,-928</points>
<connection>
<GID>1880</GID>
<name>IN_0</name></connection>
<intersection>-928 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86,-928,87.5,-928</points>
<connection>
<GID>1879</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-934.5,137,-928</points>
<intersection>-934.5 1</intersection>
<intersection>-928 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-934.5,138,-934.5</points>
<connection>
<GID>1882</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>135.5,-928,137,-928</points>
<connection>
<GID>1881</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-934,185.5,-928</points>
<intersection>-934 5</intersection>
<intersection>-928 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>183.5,-928,185.5,-928</points>
<connection>
<GID>1883</GID>
<name>OUT_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>185.5,-934,186,-934</points>
<connection>
<GID>1884</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-936,244,-928</points>
<intersection>-936 1</intersection>
<intersection>-928 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-936,244.5,-936</points>
<connection>
<GID>1886</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241,-928,244,-928</points>
<connection>
<GID>1885</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-935,297.5,-928</points>
<intersection>-935 4</intersection>
<intersection>-928 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>296,-928,297.5,-928</points>
<connection>
<GID>1887</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>297.5,-935,298,-935</points>
<connection>
<GID>1888</GID>
<name>IN_0</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-935.5,356,-928</points>
<intersection>-935.5 1</intersection>
<intersection>-928 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-935.5,356.5,-935.5</points>
<connection>
<GID>1890</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-928,356,-928</points>
<connection>
<GID>1889</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-948.5,-10,-942</points>
<intersection>-948.5 1</intersection>
<intersection>-942 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-948.5,-7.5,-948.5</points>
<connection>
<GID>1893</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-942,-10,-942</points>
<connection>
<GID>1892</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-949.5,39,-942</points>
<intersection>-949.5 1</intersection>
<intersection>-942 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-949.5,41,-949.5</points>
<connection>
<GID>1895</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-942,39,-942</points>
<connection>
<GID>1894</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-943,356.5,-943</points>
<connection>
<GID>1908</GID>
<name>OUT</name></connection>
<intersection>-17.5 107</intersection>
<intersection>-9 4</intersection>
<intersection>32 108</intersection>
<intersection>39.5 16</intersection>
<intersection>80 109</intersection>
<intersection>87 23</intersection>
<intersection>129.5 110</intersection>
<intersection>137.5 31</intersection>
<intersection>177.5 111</intersection>
<intersection>186 55</intersection>
<intersection>235 112</intersection>
<intersection>244.5 56</intersection>
<intersection>290 113</intersection>
<intersection>298.5 66</intersection>
<intersection>347 114</intersection>
<intersection>356.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-9,-950.5,-9,-943</points>
<intersection>-950.5 5</intersection>
<intersection>-943 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-9,-950.5,-7.5,-950.5</points>
<connection>
<GID>1893</GID>
<name>IN_1</name></connection>
<intersection>-9 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>39.5,-951.5,39.5,-943</points>
<intersection>-951.5 21</intersection>
<intersection>-943 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>39.5,-951.5,41,-951.5</points>
<connection>
<GID>1895</GID>
<name>IN_1</name></connection>
<intersection>39.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>87,-950.5,87,-943</points>
<intersection>-950.5 53</intersection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>137.5,-950.5,137.5,-943</points>
<intersection>-950.5 115</intersection>
<intersection>-943 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>87,-950.5,87.5,-950.5</points>
<connection>
<GID>1897</GID>
<name>IN_1</name></connection>
<intersection>87 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>186,-950,186,-943</points>
<connection>
<GID>1901</GID>
<name>IN_1</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>244.5,-952,244.5,-943</points>
<connection>
<GID>1903</GID>
<name>IN_1</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>298.5,-951,298.5,-943</points>
<intersection>-951 118</intersection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>356.5,-951.5,356.5,-943</points>
<connection>
<GID>1907</GID>
<name>IN_1</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-17.5,-945,-17.5,-943</points>
<connection>
<GID>1892</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>32,-945,32,-943</points>
<connection>
<GID>1894</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>80,-945,80,-943</points>
<connection>
<GID>1896</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>129.5,-945,129.5,-943</points>
<connection>
<GID>1898</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>177.5,-945,177.5,-943</points>
<connection>
<GID>1900</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>235,-945,235,-943</points>
<connection>
<GID>1902</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>290,-945,290,-943</points>
<connection>
<GID>1904</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>347,-945,347,-943</points>
<connection>
<GID>1906</GID>
<name>clock</name></connection>
<intersection>-943 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>137.5,-950.5,138,-950.5</points>
<connection>
<GID>1899</GID>
<name>IN_1</name></connection>
<intersection>137.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>298,-951,298.5,-951</points>
<connection>
<GID>1905</GID>
<name>IN_1</name></connection>
<intersection>298.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-948.5,87.5,-942</points>
<connection>
<GID>1897</GID>
<name>IN_0</name></connection>
<intersection>-942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86,-942,87.5,-942</points>
<connection>
<GID>1896</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-948.5,137,-942</points>
<intersection>-948.5 1</intersection>
<intersection>-942 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-948.5,138,-948.5</points>
<connection>
<GID>1899</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>135.5,-942,137,-942</points>
<connection>
<GID>1898</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-948,185.5,-942</points>
<intersection>-948 5</intersection>
<intersection>-942 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>183.5,-942,185.5,-942</points>
<connection>
<GID>1900</GID>
<name>OUT_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>185.5,-948,186,-948</points>
<connection>
<GID>1901</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-950,244,-942</points>
<intersection>-950 1</intersection>
<intersection>-942 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-950,244.5,-950</points>
<connection>
<GID>1903</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241,-942,244,-942</points>
<connection>
<GID>1902</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-949,297.5,-942</points>
<intersection>-949 4</intersection>
<intersection>-942 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>296,-942,297.5,-942</points>
<connection>
<GID>1904</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>297.5,-949,298,-949</points>
<connection>
<GID>1905</GID>
<name>IN_0</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-949.5,356,-942</points>
<intersection>-949.5 1</intersection>
<intersection>-942 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-949.5,356.5,-949.5</points>
<connection>
<GID>1907</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-942,356,-942</points>
<connection>
<GID>1906</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment></shape></wire>
<wire>
<ID>1141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-966,-10.5,-959.5</points>
<intersection>-966 1</intersection>
<intersection>-959.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10.5,-966,-8,-966</points>
<connection>
<GID>1910</GID>
<name>IN_0</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12,-959.5,-10.5,-959.5</points>
<connection>
<GID>1909</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-967,38.5,-959.5</points>
<intersection>-967 1</intersection>
<intersection>-959.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-967,40.5,-967</points>
<connection>
<GID>1912</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>37.5,-959.5,38.5,-959.5</points>
<connection>
<GID>1911</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43.5,-960.5,356,-960.5</points>
<connection>
<GID>1925</GID>
<name>OUT</name></connection>
<intersection>-18 107</intersection>
<intersection>-9.5 4</intersection>
<intersection>31.5 108</intersection>
<intersection>39 16</intersection>
<intersection>79.5 109</intersection>
<intersection>86.5 23</intersection>
<intersection>129 110</intersection>
<intersection>137 31</intersection>
<intersection>177 111</intersection>
<intersection>185.5 55</intersection>
<intersection>234.5 112</intersection>
<intersection>244 56</intersection>
<intersection>289.5 113</intersection>
<intersection>298 66</intersection>
<intersection>346.5 114</intersection>
<intersection>356 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-9.5,-968,-9.5,-960.5</points>
<intersection>-968 5</intersection>
<intersection>-960.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-9.5,-968,-8,-968</points>
<connection>
<GID>1910</GID>
<name>IN_1</name></connection>
<intersection>-9.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>39,-969,39,-960.5</points>
<intersection>-969 21</intersection>
<intersection>-960.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>39,-969,40.5,-969</points>
<connection>
<GID>1912</GID>
<name>IN_1</name></connection>
<intersection>39 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>86.5,-968,86.5,-960.5</points>
<intersection>-968 53</intersection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>137,-968,137,-960.5</points>
<intersection>-968 115</intersection>
<intersection>-960.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>86.5,-968,87,-968</points>
<connection>
<GID>1914</GID>
<name>IN_1</name></connection>
<intersection>86.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>185.5,-967.5,185.5,-960.5</points>
<connection>
<GID>1918</GID>
<name>IN_1</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>244,-969.5,244,-960.5</points>
<connection>
<GID>1920</GID>
<name>IN_1</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>298,-968.5,298,-960.5</points>
<intersection>-968.5 118</intersection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>356,-969,356,-960.5</points>
<connection>
<GID>1924</GID>
<name>IN_1</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-18,-962.5,-18,-960.5</points>
<connection>
<GID>1909</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>31.5,-962.5,31.5,-960.5</points>
<connection>
<GID>1911</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>79.5,-962.5,79.5,-960.5</points>
<connection>
<GID>1913</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>129,-962.5,129,-960.5</points>
<connection>
<GID>1915</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>177,-962.5,177,-960.5</points>
<connection>
<GID>1917</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>234.5,-962.5,234.5,-960.5</points>
<connection>
<GID>1919</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>289.5,-962.5,289.5,-960.5</points>
<connection>
<GID>1921</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>346.5,-962.5,346.5,-960.5</points>
<connection>
<GID>1923</GID>
<name>clock</name></connection>
<intersection>-960.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>137,-968,137.5,-968</points>
<connection>
<GID>1916</GID>
<name>IN_1</name></connection>
<intersection>137 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>297.5,-968.5,298,-968.5</points>
<connection>
<GID>1922</GID>
<name>IN_1</name></connection>
<intersection>298 66</intersection></hsegment></shape></wire>
<wire>
<ID>1144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-966,87,-959.5</points>
<connection>
<GID>1914</GID>
<name>IN_0</name></connection>
<intersection>-959.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>85.5,-959.5,87,-959.5</points>
<connection>
<GID>1913</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>1145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-966,136.5,-959.5</points>
<intersection>-966 1</intersection>
<intersection>-959.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-966,137.5,-966</points>
<connection>
<GID>1916</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>135,-959.5,136.5,-959.5</points>
<connection>
<GID>1915</GID>
<name>OUT_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-965.5,185,-959.5</points>
<intersection>-965.5 5</intersection>
<intersection>-959.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>183,-959.5,185,-959.5</points>
<connection>
<GID>1917</GID>
<name>OUT_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>185,-965.5,185.5,-965.5</points>
<connection>
<GID>1918</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>1147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243.5,-967.5,243.5,-959.5</points>
<intersection>-967.5 1</intersection>
<intersection>-959.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243.5,-967.5,244,-967.5</points>
<connection>
<GID>1920</GID>
<name>IN_0</name></connection>
<intersection>243.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>240.5,-959.5,243.5,-959.5</points>
<connection>
<GID>1919</GID>
<name>OUT_0</name></connection>
<intersection>243.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297,-966.5,297,-959.5</points>
<intersection>-966.5 4</intersection>
<intersection>-959.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>295.5,-959.5,297,-959.5</points>
<connection>
<GID>1921</GID>
<name>OUT_0</name></connection>
<intersection>297 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>297,-966.5,297.5,-966.5</points>
<connection>
<GID>1922</GID>
<name>IN_0</name></connection>
<intersection>297 0</intersection></hsegment></shape></wire>
<wire>
<ID>1149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355.5,-967,355.5,-959.5</points>
<intersection>-967 1</intersection>
<intersection>-959.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,-967,356,-967</points>
<connection>
<GID>1924</GID>
<name>IN_0</name></connection>
<intersection>355.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352.5,-959.5,355.5,-959.5</points>
<connection>
<GID>1923</GID>
<name>OUT_0</name></connection>
<intersection>355.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-917,-60,-860</points>
<intersection>-917 2</intersection>
<intersection>-860 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,-860,-48,-860</points>
<connection>
<GID>1942</GID>
<name>IN_0</name></connection>
<intersection>-60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-917,-60,-917</points>
<connection>
<GID>469</GID>
<name>OUT_7</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>1151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,-918,-59,-873</points>
<intersection>-918 2</intersection>
<intersection>-873 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59,-873,-48,-873</points>
<connection>
<GID>1959</GID>
<name>IN_0</name></connection>
<intersection>-59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-918,-59,-918</points>
<connection>
<GID>469</GID>
<name>OUT_6</name></connection>
<intersection>-59 0</intersection></hsegment></shape></wire>
<wire>
<ID>1152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-919,-58,-887.5</points>
<intersection>-919 2</intersection>
<intersection>-887.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-887.5,-48,-887.5</points>
<connection>
<GID>1976</GID>
<name>IN_0</name></connection>
<intersection>-58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-919,-58,-919</points>
<connection>
<GID>469</GID>
<name>OUT_5</name></connection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>1153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-920,-57,-900</points>
<intersection>-920 2</intersection>
<intersection>-900 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,-900,-48.5,-900</points>
<connection>
<GID>1993</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-920,-57,-920</points>
<connection>
<GID>469</GID>
<name>OUT_4</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>1154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-921,-56,-913</points>
<intersection>-921 2</intersection>
<intersection>-913 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-913,-49,-913</points>
<connection>
<GID>2010</GID>
<name>IN_0</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-921,-56,-921</points>
<connection>
<GID>469</GID>
<name>OUT_3</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>1155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-928,-56,-922</points>
<intersection>-928 1</intersection>
<intersection>-922 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-928,-49,-928</points>
<connection>
<GID>1891</GID>
<name>IN_0</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-922,-56,-922</points>
<connection>
<GID>469</GID>
<name>OUT_2</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>1156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-942,-57,-923</points>
<intersection>-942 1</intersection>
<intersection>-923 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,-942,-49,-942</points>
<connection>
<GID>1908</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-923,-57,-923</points>
<connection>
<GID>469</GID>
<name>OUT_1</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>1157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-959.5,-58.5,-924</points>
<intersection>-959.5 1</intersection>
<intersection>-924 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,-959.5,-49.5,-959.5</points>
<connection>
<GID>1925</GID>
<name>IN_0</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-924,-58.5,-924</points>
<connection>
<GID>469</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-1192,-13,-1185.5</points>
<intersection>-1192 1</intersection>
<intersection>-1185.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-1192,-10.5,-1192</points>
<connection>
<GID>2063</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14.5,-1185.5,-13,-1185.5</points>
<connection>
<GID>2062</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>1159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-1193,36,-1185.5</points>
<intersection>-1193 1</intersection>
<intersection>-1185.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-1193,38,-1193</points>
<connection>
<GID>2065</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-1185.5,36,-1185.5</points>
<connection>
<GID>2064</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-1186.5,353.5,-1186.5</points>
<connection>
<GID>2078</GID>
<name>OUT</name></connection>
<intersection>-20.5 107</intersection>
<intersection>-12 4</intersection>
<intersection>29 108</intersection>
<intersection>36.5 16</intersection>
<intersection>77 109</intersection>
<intersection>84 23</intersection>
<intersection>126.5 110</intersection>
<intersection>134.5 31</intersection>
<intersection>174.5 111</intersection>
<intersection>183 55</intersection>
<intersection>232 112</intersection>
<intersection>241.5 56</intersection>
<intersection>287 113</intersection>
<intersection>295.5 66</intersection>
<intersection>344 114</intersection>
<intersection>353.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-1194,-12,-1186.5</points>
<intersection>-1194 5</intersection>
<intersection>-1186.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-1194,-10.5,-1194</points>
<connection>
<GID>2063</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36.5,-1195,36.5,-1186.5</points>
<intersection>-1195 21</intersection>
<intersection>-1186.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36.5,-1195,38,-1195</points>
<connection>
<GID>2065</GID>
<name>IN_1</name></connection>
<intersection>36.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84,-1194,84,-1186.5</points>
<intersection>-1194 53</intersection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134.5,-1194,134.5,-1186.5</points>
<intersection>-1194 115</intersection>
<intersection>-1186.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84,-1194,84.5,-1194</points>
<connection>
<GID>2067</GID>
<name>IN_1</name></connection>
<intersection>84 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183,-1193.5,183,-1186.5</points>
<connection>
<GID>2071</GID>
<name>IN_1</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241.5,-1195.5,241.5,-1186.5</points>
<connection>
<GID>2073</GID>
<name>IN_1</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295.5,-1194.5,295.5,-1186.5</points>
<intersection>-1194.5 118</intersection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353.5,-1195,353.5,-1186.5</points>
<connection>
<GID>2077</GID>
<name>IN_1</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20.5,-1188.5,-20.5,-1186.5</points>
<connection>
<GID>2062</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29,-1188.5,29,-1186.5</points>
<connection>
<GID>2064</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77,-1188.5,77,-1186.5</points>
<connection>
<GID>2066</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126.5,-1188.5,126.5,-1186.5</points>
<connection>
<GID>2068</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174.5,-1188.5,174.5,-1186.5</points>
<connection>
<GID>2070</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232,-1188.5,232,-1186.5</points>
<connection>
<GID>2072</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287,-1188.5,287,-1186.5</points>
<connection>
<GID>2074</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344,-1188.5,344,-1186.5</points>
<connection>
<GID>2076</GID>
<name>clock</name></connection>
<intersection>-1186.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134.5,-1194,135,-1194</points>
<connection>
<GID>2069</GID>
<name>IN_1</name></connection>
<intersection>134.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295,-1194.5,295.5,-1194.5</points>
<connection>
<GID>2075</GID>
<name>IN_1</name></connection>
<intersection>295.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-1192,84.5,-1185.5</points>
<connection>
<GID>2067</GID>
<name>IN_0</name></connection>
<intersection>-1185.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83,-1185.5,84.5,-1185.5</points>
<connection>
<GID>2066</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-1192,134,-1185.5</points>
<intersection>-1192 1</intersection>
<intersection>-1185.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-1192,135,-1192</points>
<connection>
<GID>2069</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-1185.5,134,-1185.5</points>
<connection>
<GID>2068</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-1191.5,182.5,-1185.5</points>
<intersection>-1191.5 5</intersection>
<intersection>-1185.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180.5,-1185.5,182.5,-1185.5</points>
<connection>
<GID>2070</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-1191.5,183,-1191.5</points>
<connection>
<GID>2071</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-1193.5,241,-1185.5</points>
<intersection>-1193.5 1</intersection>
<intersection>-1185.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-1193.5,241.5,-1193.5</points>
<connection>
<GID>2073</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-1185.5,241,-1185.5</points>
<connection>
<GID>2072</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>1165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-1192.5,294.5,-1185.5</points>
<intersection>-1192.5 4</intersection>
<intersection>-1185.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-1185.5,294.5,-1185.5</points>
<connection>
<GID>2074</GID>
<name>OUT_0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-1192.5,295,-1192.5</points>
<connection>
<GID>2075</GID>
<name>IN_0</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-1193,353,-1185.5</points>
<intersection>-1193 1</intersection>
<intersection>-1185.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-1193,353.5,-1193</points>
<connection>
<GID>2077</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-1185.5,353,-1185.5</points>
<connection>
<GID>2076</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment></shape></wire>
<wire>
<ID>1167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-1205,-13,-1198.5</points>
<intersection>-1205 1</intersection>
<intersection>-1198.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-1205,-10.5,-1205</points>
<connection>
<GID>2080</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14.5,-1198.5,-13,-1198.5</points>
<connection>
<GID>2079</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>1168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-1206,36,-1198.5</points>
<intersection>-1206 1</intersection>
<intersection>-1198.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-1206,38,-1206</points>
<connection>
<GID>2082</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-1198.5,36,-1198.5</points>
<connection>
<GID>2081</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-1199.5,353.5,-1199.5</points>
<connection>
<GID>2095</GID>
<name>OUT</name></connection>
<intersection>-20.5 107</intersection>
<intersection>-12 4</intersection>
<intersection>29 108</intersection>
<intersection>36.5 16</intersection>
<intersection>77 109</intersection>
<intersection>84 23</intersection>
<intersection>126.5 110</intersection>
<intersection>134.5 31</intersection>
<intersection>174.5 111</intersection>
<intersection>183 55</intersection>
<intersection>232 112</intersection>
<intersection>241.5 56</intersection>
<intersection>287 113</intersection>
<intersection>295.5 66</intersection>
<intersection>344 114</intersection>
<intersection>353.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-1207,-12,-1199.5</points>
<intersection>-1207 5</intersection>
<intersection>-1199.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-1207,-10.5,-1207</points>
<connection>
<GID>2080</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36.5,-1208,36.5,-1199.5</points>
<intersection>-1208 21</intersection>
<intersection>-1199.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36.5,-1208,38,-1208</points>
<connection>
<GID>2082</GID>
<name>IN_1</name></connection>
<intersection>36.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84,-1207,84,-1199.5</points>
<intersection>-1207 53</intersection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134.5,-1207,134.5,-1199.5</points>
<intersection>-1207 115</intersection>
<intersection>-1199.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84,-1207,84.5,-1207</points>
<connection>
<GID>2084</GID>
<name>IN_1</name></connection>
<intersection>84 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183,-1206.5,183,-1199.5</points>
<connection>
<GID>2088</GID>
<name>IN_1</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241.5,-1208.5,241.5,-1199.5</points>
<connection>
<GID>2090</GID>
<name>IN_1</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295.5,-1207.5,295.5,-1199.5</points>
<intersection>-1207.5 118</intersection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353.5,-1208,353.5,-1199.5</points>
<connection>
<GID>2094</GID>
<name>IN_1</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20.5,-1201.5,-20.5,-1199.5</points>
<connection>
<GID>2079</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29,-1201.5,29,-1199.5</points>
<connection>
<GID>2081</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77,-1201.5,77,-1199.5</points>
<connection>
<GID>2083</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126.5,-1201.5,126.5,-1199.5</points>
<connection>
<GID>2085</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174.5,-1201.5,174.5,-1199.5</points>
<connection>
<GID>2087</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232,-1201.5,232,-1199.5</points>
<connection>
<GID>2089</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287,-1201.5,287,-1199.5</points>
<connection>
<GID>2091</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344,-1201.5,344,-1199.5</points>
<connection>
<GID>2093</GID>
<name>clock</name></connection>
<intersection>-1199.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134.5,-1207,135,-1207</points>
<connection>
<GID>2086</GID>
<name>IN_1</name></connection>
<intersection>134.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295,-1207.5,295.5,-1207.5</points>
<connection>
<GID>2092</GID>
<name>IN_1</name></connection>
<intersection>295.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-1205,84.5,-1198.5</points>
<connection>
<GID>2084</GID>
<name>IN_0</name></connection>
<intersection>-1198.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83,-1198.5,84.5,-1198.5</points>
<connection>
<GID>2083</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-1205,134,-1198.5</points>
<intersection>-1205 1</intersection>
<intersection>-1198.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-1205,135,-1205</points>
<connection>
<GID>2086</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-1198.5,134,-1198.5</points>
<connection>
<GID>2085</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-1204.5,182.5,-1198.5</points>
<intersection>-1204.5 5</intersection>
<intersection>-1198.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180.5,-1198.5,182.5,-1198.5</points>
<connection>
<GID>2087</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-1204.5,183,-1204.5</points>
<connection>
<GID>2088</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-1206.5,241,-1198.5</points>
<intersection>-1206.5 1</intersection>
<intersection>-1198.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-1206.5,241.5,-1206.5</points>
<connection>
<GID>2090</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-1198.5,241,-1198.5</points>
<connection>
<GID>2089</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>1174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-1205.5,294.5,-1198.5</points>
<intersection>-1205.5 4</intersection>
<intersection>-1198.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-1198.5,294.5,-1198.5</points>
<connection>
<GID>2091</GID>
<name>OUT_0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-1205.5,295,-1205.5</points>
<connection>
<GID>2092</GID>
<name>IN_0</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-1206,353,-1198.5</points>
<intersection>-1206 1</intersection>
<intersection>-1198.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-1206,353.5,-1206</points>
<connection>
<GID>2094</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-1198.5,353,-1198.5</points>
<connection>
<GID>2093</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment></shape></wire>
<wire>
<ID>1176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-1219.5,-13,-1213</points>
<intersection>-1219.5 1</intersection>
<intersection>-1213 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-1219.5,-10.5,-1219.5</points>
<connection>
<GID>2097</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14.5,-1213,-13,-1213</points>
<connection>
<GID>2096</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>1177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-1220.5,36,-1213</points>
<intersection>-1220.5 1</intersection>
<intersection>-1213 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-1220.5,38,-1220.5</points>
<connection>
<GID>2099</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-1213,36,-1213</points>
<connection>
<GID>2098</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-1214,353.5,-1214</points>
<connection>
<GID>2112</GID>
<name>OUT</name></connection>
<intersection>-20.5 107</intersection>
<intersection>-12 4</intersection>
<intersection>29 108</intersection>
<intersection>36.5 16</intersection>
<intersection>77 109</intersection>
<intersection>84 23</intersection>
<intersection>126.5 110</intersection>
<intersection>134.5 31</intersection>
<intersection>174.5 111</intersection>
<intersection>183 55</intersection>
<intersection>232 112</intersection>
<intersection>241.5 56</intersection>
<intersection>287 113</intersection>
<intersection>295.5 66</intersection>
<intersection>344 114</intersection>
<intersection>353.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-1221.5,-12,-1214</points>
<intersection>-1221.5 5</intersection>
<intersection>-1214 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12,-1221.5,-10.5,-1221.5</points>
<connection>
<GID>2097</GID>
<name>IN_1</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36.5,-1222.5,36.5,-1214</points>
<intersection>-1222.5 21</intersection>
<intersection>-1214 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36.5,-1222.5,38,-1222.5</points>
<connection>
<GID>2099</GID>
<name>IN_1</name></connection>
<intersection>36.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84,-1221.5,84,-1214</points>
<intersection>-1221.5 53</intersection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134.5,-1221.5,134.5,-1214</points>
<intersection>-1221.5 115</intersection>
<intersection>-1214 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84,-1221.5,84.5,-1221.5</points>
<connection>
<GID>2101</GID>
<name>IN_1</name></connection>
<intersection>84 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183,-1221,183,-1214</points>
<connection>
<GID>2105</GID>
<name>IN_1</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241.5,-1223,241.5,-1214</points>
<connection>
<GID>2107</GID>
<name>IN_1</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295.5,-1222,295.5,-1214</points>
<intersection>-1222 118</intersection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353.5,-1222.5,353.5,-1214</points>
<connection>
<GID>2111</GID>
<name>IN_1</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20.5,-1216,-20.5,-1214</points>
<connection>
<GID>2096</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29,-1216,29,-1214</points>
<connection>
<GID>2098</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77,-1216,77,-1214</points>
<connection>
<GID>2100</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126.5,-1216,126.5,-1214</points>
<connection>
<GID>2102</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174.5,-1216,174.5,-1214</points>
<connection>
<GID>2104</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232,-1216,232,-1214</points>
<connection>
<GID>2106</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287,-1216,287,-1214</points>
<connection>
<GID>2108</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344,-1216,344,-1214</points>
<connection>
<GID>2110</GID>
<name>clock</name></connection>
<intersection>-1214 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134.5,-1221.5,135,-1221.5</points>
<connection>
<GID>2103</GID>
<name>IN_1</name></connection>
<intersection>134.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295,-1222,295.5,-1222</points>
<connection>
<GID>2109</GID>
<name>IN_1</name></connection>
<intersection>295.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-1219.5,84.5,-1213</points>
<connection>
<GID>2101</GID>
<name>IN_0</name></connection>
<intersection>-1213 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>83,-1213,84.5,-1213</points>
<connection>
<GID>2100</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-1219.5,134,-1213</points>
<intersection>-1219.5 1</intersection>
<intersection>-1213 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-1219.5,135,-1219.5</points>
<connection>
<GID>2103</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-1213,134,-1213</points>
<connection>
<GID>2102</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-1219,182.5,-1213</points>
<intersection>-1219 5</intersection>
<intersection>-1213 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180.5,-1213,182.5,-1213</points>
<connection>
<GID>2104</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-1219,183,-1219</points>
<connection>
<GID>2105</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-1221,241,-1213</points>
<intersection>-1221 1</intersection>
<intersection>-1213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-1221,241.5,-1221</points>
<connection>
<GID>2107</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,-1213,241,-1213</points>
<connection>
<GID>2106</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>1183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-1220,294.5,-1213</points>
<intersection>-1220 4</intersection>
<intersection>-1213 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>293,-1213,294.5,-1213</points>
<connection>
<GID>2108</GID>
<name>OUT_0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-1220,295,-1220</points>
<connection>
<GID>2109</GID>
<name>IN_0</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-1220.5,353,-1213</points>
<intersection>-1220.5 1</intersection>
<intersection>-1213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-1220.5,353.5,-1220.5</points>
<connection>
<GID>2111</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-1213,353,-1213</points>
<connection>
<GID>2110</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment></shape></wire>
<wire>
<ID>1185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-1232,-13.5,-1225.5</points>
<intersection>-1232 1</intersection>
<intersection>-1225.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-1232,-11,-1232</points>
<connection>
<GID>2114</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15,-1225.5,-13.5,-1225.5</points>
<connection>
<GID>2113</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-1233,35.5,-1225.5</points>
<intersection>-1233 1</intersection>
<intersection>-1225.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-1233,37.5,-1233</points>
<connection>
<GID>2116</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34.5,-1225.5,35.5,-1225.5</points>
<connection>
<GID>2115</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46.5,-1226.5,353,-1226.5</points>
<connection>
<GID>2129</GID>
<name>OUT</name></connection>
<intersection>-21 107</intersection>
<intersection>-12.5 4</intersection>
<intersection>28.5 108</intersection>
<intersection>36 16</intersection>
<intersection>76.5 109</intersection>
<intersection>83.5 23</intersection>
<intersection>126 110</intersection>
<intersection>134 31</intersection>
<intersection>174 111</intersection>
<intersection>182.5 55</intersection>
<intersection>231.5 112</intersection>
<intersection>241 56</intersection>
<intersection>286.5 113</intersection>
<intersection>295 66</intersection>
<intersection>343.5 114</intersection>
<intersection>353 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12.5,-1234,-12.5,-1226.5</points>
<intersection>-1234 5</intersection>
<intersection>-1226.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,-1234,-11,-1234</points>
<connection>
<GID>2114</GID>
<name>IN_1</name></connection>
<intersection>-12.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>36,-1235,36,-1226.5</points>
<intersection>-1235 21</intersection>
<intersection>-1226.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>36,-1235,37.5,-1235</points>
<connection>
<GID>2116</GID>
<name>IN_1</name></connection>
<intersection>36 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83.5,-1234,83.5,-1226.5</points>
<intersection>-1234 53</intersection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>134,-1234,134,-1226.5</points>
<intersection>-1234 115</intersection>
<intersection>-1226.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83.5,-1234,84,-1234</points>
<connection>
<GID>2118</GID>
<name>IN_1</name></connection>
<intersection>83.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182.5,-1233.5,182.5,-1226.5</points>
<connection>
<GID>2122</GID>
<name>IN_1</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>241,-1235.5,241,-1226.5</points>
<connection>
<GID>2124</GID>
<name>IN_1</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>295,-1234.5,295,-1226.5</points>
<intersection>-1234.5 118</intersection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>353,-1235,353,-1226.5</points>
<connection>
<GID>2128</GID>
<name>IN_1</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21,-1228.5,-21,-1226.5</points>
<connection>
<GID>2113</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28.5,-1228.5,28.5,-1226.5</points>
<connection>
<GID>2115</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76.5,-1228.5,76.5,-1226.5</points>
<connection>
<GID>2117</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>126,-1228.5,126,-1226.5</points>
<connection>
<GID>2119</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>174,-1228.5,174,-1226.5</points>
<connection>
<GID>2121</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231.5,-1228.5,231.5,-1226.5</points>
<connection>
<GID>2123</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286.5,-1228.5,286.5,-1226.5</points>
<connection>
<GID>2125</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343.5,-1228.5,343.5,-1226.5</points>
<connection>
<GID>2127</GID>
<name>clock</name></connection>
<intersection>-1226.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>134,-1234,134.5,-1234</points>
<connection>
<GID>2120</GID>
<name>IN_1</name></connection>
<intersection>134 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294.5,-1234.5,295,-1234.5</points>
<connection>
<GID>2126</GID>
<name>IN_1</name></connection>
<intersection>295 66</intersection></hsegment></shape></wire>
<wire>
<ID>1188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-1232,84,-1225.5</points>
<connection>
<GID>2118</GID>
<name>IN_0</name></connection>
<intersection>-1225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82.5,-1225.5,84,-1225.5</points>
<connection>
<GID>2117</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>1189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-1232,133.5,-1225.5</points>
<intersection>-1232 1</intersection>
<intersection>-1225.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-1232,134.5,-1232</points>
<connection>
<GID>2120</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,-1225.5,133.5,-1225.5</points>
<connection>
<GID>2119</GID>
<name>OUT_0</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-1231.5,182,-1225.5</points>
<intersection>-1231.5 5</intersection>
<intersection>-1225.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>180,-1225.5,182,-1225.5</points>
<connection>
<GID>2121</GID>
<name>OUT_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182,-1231.5,182.5,-1231.5</points>
<connection>
<GID>2122</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>1191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-1233.5,240.5,-1225.5</points>
<intersection>-1233.5 1</intersection>
<intersection>-1225.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240.5,-1233.5,241,-1233.5</points>
<connection>
<GID>2124</GID>
<name>IN_0</name></connection>
<intersection>240.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237.5,-1225.5,240.5,-1225.5</points>
<connection>
<GID>2123</GID>
<name>OUT_0</name></connection>
<intersection>240.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-1232.5,294,-1225.5</points>
<intersection>-1232.5 4</intersection>
<intersection>-1225.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292.5,-1225.5,294,-1225.5</points>
<connection>
<GID>2125</GID>
<name>OUT_0</name></connection>
<intersection>294 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294,-1232.5,294.5,-1232.5</points>
<connection>
<GID>2126</GID>
<name>IN_0</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>1193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352.5,-1233,352.5,-1225.5</points>
<intersection>-1233 1</intersection>
<intersection>-1225.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352.5,-1233,353,-1233</points>
<connection>
<GID>2128</GID>
<name>IN_0</name></connection>
<intersection>352.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-1225.5,352.5,-1225.5</points>
<connection>
<GID>2127</GID>
<name>OUT_0</name></connection>
<intersection>352.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-1245,-14,-1238.5</points>
<intersection>-1245 1</intersection>
<intersection>-1238.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-1245,-11.5,-1245</points>
<connection>
<GID>2131</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-1238.5,-14,-1238.5</points>
<connection>
<GID>2130</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1246,35,-1238.5</points>
<intersection>-1246 1</intersection>
<intersection>-1238.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1246,37,-1246</points>
<connection>
<GID>2133</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-1238.5,35,-1238.5</points>
<connection>
<GID>2132</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-1239.5,352.5,-1239.5</points>
<connection>
<GID>2146</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-1247,-13,-1239.5</points>
<intersection>-1247 5</intersection>
<intersection>-1239.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-1247,-11.5,-1247</points>
<connection>
<GID>2131</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-1248,35.5,-1239.5</points>
<intersection>-1248 21</intersection>
<intersection>-1239.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-1248,37,-1248</points>
<connection>
<GID>2133</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-1247,83,-1239.5</points>
<intersection>-1247 53</intersection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-1247,133.5,-1239.5</points>
<intersection>-1247 115</intersection>
<intersection>-1239.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-1247,83.5,-1247</points>
<connection>
<GID>2135</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-1246.5,182,-1239.5</points>
<connection>
<GID>2139</GID>
<name>IN_1</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-1248.5,240.5,-1239.5</points>
<connection>
<GID>2141</GID>
<name>IN_1</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-1247.5,294.5,-1239.5</points>
<intersection>-1247.5 118</intersection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-1248,352.5,-1239.5</points>
<connection>
<GID>2145</GID>
<name>IN_1</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-1241.5,-21.5,-1239.5</points>
<connection>
<GID>2130</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-1241.5,28,-1239.5</points>
<connection>
<GID>2132</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-1241.5,76,-1239.5</points>
<connection>
<GID>2134</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-1241.5,125.5,-1239.5</points>
<connection>
<GID>2136</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-1241.5,173.5,-1239.5</points>
<connection>
<GID>2138</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-1241.5,231,-1239.5</points>
<connection>
<GID>2140</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-1241.5,286,-1239.5</points>
<connection>
<GID>2142</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-1241.5,343,-1239.5</points>
<connection>
<GID>2144</GID>
<name>clock</name></connection>
<intersection>-1239.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-1247,134,-1247</points>
<connection>
<GID>2137</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-1247.5,294.5,-1247.5</points>
<connection>
<GID>2143</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1245,83.5,-1238.5</points>
<connection>
<GID>2135</GID>
<name>IN_0</name></connection>
<intersection>-1238.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-1238.5,83.5,-1238.5</points>
<connection>
<GID>2134</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1245,133,-1238.5</points>
<intersection>-1245 1</intersection>
<intersection>-1238.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-1245,134,-1245</points>
<connection>
<GID>2137</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-1238.5,133,-1238.5</points>
<connection>
<GID>2136</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1244.5,181.5,-1238.5</points>
<intersection>-1244.5 5</intersection>
<intersection>-1238.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-1238.5,181.5,-1238.5</points>
<connection>
<GID>2138</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-1244.5,182,-1244.5</points>
<connection>
<GID>2139</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-1246.5,240,-1238.5</points>
<intersection>-1246.5 1</intersection>
<intersection>-1238.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-1246.5,240.5,-1246.5</points>
<connection>
<GID>2141</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-1238.5,240,-1238.5</points>
<connection>
<GID>2140</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1245.5,293.5,-1238.5</points>
<intersection>-1245.5 4</intersection>
<intersection>-1238.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-1238.5,293.5,-1238.5</points>
<connection>
<GID>2142</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-1245.5,294,-1245.5</points>
<connection>
<GID>2143</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-1246,352,-1238.5</points>
<intersection>-1246 1</intersection>
<intersection>-1238.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-1246,352.5,-1246</points>
<connection>
<GID>2145</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-1238.5,352,-1238.5</points>
<connection>
<GID>2144</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-1260,-14,-1253.5</points>
<intersection>-1260 1</intersection>
<intersection>-1253.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-1260,-11.5,-1260</points>
<connection>
<GID>2012</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-1253.5,-14,-1253.5</points>
<connection>
<GID>2011</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1261,35,-1253.5</points>
<intersection>-1261 1</intersection>
<intersection>-1253.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1261,37,-1261</points>
<connection>
<GID>2014</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-1253.5,35,-1253.5</points>
<connection>
<GID>2013</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-1254.5,352.5,-1254.5</points>
<connection>
<GID>2027</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-1262,-13,-1254.5</points>
<intersection>-1262 5</intersection>
<intersection>-1254.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-1262,-11.5,-1262</points>
<connection>
<GID>2012</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-1263,35.5,-1254.5</points>
<intersection>-1263 21</intersection>
<intersection>-1254.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-1263,37,-1263</points>
<connection>
<GID>2014</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-1262,83,-1254.5</points>
<intersection>-1262 53</intersection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-1262,133.5,-1254.5</points>
<intersection>-1262 115</intersection>
<intersection>-1254.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-1262,83.5,-1262</points>
<connection>
<GID>2016</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-1261.5,182,-1254.5</points>
<connection>
<GID>2020</GID>
<name>IN_1</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-1263.5,240.5,-1254.5</points>
<connection>
<GID>2022</GID>
<name>IN_1</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-1262.5,294.5,-1254.5</points>
<intersection>-1262.5 118</intersection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-1263,352.5,-1254.5</points>
<connection>
<GID>2026</GID>
<name>IN_1</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-1256.5,-21.5,-1254.5</points>
<connection>
<GID>2011</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-1256.5,28,-1254.5</points>
<connection>
<GID>2013</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-1256.5,76,-1254.5</points>
<connection>
<GID>2015</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-1256.5,125.5,-1254.5</points>
<connection>
<GID>2017</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-1256.5,173.5,-1254.5</points>
<connection>
<GID>2019</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-1256.5,231,-1254.5</points>
<connection>
<GID>2021</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-1256.5,286,-1254.5</points>
<connection>
<GID>2023</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-1256.5,343,-1254.5</points>
<connection>
<GID>2025</GID>
<name>clock</name></connection>
<intersection>-1254.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-1262,134,-1262</points>
<connection>
<GID>2018</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-1262.5,294.5,-1262.5</points>
<connection>
<GID>2024</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1260,83.5,-1253.5</points>
<connection>
<GID>2016</GID>
<name>IN_0</name></connection>
<intersection>-1253.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-1253.5,83.5,-1253.5</points>
<connection>
<GID>2015</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1260,133,-1253.5</points>
<intersection>-1260 1</intersection>
<intersection>-1253.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-1260,134,-1260</points>
<connection>
<GID>2018</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-1253.5,133,-1253.5</points>
<connection>
<GID>2017</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1259.5,181.5,-1253.5</points>
<intersection>-1259.5 5</intersection>
<intersection>-1253.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-1253.5,181.5,-1253.5</points>
<connection>
<GID>2019</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-1259.5,182,-1259.5</points>
<connection>
<GID>2020</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-1261.5,240,-1253.5</points>
<intersection>-1261.5 1</intersection>
<intersection>-1253.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-1261.5,240.5,-1261.5</points>
<connection>
<GID>2022</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-1253.5,240,-1253.5</points>
<connection>
<GID>2021</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1260.5,293.5,-1253.5</points>
<intersection>-1260.5 4</intersection>
<intersection>-1253.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-1253.5,293.5,-1253.5</points>
<connection>
<GID>2023</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-1260.5,294,-1260.5</points>
<connection>
<GID>2024</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-1261,352,-1253.5</points>
<intersection>-1261 1</intersection>
<intersection>-1253.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-1261,352.5,-1261</points>
<connection>
<GID>2026</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-1253.5,352,-1253.5</points>
<connection>
<GID>2025</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-1274,-14,-1267.5</points>
<intersection>-1274 1</intersection>
<intersection>-1267.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-1274,-11.5,-1274</points>
<connection>
<GID>2029</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-1267.5,-14,-1267.5</points>
<connection>
<GID>2028</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1275,35,-1267.5</points>
<intersection>-1275 1</intersection>
<intersection>-1267.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1275,37,-1275</points>
<connection>
<GID>2031</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-1267.5,35,-1267.5</points>
<connection>
<GID>2030</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-1268.5,352.5,-1268.5</points>
<connection>
<GID>2044</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-1276,-13,-1268.5</points>
<intersection>-1276 5</intersection>
<intersection>-1268.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-1276,-11.5,-1276</points>
<connection>
<GID>2029</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-1277,35.5,-1268.5</points>
<intersection>-1277 21</intersection>
<intersection>-1268.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-1277,37,-1277</points>
<connection>
<GID>2031</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-1276,83,-1268.5</points>
<intersection>-1276 53</intersection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-1276,133.5,-1268.5</points>
<intersection>-1276 115</intersection>
<intersection>-1268.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-1276,83.5,-1276</points>
<connection>
<GID>2033</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-1275.5,182,-1268.5</points>
<connection>
<GID>2037</GID>
<name>IN_1</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-1277.5,240.5,-1268.5</points>
<connection>
<GID>2039</GID>
<name>IN_1</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-1276.5,294.5,-1268.5</points>
<intersection>-1276.5 118</intersection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-1277,352.5,-1268.5</points>
<connection>
<GID>2043</GID>
<name>IN_1</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-1270.5,-21.5,-1268.5</points>
<connection>
<GID>2028</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-1270.5,28,-1268.5</points>
<connection>
<GID>2030</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-1270.5,76,-1268.5</points>
<connection>
<GID>2032</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-1270.5,125.5,-1268.5</points>
<connection>
<GID>2034</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-1270.5,173.5,-1268.5</points>
<connection>
<GID>2036</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-1270.5,231,-1268.5</points>
<connection>
<GID>2038</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-1270.5,286,-1268.5</points>
<connection>
<GID>2040</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-1270.5,343,-1268.5</points>
<connection>
<GID>2042</GID>
<name>clock</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-1276,134,-1276</points>
<connection>
<GID>2035</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-1276.5,294.5,-1276.5</points>
<connection>
<GID>2041</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1274,83.5,-1267.5</points>
<connection>
<GID>2033</GID>
<name>IN_0</name></connection>
<intersection>-1267.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-1267.5,83.5,-1267.5</points>
<connection>
<GID>2032</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1274,133,-1267.5</points>
<intersection>-1274 1</intersection>
<intersection>-1267.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-1274,134,-1274</points>
<connection>
<GID>2035</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-1267.5,133,-1267.5</points>
<connection>
<GID>2034</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1273.5,181.5,-1267.5</points>
<intersection>-1273.5 5</intersection>
<intersection>-1267.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-1267.5,181.5,-1267.5</points>
<connection>
<GID>2036</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-1273.5,182,-1273.5</points>
<connection>
<GID>2037</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-1275.5,240,-1267.5</points>
<intersection>-1275.5 1</intersection>
<intersection>-1267.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-1275.5,240.5,-1275.5</points>
<connection>
<GID>2039</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-1267.5,240,-1267.5</points>
<connection>
<GID>2038</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1274.5,293.5,-1267.5</points>
<intersection>-1274.5 4</intersection>
<intersection>-1267.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-1267.5,293.5,-1267.5</points>
<connection>
<GID>2040</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-1274.5,294,-1274.5</points>
<connection>
<GID>2041</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-1275,352,-1267.5</points>
<intersection>-1275 1</intersection>
<intersection>-1267.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-1275,352.5,-1275</points>
<connection>
<GID>2043</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-1267.5,352,-1267.5</points>
<connection>
<GID>2042</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-1291.5,-14.5,-1285</points>
<intersection>-1291.5 1</intersection>
<intersection>-1285 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-1291.5,-12,-1291.5</points>
<connection>
<GID>2046</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-1285,-14.5,-1285</points>
<connection>
<GID>2045</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-1292.5,34.5,-1285</points>
<intersection>-1292.5 1</intersection>
<intersection>-1285 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-1292.5,36.5,-1292.5</points>
<connection>
<GID>2048</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-1285,34.5,-1285</points>
<connection>
<GID>2047</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47.5,-1286,352,-1286</points>
<connection>
<GID>2061</GID>
<name>OUT</name></connection>
<intersection>-22 107</intersection>
<intersection>-13.5 4</intersection>
<intersection>27.5 108</intersection>
<intersection>35 16</intersection>
<intersection>75.5 109</intersection>
<intersection>82.5 23</intersection>
<intersection>125 110</intersection>
<intersection>133 31</intersection>
<intersection>173 111</intersection>
<intersection>181.5 55</intersection>
<intersection>230.5 112</intersection>
<intersection>240 56</intersection>
<intersection>285.5 113</intersection>
<intersection>294 66</intersection>
<intersection>342.5 114</intersection>
<intersection>352 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13.5,-1293.5,-13.5,-1286</points>
<intersection>-1293.5 5</intersection>
<intersection>-1286 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13.5,-1293.5,-12,-1293.5</points>
<connection>
<GID>2046</GID>
<name>IN_1</name></connection>
<intersection>-13.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35,-1294.5,35,-1286</points>
<intersection>-1294.5 21</intersection>
<intersection>-1286 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35,-1294.5,36.5,-1294.5</points>
<connection>
<GID>2048</GID>
<name>IN_1</name></connection>
<intersection>35 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>82.5,-1293.5,82.5,-1286</points>
<intersection>-1293.5 53</intersection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133,-1293.5,133,-1286</points>
<intersection>-1293.5 115</intersection>
<intersection>-1286 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>82.5,-1293.5,83,-1293.5</points>
<connection>
<GID>2050</GID>
<name>IN_1</name></connection>
<intersection>82.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>181.5,-1293,181.5,-1286</points>
<connection>
<GID>2054</GID>
<name>IN_1</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240,-1295,240,-1286</points>
<connection>
<GID>2056</GID>
<name>IN_1</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294,-1294,294,-1286</points>
<intersection>-1294 118</intersection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352,-1294.5,352,-1286</points>
<connection>
<GID>2060</GID>
<name>IN_1</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-22,-1288,-22,-1286</points>
<connection>
<GID>2045</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>27.5,-1288,27.5,-1286</points>
<connection>
<GID>2047</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>75.5,-1288,75.5,-1286</points>
<connection>
<GID>2049</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125,-1288,125,-1286</points>
<connection>
<GID>2051</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173,-1288,173,-1286</points>
<connection>
<GID>2053</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>230.5,-1288,230.5,-1286</points>
<connection>
<GID>2055</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>285.5,-1288,285.5,-1286</points>
<connection>
<GID>2057</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>342.5,-1288,342.5,-1286</points>
<connection>
<GID>2059</GID>
<name>clock</name></connection>
<intersection>-1286 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133,-1293.5,133.5,-1293.5</points>
<connection>
<GID>2052</GID>
<name>IN_1</name></connection>
<intersection>133 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>293.5,-1294,294,-1294</points>
<connection>
<GID>2058</GID>
<name>IN_1</name></connection>
<intersection>294 66</intersection></hsegment></shape></wire>
<wire>
<ID>1224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-1291.5,83,-1285</points>
<connection>
<GID>2050</GID>
<name>IN_0</name></connection>
<intersection>-1285 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-1285,83,-1285</points>
<connection>
<GID>2049</GID>
<name>OUT_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>1225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-1291.5,132.5,-1285</points>
<intersection>-1291.5 1</intersection>
<intersection>-1285 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-1291.5,133.5,-1291.5</points>
<connection>
<GID>2052</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-1285,132.5,-1285</points>
<connection>
<GID>2051</GID>
<name>OUT_0</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-1291,181,-1285</points>
<intersection>-1291 5</intersection>
<intersection>-1285 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179,-1285,181,-1285</points>
<connection>
<GID>2053</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181,-1291,181.5,-1291</points>
<connection>
<GID>2054</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>1227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-1293,239.5,-1285</points>
<intersection>-1293 1</intersection>
<intersection>-1285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-1293,240,-1293</points>
<connection>
<GID>2056</GID>
<name>IN_0</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-1285,239.5,-1285</points>
<connection>
<GID>2055</GID>
<name>OUT_0</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-1292,293,-1285</points>
<intersection>-1292 4</intersection>
<intersection>-1285 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-1285,293,-1285</points>
<connection>
<GID>2057</GID>
<name>OUT_0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-1292,293.5,-1292</points>
<connection>
<GID>2058</GID>
<name>IN_0</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>1229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,-1292.5,351.5,-1285</points>
<intersection>-1292.5 1</intersection>
<intersection>-1285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,-1292.5,352,-1292.5</points>
<connection>
<GID>2060</GID>
<name>IN_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,-1285,351.5,-1285</points>
<connection>
<GID>2059</GID>
<name>OUT_0</name></connection>
<intersection>351.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70,-1234.5,-70,-1185.5</points>
<intersection>-1234.5 2</intersection>
<intersection>-1185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70,-1185.5,-52,-1185.5</points>
<connection>
<GID>2078</GID>
<name>IN_0</name></connection>
<intersection>-70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1234.5,-70,-1234.5</points>
<connection>
<GID>606</GID>
<name>OUT_7</name></connection>
<intersection>-70 0</intersection></hsegment></shape></wire>
<wire>
<ID>1231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-1235.5,-69,-1198.5</points>
<intersection>-1235.5 2</intersection>
<intersection>-1198.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-1198.5,-52,-1198.5</points>
<connection>
<GID>2095</GID>
<name>IN_0</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1235.5,-69,-1235.5</points>
<connection>
<GID>606</GID>
<name>OUT_6</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>1232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,-1236.5,-68,-1213</points>
<intersection>-1236.5 2</intersection>
<intersection>-1213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-1213,-52,-1213</points>
<connection>
<GID>2112</GID>
<name>IN_0</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1236.5,-68,-1236.5</points>
<connection>
<GID>606</GID>
<name>OUT_5</name></connection>
<intersection>-68 0</intersection></hsegment></shape></wire>
<wire>
<ID>1233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-1237.5,-67,-1225.5</points>
<intersection>-1237.5 2</intersection>
<intersection>-1225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,-1225.5,-52.5,-1225.5</points>
<connection>
<GID>2129</GID>
<name>IN_0</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1237.5,-67,-1237.5</points>
<connection>
<GID>606</GID>
<name>OUT_4</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>1234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-86,-1238.5,-53,-1238.5</points>
<connection>
<GID>2146</GID>
<name>IN_0</name></connection>
<connection>
<GID>606</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-1253.5,-67.5,-1239.5</points>
<intersection>-1253.5 1</intersection>
<intersection>-1239.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-1253.5,-53,-1253.5</points>
<connection>
<GID>2027</GID>
<name>IN_0</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1239.5,-67.5,-1239.5</points>
<connection>
<GID>606</GID>
<name>OUT_2</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-1267.5,-68.5,-1240.5</points>
<intersection>-1267.5 1</intersection>
<intersection>-1240.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,-1267.5,-53,-1267.5</points>
<connection>
<GID>2044</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1240.5,-68.5,-1240.5</points>
<connection>
<GID>606</GID>
<name>OUT_1</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-1285,-69.5,-1241.5</points>
<intersection>-1285 1</intersection>
<intersection>-1241.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-1285,-53.5,-1285</points>
<connection>
<GID>2061</GID>
<name>IN_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-1241.5,-69.5,-1241.5</points>
<connection>
<GID>606</GID>
<name>OUT_0</name></connection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-1435,-14,-1428.5</points>
<intersection>-1435 1</intersection>
<intersection>-1428.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-1435,-11.5,-1435</points>
<connection>
<GID>2335</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-1428.5,-14,-1428.5</points>
<connection>
<GID>2334</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1436,35,-1428.5</points>
<intersection>-1436 1</intersection>
<intersection>-1428.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1436,37,-1436</points>
<connection>
<GID>2337</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-1428.5,35,-1428.5</points>
<connection>
<GID>2336</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-1429.5,352.5,-1429.5</points>
<connection>
<GID>2350</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-1437,-13,-1429.5</points>
<intersection>-1437 5</intersection>
<intersection>-1429.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-1437,-11.5,-1437</points>
<connection>
<GID>2335</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-1438,35.5,-1429.5</points>
<intersection>-1438 21</intersection>
<intersection>-1429.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-1438,37,-1438</points>
<connection>
<GID>2337</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-1437,83,-1429.5</points>
<intersection>-1437 53</intersection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-1437,133.5,-1429.5</points>
<intersection>-1437 115</intersection>
<intersection>-1429.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-1437,83.5,-1437</points>
<connection>
<GID>2339</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-1436.5,182,-1429.5</points>
<connection>
<GID>2343</GID>
<name>IN_1</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-1438.5,240.5,-1429.5</points>
<connection>
<GID>2345</GID>
<name>IN_1</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-1437.5,294.5,-1429.5</points>
<intersection>-1437.5 118</intersection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-1438,352.5,-1429.5</points>
<connection>
<GID>2349</GID>
<name>IN_1</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-1431.5,-21.5,-1429.5</points>
<connection>
<GID>2334</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-1431.5,28,-1429.5</points>
<connection>
<GID>2336</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-1431.5,76,-1429.5</points>
<connection>
<GID>2338</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-1431.5,125.5,-1429.5</points>
<connection>
<GID>2340</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-1431.5,173.5,-1429.5</points>
<connection>
<GID>2342</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-1431.5,231,-1429.5</points>
<connection>
<GID>2344</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-1431.5,286,-1429.5</points>
<connection>
<GID>2346</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-1431.5,343,-1429.5</points>
<connection>
<GID>2348</GID>
<name>clock</name></connection>
<intersection>-1429.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-1437,134,-1437</points>
<connection>
<GID>2341</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-1437.5,294.5,-1437.5</points>
<connection>
<GID>2347</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1435,83.5,-1428.5</points>
<connection>
<GID>2339</GID>
<name>IN_0</name></connection>
<intersection>-1428.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-1428.5,83.5,-1428.5</points>
<connection>
<GID>2338</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1435,133,-1428.5</points>
<intersection>-1435 1</intersection>
<intersection>-1428.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-1435,134,-1435</points>
<connection>
<GID>2341</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-1428.5,133,-1428.5</points>
<connection>
<GID>2340</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1434.5,181.5,-1428.5</points>
<intersection>-1434.5 5</intersection>
<intersection>-1428.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-1428.5,181.5,-1428.5</points>
<connection>
<GID>2342</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-1434.5,182,-1434.5</points>
<connection>
<GID>2343</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-1436.5,240,-1428.5</points>
<intersection>-1436.5 1</intersection>
<intersection>-1428.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-1436.5,240.5,-1436.5</points>
<connection>
<GID>2345</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-1428.5,240,-1428.5</points>
<connection>
<GID>2344</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1435.5,293.5,-1428.5</points>
<intersection>-1435.5 4</intersection>
<intersection>-1428.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-1428.5,293.5,-1428.5</points>
<connection>
<GID>2346</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-1435.5,294,-1435.5</points>
<connection>
<GID>2347</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-1436,352,-1428.5</points>
<intersection>-1436 1</intersection>
<intersection>-1428.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-1436,352.5,-1436</points>
<connection>
<GID>2349</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-1428.5,352,-1428.5</points>
<connection>
<GID>2348</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-1448,-14,-1441.5</points>
<intersection>-1448 1</intersection>
<intersection>-1441.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-1448,-11.5,-1448</points>
<connection>
<GID>2352</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-1441.5,-14,-1441.5</points>
<connection>
<GID>2351</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1449,35,-1441.5</points>
<intersection>-1449 1</intersection>
<intersection>-1441.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1449,37,-1449</points>
<connection>
<GID>2354</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-1441.5,35,-1441.5</points>
<connection>
<GID>2353</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-1442.5,352.5,-1442.5</points>
<connection>
<GID>2367</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-1450,-13,-1442.5</points>
<intersection>-1450 5</intersection>
<intersection>-1442.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-1450,-11.5,-1450</points>
<connection>
<GID>2352</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-1451,35.5,-1442.5</points>
<intersection>-1451 21</intersection>
<intersection>-1442.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-1451,37,-1451</points>
<connection>
<GID>2354</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-1450,83,-1442.5</points>
<intersection>-1450 53</intersection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-1450,133.5,-1442.5</points>
<intersection>-1450 115</intersection>
<intersection>-1442.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-1450,83.5,-1450</points>
<connection>
<GID>2356</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-1449.5,182,-1442.5</points>
<connection>
<GID>2360</GID>
<name>IN_1</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-1451.5,240.5,-1442.5</points>
<connection>
<GID>2362</GID>
<name>IN_1</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-1450.5,294.5,-1442.5</points>
<intersection>-1450.5 118</intersection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-1451,352.5,-1442.5</points>
<connection>
<GID>2366</GID>
<name>IN_1</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-1444.5,-21.5,-1442.5</points>
<connection>
<GID>2351</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-1444.5,28,-1442.5</points>
<connection>
<GID>2353</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-1444.5,76,-1442.5</points>
<connection>
<GID>2355</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-1444.5,125.5,-1442.5</points>
<connection>
<GID>2357</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-1444.5,173.5,-1442.5</points>
<connection>
<GID>2359</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-1444.5,231,-1442.5</points>
<connection>
<GID>2361</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-1444.5,286,-1442.5</points>
<connection>
<GID>2363</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-1444.5,343,-1442.5</points>
<connection>
<GID>2365</GID>
<name>clock</name></connection>
<intersection>-1442.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-1450,134,-1450</points>
<connection>
<GID>2358</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-1450.5,294.5,-1450.5</points>
<connection>
<GID>2364</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1448,83.5,-1441.5</points>
<connection>
<GID>2356</GID>
<name>IN_0</name></connection>
<intersection>-1441.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-1441.5,83.5,-1441.5</points>
<connection>
<GID>2355</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1448,133,-1441.5</points>
<intersection>-1448 1</intersection>
<intersection>-1441.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-1448,134,-1448</points>
<connection>
<GID>2358</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-1441.5,133,-1441.5</points>
<connection>
<GID>2357</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1447.5,181.5,-1441.5</points>
<intersection>-1447.5 5</intersection>
<intersection>-1441.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-1441.5,181.5,-1441.5</points>
<connection>
<GID>2359</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-1447.5,182,-1447.5</points>
<connection>
<GID>2360</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-1449.5,240,-1441.5</points>
<intersection>-1449.5 1</intersection>
<intersection>-1441.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-1449.5,240.5,-1449.5</points>
<connection>
<GID>2362</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-1441.5,240,-1441.5</points>
<connection>
<GID>2361</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1448.5,293.5,-1441.5</points>
<intersection>-1448.5 4</intersection>
<intersection>-1441.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-1441.5,293.5,-1441.5</points>
<connection>
<GID>2363</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-1448.5,294,-1448.5</points>
<connection>
<GID>2364</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-1449,352,-1441.5</points>
<intersection>-1449 1</intersection>
<intersection>-1441.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-1449,352.5,-1449</points>
<connection>
<GID>2366</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-1441.5,352,-1441.5</points>
<connection>
<GID>2365</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-1462.5,-14,-1456</points>
<intersection>-1462.5 1</intersection>
<intersection>-1456 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-1462.5,-11.5,-1462.5</points>
<connection>
<GID>2369</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-1456,-14,-1456</points>
<connection>
<GID>2368</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>1331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1463.5,35,-1456</points>
<intersection>-1463.5 1</intersection>
<intersection>-1456 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1463.5,37,-1463.5</points>
<connection>
<GID>2371</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-1456,35,-1456</points>
<connection>
<GID>2370</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-1457,352.5,-1457</points>
<connection>
<GID>2384</GID>
<name>OUT</name></connection>
<intersection>-21.5 107</intersection>
<intersection>-13 4</intersection>
<intersection>28 108</intersection>
<intersection>35.5 16</intersection>
<intersection>76 109</intersection>
<intersection>83 23</intersection>
<intersection>125.5 110</intersection>
<intersection>133.5 31</intersection>
<intersection>173.5 111</intersection>
<intersection>182 55</intersection>
<intersection>231 112</intersection>
<intersection>240.5 56</intersection>
<intersection>286 113</intersection>
<intersection>294.5 66</intersection>
<intersection>343 114</intersection>
<intersection>352.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-1464.5,-13,-1457</points>
<intersection>-1464.5 5</intersection>
<intersection>-1457 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13,-1464.5,-11.5,-1464.5</points>
<connection>
<GID>2369</GID>
<name>IN_1</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35.5,-1465.5,35.5,-1457</points>
<intersection>-1465.5 21</intersection>
<intersection>-1457 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35.5,-1465.5,37,-1465.5</points>
<connection>
<GID>2371</GID>
<name>IN_1</name></connection>
<intersection>35.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>83,-1464.5,83,-1457</points>
<intersection>-1464.5 53</intersection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133.5,-1464.5,133.5,-1457</points>
<intersection>-1464.5 115</intersection>
<intersection>-1457 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>83,-1464.5,83.5,-1464.5</points>
<connection>
<GID>2373</GID>
<name>IN_1</name></connection>
<intersection>83 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>182,-1464,182,-1457</points>
<connection>
<GID>2377</GID>
<name>IN_1</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240.5,-1466,240.5,-1457</points>
<connection>
<GID>2379</GID>
<name>IN_1</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294.5,-1465,294.5,-1457</points>
<intersection>-1465 118</intersection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352.5,-1465.5,352.5,-1457</points>
<connection>
<GID>2383</GID>
<name>IN_1</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-21.5,-1459,-21.5,-1457</points>
<connection>
<GID>2368</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>28,-1459,28,-1457</points>
<connection>
<GID>2370</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>76,-1459,76,-1457</points>
<connection>
<GID>2372</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125.5,-1459,125.5,-1457</points>
<connection>
<GID>2374</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173.5,-1459,173.5,-1457</points>
<connection>
<GID>2376</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>231,-1459,231,-1457</points>
<connection>
<GID>2378</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>286,-1459,286,-1457</points>
<connection>
<GID>2380</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>343,-1459,343,-1457</points>
<connection>
<GID>2382</GID>
<name>clock</name></connection>
<intersection>-1457 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133.5,-1464.5,134,-1464.5</points>
<connection>
<GID>2375</GID>
<name>IN_1</name></connection>
<intersection>133.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>294,-1465,294.5,-1465</points>
<connection>
<GID>2381</GID>
<name>IN_1</name></connection>
<intersection>294.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1462.5,83.5,-1456</points>
<connection>
<GID>2373</GID>
<name>IN_0</name></connection>
<intersection>-1456 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82,-1456,83.5,-1456</points>
<connection>
<GID>2372</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-1462.5,133,-1456</points>
<intersection>-1462.5 1</intersection>
<intersection>-1456 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-1462.5,134,-1462.5</points>
<connection>
<GID>2375</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131.5,-1456,133,-1456</points>
<connection>
<GID>2374</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-1462,181.5,-1456</points>
<intersection>-1462 5</intersection>
<intersection>-1456 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179.5,-1456,181.5,-1456</points>
<connection>
<GID>2376</GID>
<name>OUT_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,-1462,182,-1462</points>
<connection>
<GID>2377</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-1464,240,-1456</points>
<intersection>-1464 1</intersection>
<intersection>-1456 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-1464,240.5,-1464</points>
<connection>
<GID>2379</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-1456,240,-1456</points>
<connection>
<GID>2378</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>1337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1463,293.5,-1456</points>
<intersection>-1463 4</intersection>
<intersection>-1456 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>292,-1456,293.5,-1456</points>
<connection>
<GID>2380</GID>
<name>OUT_0</name></connection>
<intersection>293.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-1463,294,-1463</points>
<connection>
<GID>2381</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-1463.5,352,-1456</points>
<intersection>-1463.5 1</intersection>
<intersection>-1456 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-1463.5,352.5,-1463.5</points>
<connection>
<GID>2383</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-1456,352,-1456</points>
<connection>
<GID>2382</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>1339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-1475,-14.5,-1468.5</points>
<intersection>-1475 1</intersection>
<intersection>-1468.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-1475,-12,-1475</points>
<connection>
<GID>2386</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-1468.5,-14.5,-1468.5</points>
<connection>
<GID>2385</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-1476,34.5,-1468.5</points>
<intersection>-1476 1</intersection>
<intersection>-1468.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-1476,36.5,-1476</points>
<connection>
<GID>2388</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-1468.5,34.5,-1468.5</points>
<connection>
<GID>2387</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47.5,-1469.5,352,-1469.5</points>
<connection>
<GID>2401</GID>
<name>OUT</name></connection>
<intersection>-22 107</intersection>
<intersection>-13.5 4</intersection>
<intersection>27.5 108</intersection>
<intersection>35 16</intersection>
<intersection>75.5 109</intersection>
<intersection>82.5 23</intersection>
<intersection>125 110</intersection>
<intersection>133 31</intersection>
<intersection>173 111</intersection>
<intersection>181.5 55</intersection>
<intersection>230.5 112</intersection>
<intersection>240 56</intersection>
<intersection>285.5 113</intersection>
<intersection>294 66</intersection>
<intersection>342.5 114</intersection>
<intersection>352 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13.5,-1477,-13.5,-1469.5</points>
<intersection>-1477 5</intersection>
<intersection>-1469.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13.5,-1477,-12,-1477</points>
<connection>
<GID>2386</GID>
<name>IN_1</name></connection>
<intersection>-13.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>35,-1478,35,-1469.5</points>
<intersection>-1478 21</intersection>
<intersection>-1469.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>35,-1478,36.5,-1478</points>
<connection>
<GID>2388</GID>
<name>IN_1</name></connection>
<intersection>35 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>82.5,-1477,82.5,-1469.5</points>
<intersection>-1477 53</intersection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>133,-1477,133,-1469.5</points>
<intersection>-1477 115</intersection>
<intersection>-1469.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>82.5,-1477,83,-1477</points>
<connection>
<GID>2390</GID>
<name>IN_1</name></connection>
<intersection>82.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>181.5,-1476.5,181.5,-1469.5</points>
<connection>
<GID>2394</GID>
<name>IN_1</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>240,-1478.5,240,-1469.5</points>
<connection>
<GID>2396</GID>
<name>IN_1</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>294,-1477.5,294,-1469.5</points>
<intersection>-1477.5 118</intersection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>352,-1478,352,-1469.5</points>
<connection>
<GID>2400</GID>
<name>IN_1</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-22,-1471.5,-22,-1469.5</points>
<connection>
<GID>2385</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>27.5,-1471.5,27.5,-1469.5</points>
<connection>
<GID>2387</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>75.5,-1471.5,75.5,-1469.5</points>
<connection>
<GID>2389</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>125,-1471.5,125,-1469.5</points>
<connection>
<GID>2391</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>173,-1471.5,173,-1469.5</points>
<connection>
<GID>2393</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>230.5,-1471.5,230.5,-1469.5</points>
<connection>
<GID>2395</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>285.5,-1471.5,285.5,-1469.5</points>
<connection>
<GID>2397</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>342.5,-1471.5,342.5,-1469.5</points>
<connection>
<GID>2399</GID>
<name>clock</name></connection>
<intersection>-1469.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>133,-1477,133.5,-1477</points>
<connection>
<GID>2392</GID>
<name>IN_1</name></connection>
<intersection>133 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>293.5,-1477.5,294,-1477.5</points>
<connection>
<GID>2398</GID>
<name>IN_1</name></connection>
<intersection>294 66</intersection></hsegment></shape></wire>
<wire>
<ID>1342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-1475,83,-1468.5</points>
<connection>
<GID>2390</GID>
<name>IN_0</name></connection>
<intersection>-1468.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-1468.5,83,-1468.5</points>
<connection>
<GID>2389</GID>
<name>OUT_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>1343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-1475,132.5,-1468.5</points>
<intersection>-1475 1</intersection>
<intersection>-1468.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-1475,133.5,-1475</points>
<connection>
<GID>2392</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-1468.5,132.5,-1468.5</points>
<connection>
<GID>2391</GID>
<name>OUT_0</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-1474.5,181,-1468.5</points>
<intersection>-1474.5 5</intersection>
<intersection>-1468.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>179,-1468.5,181,-1468.5</points>
<connection>
<GID>2393</GID>
<name>OUT_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181,-1474.5,181.5,-1474.5</points>
<connection>
<GID>2394</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>1345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239.5,-1476.5,239.5,-1468.5</points>
<intersection>-1476.5 1</intersection>
<intersection>-1468.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239.5,-1476.5,240,-1476.5</points>
<connection>
<GID>2396</GID>
<name>IN_0</name></connection>
<intersection>239.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236.5,-1468.5,239.5,-1468.5</points>
<connection>
<GID>2395</GID>
<name>OUT_0</name></connection>
<intersection>239.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-1475.5,293,-1468.5</points>
<intersection>-1475.5 4</intersection>
<intersection>-1468.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-1468.5,293,-1468.5</points>
<connection>
<GID>2397</GID>
<name>OUT_0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>293,-1475.5,293.5,-1475.5</points>
<connection>
<GID>2398</GID>
<name>IN_0</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>1347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,-1476,351.5,-1468.5</points>
<intersection>-1476 1</intersection>
<intersection>-1468.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,-1476,352,-1476</points>
<connection>
<GID>2400</GID>
<name>IN_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,-1468.5,351.5,-1468.5</points>
<connection>
<GID>2399</GID>
<name>OUT_0</name></connection>
<intersection>351.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-1488,-15,-1481.5</points>
<intersection>-1488 1</intersection>
<intersection>-1481.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-1488,-12.5,-1488</points>
<connection>
<GID>2403</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16.5,-1481.5,-15,-1481.5</points>
<connection>
<GID>2402</GID>
<name>OUT_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>1349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-1489,34,-1481.5</points>
<intersection>-1489 1</intersection>
<intersection>-1481.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-1489,36,-1489</points>
<connection>
<GID>2405</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-1481.5,34,-1481.5</points>
<connection>
<GID>2404</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>1350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-1482.5,351.5,-1482.5</points>
<connection>
<GID>2418</GID>
<name>OUT</name></connection>
<intersection>-22.5 107</intersection>
<intersection>-14 4</intersection>
<intersection>27 108</intersection>
<intersection>34.5 16</intersection>
<intersection>75 109</intersection>
<intersection>82 23</intersection>
<intersection>124.5 110</intersection>
<intersection>132.5 31</intersection>
<intersection>172.5 111</intersection>
<intersection>181 55</intersection>
<intersection>230 112</intersection>
<intersection>239.5 56</intersection>
<intersection>285 113</intersection>
<intersection>293.5 66</intersection>
<intersection>342 114</intersection>
<intersection>351.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-14,-1490,-14,-1482.5</points>
<intersection>-1490 5</intersection>
<intersection>-1482.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-14,-1490,-12.5,-1490</points>
<connection>
<GID>2403</GID>
<name>IN_1</name></connection>
<intersection>-14 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>34.5,-1491,34.5,-1482.5</points>
<intersection>-1491 21</intersection>
<intersection>-1482.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>34.5,-1491,36,-1491</points>
<connection>
<GID>2405</GID>
<name>IN_1</name></connection>
<intersection>34.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>82,-1490,82,-1482.5</points>
<intersection>-1490 53</intersection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>132.5,-1490,132.5,-1482.5</points>
<intersection>-1490 115</intersection>
<intersection>-1482.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>82,-1490,82.5,-1490</points>
<connection>
<GID>2407</GID>
<name>IN_1</name></connection>
<intersection>82 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>181,-1489.5,181,-1482.5</points>
<connection>
<GID>2411</GID>
<name>IN_1</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>239.5,-1491.5,239.5,-1482.5</points>
<connection>
<GID>2413</GID>
<name>IN_1</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>293.5,-1490.5,293.5,-1482.5</points>
<intersection>-1490.5 118</intersection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>351.5,-1491,351.5,-1482.5</points>
<connection>
<GID>2417</GID>
<name>IN_1</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-22.5,-1484.5,-22.5,-1482.5</points>
<connection>
<GID>2402</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>27,-1484.5,27,-1482.5</points>
<connection>
<GID>2404</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>75,-1484.5,75,-1482.5</points>
<connection>
<GID>2406</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>124.5,-1484.5,124.5,-1482.5</points>
<connection>
<GID>2408</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>172.5,-1484.5,172.5,-1482.5</points>
<connection>
<GID>2410</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>230,-1484.5,230,-1482.5</points>
<connection>
<GID>2412</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>285,-1484.5,285,-1482.5</points>
<connection>
<GID>2414</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>342,-1484.5,342,-1482.5</points>
<connection>
<GID>2416</GID>
<name>clock</name></connection>
<intersection>-1482.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>132.5,-1490,133,-1490</points>
<connection>
<GID>2409</GID>
<name>IN_1</name></connection>
<intersection>132.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>293,-1490.5,293.5,-1490.5</points>
<connection>
<GID>2415</GID>
<name>IN_1</name></connection>
<intersection>293.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-1488,82.5,-1481.5</points>
<connection>
<GID>2407</GID>
<name>IN_0</name></connection>
<intersection>-1481.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81,-1481.5,82.5,-1481.5</points>
<connection>
<GID>2406</GID>
<name>OUT_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-1488,132,-1481.5</points>
<intersection>-1488 1</intersection>
<intersection>-1481.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-1488,133,-1488</points>
<connection>
<GID>2409</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130.5,-1481.5,132,-1481.5</points>
<connection>
<GID>2408</GID>
<name>OUT_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>1353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-1487.5,180.5,-1481.5</points>
<intersection>-1487.5 5</intersection>
<intersection>-1481.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>178.5,-1481.5,180.5,-1481.5</points>
<connection>
<GID>2410</GID>
<name>OUT_0</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>180.5,-1487.5,181,-1487.5</points>
<connection>
<GID>2411</GID>
<name>IN_0</name></connection>
<intersection>180.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-1489.5,239,-1481.5</points>
<intersection>-1489.5 1</intersection>
<intersection>-1481.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-1489.5,239.5,-1489.5</points>
<connection>
<GID>2413</GID>
<name>IN_0</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236,-1481.5,239,-1481.5</points>
<connection>
<GID>2412</GID>
<name>OUT_0</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>1355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-1488.5,292.5,-1481.5</points>
<intersection>-1488.5 4</intersection>
<intersection>-1481.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291,-1481.5,292.5,-1481.5</points>
<connection>
<GID>2414</GID>
<name>OUT_0</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-1488.5,293,-1488.5</points>
<connection>
<GID>2415</GID>
<name>IN_0</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-1489,351,-1481.5</points>
<intersection>-1489 1</intersection>
<intersection>-1481.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,-1489,351.5,-1489</points>
<connection>
<GID>2417</GID>
<name>IN_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348,-1481.5,351,-1481.5</points>
<connection>
<GID>2416</GID>
<name>OUT_0</name></connection>
<intersection>351 0</intersection></hsegment></shape></wire>
<wire>
<ID>1357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-1503,-15,-1496.5</points>
<intersection>-1503 1</intersection>
<intersection>-1496.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-1503,-12.5,-1503</points>
<connection>
<GID>2284</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16.5,-1496.5,-15,-1496.5</points>
<connection>
<GID>2283</GID>
<name>OUT_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>1358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-1504,34,-1496.5</points>
<intersection>-1504 1</intersection>
<intersection>-1496.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-1504,36,-1504</points>
<connection>
<GID>2286</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-1496.5,34,-1496.5</points>
<connection>
<GID>2285</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>1359</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-1497.5,351.5,-1497.5</points>
<connection>
<GID>2299</GID>
<name>OUT</name></connection>
<intersection>-22.5 107</intersection>
<intersection>-14 4</intersection>
<intersection>27 108</intersection>
<intersection>34.5 16</intersection>
<intersection>75 109</intersection>
<intersection>82 23</intersection>
<intersection>124.5 110</intersection>
<intersection>132.5 31</intersection>
<intersection>172.5 111</intersection>
<intersection>181 55</intersection>
<intersection>230 112</intersection>
<intersection>239.5 56</intersection>
<intersection>285 113</intersection>
<intersection>293.5 66</intersection>
<intersection>342 114</intersection>
<intersection>351.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-14,-1505,-14,-1497.5</points>
<intersection>-1505 5</intersection>
<intersection>-1497.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-14,-1505,-12.5,-1505</points>
<connection>
<GID>2284</GID>
<name>IN_1</name></connection>
<intersection>-14 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>34.5,-1506,34.5,-1497.5</points>
<intersection>-1506 21</intersection>
<intersection>-1497.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>34.5,-1506,36,-1506</points>
<connection>
<GID>2286</GID>
<name>IN_1</name></connection>
<intersection>34.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>82,-1505,82,-1497.5</points>
<intersection>-1505 53</intersection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>132.5,-1505,132.5,-1497.5</points>
<intersection>-1505 115</intersection>
<intersection>-1497.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>82,-1505,82.5,-1505</points>
<connection>
<GID>2288</GID>
<name>IN_1</name></connection>
<intersection>82 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>181,-1504.5,181,-1497.5</points>
<connection>
<GID>2292</GID>
<name>IN_1</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>239.5,-1506.5,239.5,-1497.5</points>
<connection>
<GID>2294</GID>
<name>IN_1</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>293.5,-1505.5,293.5,-1497.5</points>
<intersection>-1505.5 118</intersection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>351.5,-1506,351.5,-1497.5</points>
<connection>
<GID>2298</GID>
<name>IN_1</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-22.5,-1499.5,-22.5,-1497.5</points>
<connection>
<GID>2283</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>27,-1499.5,27,-1497.5</points>
<connection>
<GID>2285</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>75,-1499.5,75,-1497.5</points>
<connection>
<GID>2287</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>124.5,-1499.5,124.5,-1497.5</points>
<connection>
<GID>2289</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>172.5,-1499.5,172.5,-1497.5</points>
<connection>
<GID>2291</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>230,-1499.5,230,-1497.5</points>
<connection>
<GID>2293</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>285,-1499.5,285,-1497.5</points>
<connection>
<GID>2295</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>342,-1499.5,342,-1497.5</points>
<connection>
<GID>2297</GID>
<name>clock</name></connection>
<intersection>-1497.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>132.5,-1505,133,-1505</points>
<connection>
<GID>2290</GID>
<name>IN_1</name></connection>
<intersection>132.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>293,-1505.5,293.5,-1505.5</points>
<connection>
<GID>2296</GID>
<name>IN_1</name></connection>
<intersection>293.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-1503,82.5,-1496.5</points>
<connection>
<GID>2288</GID>
<name>IN_0</name></connection>
<intersection>-1496.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81,-1496.5,82.5,-1496.5</points>
<connection>
<GID>2287</GID>
<name>OUT_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-1503,132,-1496.5</points>
<intersection>-1503 1</intersection>
<intersection>-1496.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-1503,133,-1503</points>
<connection>
<GID>2290</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130.5,-1496.5,132,-1496.5</points>
<connection>
<GID>2289</GID>
<name>OUT_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>1362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-1502.5,180.5,-1496.5</points>
<intersection>-1502.5 5</intersection>
<intersection>-1496.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>178.5,-1496.5,180.5,-1496.5</points>
<connection>
<GID>2291</GID>
<name>OUT_0</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>180.5,-1502.5,181,-1502.5</points>
<connection>
<GID>2292</GID>
<name>IN_0</name></connection>
<intersection>180.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-1504.5,239,-1496.5</points>
<intersection>-1504.5 1</intersection>
<intersection>-1496.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-1504.5,239.5,-1504.5</points>
<connection>
<GID>2294</GID>
<name>IN_0</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236,-1496.5,239,-1496.5</points>
<connection>
<GID>2293</GID>
<name>OUT_0</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>1364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-1503.5,292.5,-1496.5</points>
<intersection>-1503.5 4</intersection>
<intersection>-1496.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291,-1496.5,292.5,-1496.5</points>
<connection>
<GID>2295</GID>
<name>OUT_0</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-1503.5,293,-1503.5</points>
<connection>
<GID>2296</GID>
<name>IN_0</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-1504,351,-1496.5</points>
<intersection>-1504 1</intersection>
<intersection>-1496.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,-1504,351.5,-1504</points>
<connection>
<GID>2298</GID>
<name>IN_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348,-1496.5,351,-1496.5</points>
<connection>
<GID>2297</GID>
<name>OUT_0</name></connection>
<intersection>351 0</intersection></hsegment></shape></wire>
<wire>
<ID>1366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-1517,-15,-1510.5</points>
<intersection>-1517 1</intersection>
<intersection>-1510.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-1517,-12.5,-1517</points>
<connection>
<GID>2301</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16.5,-1510.5,-15,-1510.5</points>
<connection>
<GID>2300</GID>
<name>OUT_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>1367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-1518,34,-1510.5</points>
<intersection>-1518 1</intersection>
<intersection>-1510.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-1518,36,-1518</points>
<connection>
<GID>2303</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-1510.5,34,-1510.5</points>
<connection>
<GID>2302</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>1368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-1511.5,351.5,-1511.5</points>
<connection>
<GID>2316</GID>
<name>OUT</name></connection>
<intersection>-22.5 107</intersection>
<intersection>-14 4</intersection>
<intersection>27 108</intersection>
<intersection>34.5 16</intersection>
<intersection>75 109</intersection>
<intersection>82 23</intersection>
<intersection>124.5 110</intersection>
<intersection>132.5 31</intersection>
<intersection>172.5 111</intersection>
<intersection>181 55</intersection>
<intersection>230 112</intersection>
<intersection>239.5 56</intersection>
<intersection>285 113</intersection>
<intersection>293.5 66</intersection>
<intersection>342 114</intersection>
<intersection>351.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-14,-1519,-14,-1511.5</points>
<intersection>-1519 5</intersection>
<intersection>-1511.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-14,-1519,-12.5,-1519</points>
<connection>
<GID>2301</GID>
<name>IN_1</name></connection>
<intersection>-14 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>34.5,-1520,34.5,-1511.5</points>
<intersection>-1520 21</intersection>
<intersection>-1511.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>34.5,-1520,36,-1520</points>
<connection>
<GID>2303</GID>
<name>IN_1</name></connection>
<intersection>34.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>82,-1519,82,-1511.5</points>
<intersection>-1519 53</intersection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>132.5,-1519,132.5,-1511.5</points>
<intersection>-1519 115</intersection>
<intersection>-1511.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>82,-1519,82.5,-1519</points>
<connection>
<GID>2305</GID>
<name>IN_1</name></connection>
<intersection>82 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>181,-1518.5,181,-1511.5</points>
<connection>
<GID>2309</GID>
<name>IN_1</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>239.5,-1520.5,239.5,-1511.5</points>
<connection>
<GID>2311</GID>
<name>IN_1</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>293.5,-1519.5,293.5,-1511.5</points>
<intersection>-1519.5 118</intersection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>351.5,-1520,351.5,-1511.5</points>
<connection>
<GID>2315</GID>
<name>IN_1</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-22.5,-1513.5,-22.5,-1511.5</points>
<connection>
<GID>2300</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>27,-1513.5,27,-1511.5</points>
<connection>
<GID>2302</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>75,-1513.5,75,-1511.5</points>
<connection>
<GID>2304</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>124.5,-1513.5,124.5,-1511.5</points>
<connection>
<GID>2306</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>172.5,-1513.5,172.5,-1511.5</points>
<connection>
<GID>2308</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>230,-1513.5,230,-1511.5</points>
<connection>
<GID>2310</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>285,-1513.5,285,-1511.5</points>
<connection>
<GID>2312</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>342,-1513.5,342,-1511.5</points>
<connection>
<GID>2314</GID>
<name>clock</name></connection>
<intersection>-1511.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>132.5,-1519,133,-1519</points>
<connection>
<GID>2307</GID>
<name>IN_1</name></connection>
<intersection>132.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>293,-1519.5,293.5,-1519.5</points>
<connection>
<GID>2313</GID>
<name>IN_1</name></connection>
<intersection>293.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-1517,82.5,-1510.5</points>
<connection>
<GID>2305</GID>
<name>IN_0</name></connection>
<intersection>-1510.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81,-1510.5,82.5,-1510.5</points>
<connection>
<GID>2304</GID>
<name>OUT_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-1517,132,-1510.5</points>
<intersection>-1517 1</intersection>
<intersection>-1510.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-1517,133,-1517</points>
<connection>
<GID>2307</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130.5,-1510.5,132,-1510.5</points>
<connection>
<GID>2306</GID>
<name>OUT_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>1371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-1516.5,180.5,-1510.5</points>
<intersection>-1516.5 5</intersection>
<intersection>-1510.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>178.5,-1510.5,180.5,-1510.5</points>
<connection>
<GID>2308</GID>
<name>OUT_0</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>180.5,-1516.5,181,-1516.5</points>
<connection>
<GID>2309</GID>
<name>IN_0</name></connection>
<intersection>180.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,-1518.5,239,-1510.5</points>
<intersection>-1518.5 1</intersection>
<intersection>-1510.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,-1518.5,239.5,-1518.5</points>
<connection>
<GID>2311</GID>
<name>IN_0</name></connection>
<intersection>239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236,-1510.5,239,-1510.5</points>
<connection>
<GID>2310</GID>
<name>OUT_0</name></connection>
<intersection>239 0</intersection></hsegment></shape></wire>
<wire>
<ID>1373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-1517.5,292.5,-1510.5</points>
<intersection>-1517.5 4</intersection>
<intersection>-1510.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291,-1510.5,292.5,-1510.5</points>
<connection>
<GID>2312</GID>
<name>OUT_0</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-1517.5,293,-1517.5</points>
<connection>
<GID>2313</GID>
<name>IN_0</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-1518,351,-1510.5</points>
<intersection>-1518 1</intersection>
<intersection>-1510.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,-1518,351.5,-1518</points>
<connection>
<GID>2315</GID>
<name>IN_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348,-1510.5,351,-1510.5</points>
<connection>
<GID>2314</GID>
<name>OUT_0</name></connection>
<intersection>351 0</intersection></hsegment></shape></wire>
<wire>
<ID>1375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-1534.5,-15.5,-1528</points>
<intersection>-1534.5 1</intersection>
<intersection>-1528 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-1534.5,-13,-1534.5</points>
<connection>
<GID>2318</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17,-1528,-15.5,-1528</points>
<connection>
<GID>2317</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-1535.5,33.5,-1528</points>
<intersection>-1535.5 1</intersection>
<intersection>-1528 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-1535.5,35.5,-1535.5</points>
<connection>
<GID>2320</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-1528,33.5,-1528</points>
<connection>
<GID>2319</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48.5,-1529,351,-1529</points>
<connection>
<GID>2333</GID>
<name>OUT</name></connection>
<intersection>-23 107</intersection>
<intersection>-14.5 4</intersection>
<intersection>26.5 108</intersection>
<intersection>34 16</intersection>
<intersection>74.5 109</intersection>
<intersection>81.5 23</intersection>
<intersection>124 110</intersection>
<intersection>132 31</intersection>
<intersection>172 111</intersection>
<intersection>180.5 55</intersection>
<intersection>229.5 112</intersection>
<intersection>239 56</intersection>
<intersection>284.5 113</intersection>
<intersection>293 66</intersection>
<intersection>341.5 114</intersection>
<intersection>351 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-14.5,-1536.5,-14.5,-1529</points>
<intersection>-1536.5 5</intersection>
<intersection>-1529 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-14.5,-1536.5,-13,-1536.5</points>
<connection>
<GID>2318</GID>
<name>IN_1</name></connection>
<intersection>-14.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>34,-1537.5,34,-1529</points>
<intersection>-1537.5 21</intersection>
<intersection>-1529 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>34,-1537.5,35.5,-1537.5</points>
<connection>
<GID>2320</GID>
<name>IN_1</name></connection>
<intersection>34 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>81.5,-1536.5,81.5,-1529</points>
<intersection>-1536.5 53</intersection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>132,-1536.5,132,-1529</points>
<intersection>-1536.5 115</intersection>
<intersection>-1529 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>81.5,-1536.5,82,-1536.5</points>
<connection>
<GID>2322</GID>
<name>IN_1</name></connection>
<intersection>81.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>180.5,-1536,180.5,-1529</points>
<connection>
<GID>2326</GID>
<name>IN_1</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>239,-1538,239,-1529</points>
<connection>
<GID>2328</GID>
<name>IN_1</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>293,-1537,293,-1529</points>
<intersection>-1537 118</intersection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>351,-1537.5,351,-1529</points>
<connection>
<GID>2332</GID>
<name>IN_1</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-23,-1531,-23,-1529</points>
<connection>
<GID>2317</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>26.5,-1531,26.5,-1529</points>
<connection>
<GID>2319</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>74.5,-1531,74.5,-1529</points>
<connection>
<GID>2321</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>124,-1531,124,-1529</points>
<connection>
<GID>2323</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>172,-1531,172,-1529</points>
<connection>
<GID>2325</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>229.5,-1531,229.5,-1529</points>
<connection>
<GID>2327</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>284.5,-1531,284.5,-1529</points>
<connection>
<GID>2329</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>341.5,-1531,341.5,-1529</points>
<connection>
<GID>2331</GID>
<name>clock</name></connection>
<intersection>-1529 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>132,-1536.5,132.5,-1536.5</points>
<connection>
<GID>2324</GID>
<name>IN_1</name></connection>
<intersection>132 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>292.5,-1537,293,-1537</points>
<connection>
<GID>2330</GID>
<name>IN_1</name></connection>
<intersection>293 66</intersection></hsegment></shape></wire>
<wire>
<ID>1378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-1534.5,82,-1528</points>
<connection>
<GID>2322</GID>
<name>IN_0</name></connection>
<intersection>-1528 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>80.5,-1528,82,-1528</points>
<connection>
<GID>2321</GID>
<name>OUT_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>1379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-1534.5,131.5,-1528</points>
<intersection>-1534.5 1</intersection>
<intersection>-1528 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-1534.5,132.5,-1534.5</points>
<connection>
<GID>2324</GID>
<name>IN_0</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130,-1528,131.5,-1528</points>
<connection>
<GID>2323</GID>
<name>OUT_0</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-1534,180,-1528</points>
<intersection>-1534 5</intersection>
<intersection>-1528 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>178,-1528,180,-1528</points>
<connection>
<GID>2325</GID>
<name>OUT_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>180,-1534,180.5,-1534</points>
<connection>
<GID>2326</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>1381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-1536,238.5,-1528</points>
<intersection>-1536 1</intersection>
<intersection>-1528 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,-1536,239,-1536</points>
<connection>
<GID>2328</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235.5,-1528,238.5,-1528</points>
<connection>
<GID>2327</GID>
<name>OUT_0</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-1535,292,-1528</points>
<intersection>-1535 4</intersection>
<intersection>-1528 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>290.5,-1528,292,-1528</points>
<connection>
<GID>2329</GID>
<name>OUT_0</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292,-1535,292.5,-1535</points>
<connection>
<GID>2330</GID>
<name>IN_0</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>1383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350.5,-1535.5,350.5,-1528</points>
<intersection>-1535.5 1</intersection>
<intersection>-1528 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350.5,-1535.5,351,-1535.5</points>
<connection>
<GID>2332</GID>
<name>IN_0</name></connection>
<intersection>350.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347.5,-1528,350.5,-1528</points>
<connection>
<GID>2331</GID>
<name>OUT_0</name></connection>
<intersection>350.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-1471,-67.5,-1428.5</points>
<intersection>-1471 2</intersection>
<intersection>-1428.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-1428.5,-53,-1428.5</points>
<connection>
<GID>2350</GID>
<name>IN_0</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1471,-67.5,-1471</points>
<connection>
<GID>743</GID>
<name>OUT_7</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-1472,-66.5,-1441.5</points>
<intersection>-1472 2</intersection>
<intersection>-1441.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,-1441.5,-53,-1441.5</points>
<connection>
<GID>2367</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1472,-66.5,-1472</points>
<connection>
<GID>743</GID>
<name>OUT_6</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,-1473,-65.5,-1456</points>
<intersection>-1473 2</intersection>
<intersection>-1456 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,-1456,-53,-1456</points>
<connection>
<GID>2384</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1473,-65.5,-1473</points>
<connection>
<GID>743</GID>
<name>OUT_5</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-1474,-64.5,-1468.5</points>
<intersection>-1474 2</intersection>
<intersection>-1468.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-1468.5,-53.5,-1468.5</points>
<connection>
<GID>2401</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1474,-64.5,-1474</points>
<connection>
<GID>743</GID>
<name>OUT_4</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-1481.5,-64.5,-1475</points>
<intersection>-1481.5 1</intersection>
<intersection>-1475 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-1481.5,-54,-1481.5</points>
<connection>
<GID>2418</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1475,-64.5,-1475</points>
<connection>
<GID>743</GID>
<name>OUT_3</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,-1496.5,-65.5,-1476</points>
<intersection>-1496.5 1</intersection>
<intersection>-1476 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,-1496.5,-54,-1496.5</points>
<connection>
<GID>2299</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1476,-65.5,-1476</points>
<connection>
<GID>743</GID>
<name>OUT_2</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-1510.5,-67,-1477</points>
<intersection>-1510.5 1</intersection>
<intersection>-1477 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,-1510.5,-54,-1510.5</points>
<connection>
<GID>2316</GID>
<name>IN_0</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1477,-67,-1477</points>
<connection>
<GID>743</GID>
<name>OUT_1</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>1391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,-1528,-68,-1478</points>
<intersection>-1528 1</intersection>
<intersection>-1478 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-1528,-54.5,-1528</points>
<connection>
<GID>2333</GID>
<name>IN_0</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-1478,-68,-1478</points>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection>
<intersection>-68 0</intersection></hsegment></shape></wire>
<wire>
<ID>1392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-1726.5,-16,-1720</points>
<intersection>-1726.5 1</intersection>
<intersection>-1720 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-1726.5,-13.5,-1726.5</points>
<connection>
<GID>2471</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17.5,-1720,-16,-1720</points>
<connection>
<GID>2470</GID>
<name>OUT_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>1393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-1727.5,33,-1720</points>
<intersection>-1727.5 1</intersection>
<intersection>-1720 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-1727.5,35,-1727.5</points>
<connection>
<GID>2473</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-1720,33,-1720</points>
<connection>
<GID>2472</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>1394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-1721,350.5,-1721</points>
<connection>
<GID>2486</GID>
<name>OUT</name></connection>
<intersection>-23.5 107</intersection>
<intersection>-15 4</intersection>
<intersection>26 108</intersection>
<intersection>33.5 16</intersection>
<intersection>74 109</intersection>
<intersection>81 23</intersection>
<intersection>123.5 110</intersection>
<intersection>131.5 31</intersection>
<intersection>171.5 111</intersection>
<intersection>180 55</intersection>
<intersection>229 112</intersection>
<intersection>238.5 56</intersection>
<intersection>284 113</intersection>
<intersection>292.5 66</intersection>
<intersection>341 114</intersection>
<intersection>350.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-15,-1728.5,-15,-1721</points>
<intersection>-1728.5 5</intersection>
<intersection>-1721 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-15,-1728.5,-13.5,-1728.5</points>
<connection>
<GID>2471</GID>
<name>IN_1</name></connection>
<intersection>-15 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>33.5,-1729.5,33.5,-1721</points>
<intersection>-1729.5 21</intersection>
<intersection>-1721 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>33.5,-1729.5,35,-1729.5</points>
<connection>
<GID>2473</GID>
<name>IN_1</name></connection>
<intersection>33.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>81,-1728.5,81,-1721</points>
<intersection>-1728.5 53</intersection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>131.5,-1728.5,131.5,-1721</points>
<intersection>-1728.5 115</intersection>
<intersection>-1721 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>81,-1728.5,81.5,-1728.5</points>
<connection>
<GID>2475</GID>
<name>IN_1</name></connection>
<intersection>81 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>180,-1728,180,-1721</points>
<connection>
<GID>2479</GID>
<name>IN_1</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>238.5,-1730,238.5,-1721</points>
<connection>
<GID>2481</GID>
<name>IN_1</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>292.5,-1729,292.5,-1721</points>
<intersection>-1729 118</intersection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>350.5,-1729.5,350.5,-1721</points>
<connection>
<GID>2485</GID>
<name>IN_1</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-23.5,-1723,-23.5,-1721</points>
<connection>
<GID>2470</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>26,-1723,26,-1721</points>
<connection>
<GID>2472</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>74,-1723,74,-1721</points>
<connection>
<GID>2474</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>123.5,-1723,123.5,-1721</points>
<connection>
<GID>2476</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>171.5,-1723,171.5,-1721</points>
<connection>
<GID>2478</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>229,-1723,229,-1721</points>
<connection>
<GID>2480</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>284,-1723,284,-1721</points>
<connection>
<GID>2482</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>341,-1723,341,-1721</points>
<connection>
<GID>2484</GID>
<name>clock</name></connection>
<intersection>-1721 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>131.5,-1728.5,132,-1728.5</points>
<connection>
<GID>2477</GID>
<name>IN_1</name></connection>
<intersection>131.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>292,-1729,292.5,-1729</points>
<connection>
<GID>2483</GID>
<name>IN_1</name></connection>
<intersection>292.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-1726.5,81.5,-1720</points>
<connection>
<GID>2475</GID>
<name>IN_0</name></connection>
<intersection>-1720 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>80,-1720,81.5,-1720</points>
<connection>
<GID>2474</GID>
<name>OUT_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-1726.5,131,-1720</points>
<intersection>-1726.5 1</intersection>
<intersection>-1720 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-1726.5,132,-1726.5</points>
<connection>
<GID>2477</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129.5,-1720,131,-1720</points>
<connection>
<GID>2476</GID>
<name>OUT_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>1397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-1726,179.5,-1720</points>
<intersection>-1726 5</intersection>
<intersection>-1720 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177.5,-1720,179.5,-1720</points>
<connection>
<GID>2478</GID>
<name>OUT_0</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>179.5,-1726,180,-1726</points>
<connection>
<GID>2479</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-1728,238,-1720</points>
<intersection>-1728 1</intersection>
<intersection>-1720 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,-1728,238.5,-1728</points>
<connection>
<GID>2481</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235,-1720,238,-1720</points>
<connection>
<GID>2480</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>1399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-1727,291.5,-1720</points>
<intersection>-1727 4</intersection>
<intersection>-1720 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>290,-1720,291.5,-1720</points>
<connection>
<GID>2482</GID>
<name>OUT_0</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>291.5,-1727,292,-1727</points>
<connection>
<GID>2483</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-1727.5,350,-1720</points>
<intersection>-1727.5 1</intersection>
<intersection>-1720 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-1727.5,350.5,-1727.5</points>
<connection>
<GID>2485</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347,-1720,350,-1720</points>
<connection>
<GID>2484</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>1401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-1739.5,-16,-1733</points>
<intersection>-1739.5 1</intersection>
<intersection>-1733 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-1739.5,-13.5,-1739.5</points>
<connection>
<GID>2488</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17.5,-1733,-16,-1733</points>
<connection>
<GID>2487</GID>
<name>OUT_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>1402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-1740.5,33,-1733</points>
<intersection>-1740.5 1</intersection>
<intersection>-1733 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-1740.5,35,-1740.5</points>
<connection>
<GID>2490</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-1733,33,-1733</points>
<connection>
<GID>2489</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>1403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-1734,350.5,-1734</points>
<connection>
<GID>2503</GID>
<name>OUT</name></connection>
<intersection>-23.5 107</intersection>
<intersection>-15 4</intersection>
<intersection>26 108</intersection>
<intersection>33.5 16</intersection>
<intersection>74 109</intersection>
<intersection>81 23</intersection>
<intersection>123.5 110</intersection>
<intersection>131.5 31</intersection>
<intersection>171.5 111</intersection>
<intersection>180 55</intersection>
<intersection>229 112</intersection>
<intersection>238.5 56</intersection>
<intersection>284 113</intersection>
<intersection>292.5 66</intersection>
<intersection>341 114</intersection>
<intersection>350.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-15,-1741.5,-15,-1734</points>
<intersection>-1741.5 5</intersection>
<intersection>-1734 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-15,-1741.5,-13.5,-1741.5</points>
<connection>
<GID>2488</GID>
<name>IN_1</name></connection>
<intersection>-15 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>33.5,-1742.5,33.5,-1734</points>
<intersection>-1742.5 21</intersection>
<intersection>-1734 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>33.5,-1742.5,35,-1742.5</points>
<connection>
<GID>2490</GID>
<name>IN_1</name></connection>
<intersection>33.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>81,-1741.5,81,-1734</points>
<intersection>-1741.5 53</intersection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>131.5,-1741.5,131.5,-1734</points>
<intersection>-1741.5 115</intersection>
<intersection>-1734 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>81,-1741.5,81.5,-1741.5</points>
<connection>
<GID>2492</GID>
<name>IN_1</name></connection>
<intersection>81 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>180,-1741,180,-1734</points>
<connection>
<GID>2496</GID>
<name>IN_1</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>238.5,-1743,238.5,-1734</points>
<connection>
<GID>2498</GID>
<name>IN_1</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>292.5,-1742,292.5,-1734</points>
<intersection>-1742 118</intersection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>350.5,-1742.5,350.5,-1734</points>
<connection>
<GID>2502</GID>
<name>IN_1</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-23.5,-1736,-23.5,-1734</points>
<connection>
<GID>2487</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>26,-1736,26,-1734</points>
<connection>
<GID>2489</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>74,-1736,74,-1734</points>
<connection>
<GID>2491</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>123.5,-1736,123.5,-1734</points>
<connection>
<GID>2493</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>171.5,-1736,171.5,-1734</points>
<connection>
<GID>2495</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>229,-1736,229,-1734</points>
<connection>
<GID>2497</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>284,-1736,284,-1734</points>
<connection>
<GID>2499</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>341,-1736,341,-1734</points>
<connection>
<GID>2501</GID>
<name>clock</name></connection>
<intersection>-1734 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>131.5,-1741.5,132,-1741.5</points>
<connection>
<GID>2494</GID>
<name>IN_1</name></connection>
<intersection>131.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>292,-1742,292.5,-1742</points>
<connection>
<GID>2500</GID>
<name>IN_1</name></connection>
<intersection>292.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-1739.5,81.5,-1733</points>
<connection>
<GID>2492</GID>
<name>IN_0</name></connection>
<intersection>-1733 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>80,-1733,81.5,-1733</points>
<connection>
<GID>2491</GID>
<name>OUT_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-1739.5,131,-1733</points>
<intersection>-1739.5 1</intersection>
<intersection>-1733 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-1739.5,132,-1739.5</points>
<connection>
<GID>2494</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129.5,-1733,131,-1733</points>
<connection>
<GID>2493</GID>
<name>OUT_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>1406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-1739,179.5,-1733</points>
<intersection>-1739 5</intersection>
<intersection>-1733 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177.5,-1733,179.5,-1733</points>
<connection>
<GID>2495</GID>
<name>OUT_0</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>179.5,-1739,180,-1739</points>
<connection>
<GID>2496</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-1741,238,-1733</points>
<intersection>-1741 1</intersection>
<intersection>-1733 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,-1741,238.5,-1741</points>
<connection>
<GID>2498</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235,-1733,238,-1733</points>
<connection>
<GID>2497</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>1408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-1740,291.5,-1733</points>
<intersection>-1740 4</intersection>
<intersection>-1733 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>290,-1733,291.5,-1733</points>
<connection>
<GID>2499</GID>
<name>OUT_0</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>291.5,-1740,292,-1740</points>
<connection>
<GID>2500</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-1740.5,350,-1733</points>
<intersection>-1740.5 1</intersection>
<intersection>-1733 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-1740.5,350.5,-1740.5</points>
<connection>
<GID>2502</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347,-1733,350,-1733</points>
<connection>
<GID>2501</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>1410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-1754,-16,-1747.5</points>
<intersection>-1754 1</intersection>
<intersection>-1747.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-1754,-13.5,-1754</points>
<connection>
<GID>2505</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17.5,-1747.5,-16,-1747.5</points>
<connection>
<GID>2504</GID>
<name>OUT_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>1411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-1755,33,-1747.5</points>
<intersection>-1755 1</intersection>
<intersection>-1747.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-1755,35,-1755</points>
<connection>
<GID>2507</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-1747.5,33,-1747.5</points>
<connection>
<GID>2506</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>1412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-1748.5,350.5,-1748.5</points>
<connection>
<GID>2520</GID>
<name>OUT</name></connection>
<intersection>-23.5 107</intersection>
<intersection>-15 4</intersection>
<intersection>26 108</intersection>
<intersection>33.5 16</intersection>
<intersection>74 109</intersection>
<intersection>81 23</intersection>
<intersection>123.5 110</intersection>
<intersection>131.5 31</intersection>
<intersection>171.5 111</intersection>
<intersection>180 55</intersection>
<intersection>229 112</intersection>
<intersection>238.5 56</intersection>
<intersection>284 113</intersection>
<intersection>292.5 66</intersection>
<intersection>341 114</intersection>
<intersection>350.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-15,-1756,-15,-1748.5</points>
<intersection>-1756 5</intersection>
<intersection>-1748.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-15,-1756,-13.5,-1756</points>
<connection>
<GID>2505</GID>
<name>IN_1</name></connection>
<intersection>-15 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>33.5,-1757,33.5,-1748.5</points>
<intersection>-1757 21</intersection>
<intersection>-1748.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>33.5,-1757,35,-1757</points>
<connection>
<GID>2507</GID>
<name>IN_1</name></connection>
<intersection>33.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>81,-1756,81,-1748.5</points>
<intersection>-1756 53</intersection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>131.5,-1756,131.5,-1748.5</points>
<intersection>-1756 115</intersection>
<intersection>-1748.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>81,-1756,81.5,-1756</points>
<connection>
<GID>2509</GID>
<name>IN_1</name></connection>
<intersection>81 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>180,-1755.5,180,-1748.5</points>
<connection>
<GID>2513</GID>
<name>IN_1</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>238.5,-1757.5,238.5,-1748.5</points>
<connection>
<GID>2515</GID>
<name>IN_1</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>292.5,-1756.5,292.5,-1748.5</points>
<intersection>-1756.5 118</intersection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>350.5,-1757,350.5,-1748.5</points>
<connection>
<GID>2519</GID>
<name>IN_1</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-23.5,-1750.5,-23.5,-1748.5</points>
<connection>
<GID>2504</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>26,-1750.5,26,-1748.5</points>
<connection>
<GID>2506</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>74,-1750.5,74,-1748.5</points>
<connection>
<GID>2508</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>123.5,-1750.5,123.5,-1748.5</points>
<connection>
<GID>2510</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>171.5,-1750.5,171.5,-1748.5</points>
<connection>
<GID>2512</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>229,-1750.5,229,-1748.5</points>
<connection>
<GID>2514</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>284,-1750.5,284,-1748.5</points>
<connection>
<GID>2516</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>341,-1750.5,341,-1748.5</points>
<connection>
<GID>2518</GID>
<name>clock</name></connection>
<intersection>-1748.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>131.5,-1756,132,-1756</points>
<connection>
<GID>2511</GID>
<name>IN_1</name></connection>
<intersection>131.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>292,-1756.5,292.5,-1756.5</points>
<connection>
<GID>2517</GID>
<name>IN_1</name></connection>
<intersection>292.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-1754,81.5,-1747.5</points>
<connection>
<GID>2509</GID>
<name>IN_0</name></connection>
<intersection>-1747.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>80,-1747.5,81.5,-1747.5</points>
<connection>
<GID>2508</GID>
<name>OUT_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-1754,131,-1747.5</points>
<intersection>-1754 1</intersection>
<intersection>-1747.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-1754,132,-1754</points>
<connection>
<GID>2511</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129.5,-1747.5,131,-1747.5</points>
<connection>
<GID>2510</GID>
<name>OUT_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>1415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-1753.5,179.5,-1747.5</points>
<intersection>-1753.5 5</intersection>
<intersection>-1747.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177.5,-1747.5,179.5,-1747.5</points>
<connection>
<GID>2512</GID>
<name>OUT_0</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>179.5,-1753.5,180,-1753.5</points>
<connection>
<GID>2513</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-1755.5,238,-1747.5</points>
<intersection>-1755.5 1</intersection>
<intersection>-1747.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,-1755.5,238.5,-1755.5</points>
<connection>
<GID>2515</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>235,-1747.5,238,-1747.5</points>
<connection>
<GID>2514</GID>
<name>OUT_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>1417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-1754.5,291.5,-1747.5</points>
<intersection>-1754.5 4</intersection>
<intersection>-1747.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>290,-1747.5,291.5,-1747.5</points>
<connection>
<GID>2516</GID>
<name>OUT_0</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>291.5,-1754.5,292,-1754.5</points>
<connection>
<GID>2517</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-1755,350,-1747.5</points>
<intersection>-1755 1</intersection>
<intersection>-1747.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-1755,350.5,-1755</points>
<connection>
<GID>2519</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347,-1747.5,350,-1747.5</points>
<connection>
<GID>2518</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>1419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-1766.5,-16.5,-1760</points>
<intersection>-1766.5 1</intersection>
<intersection>-1760 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-1766.5,-14,-1766.5</points>
<connection>
<GID>2522</GID>
<name>IN_0</name></connection>
<intersection>-16.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-18,-1760,-16.5,-1760</points>
<connection>
<GID>2521</GID>
<name>OUT_0</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-1767.5,32.5,-1760</points>
<intersection>-1767.5 1</intersection>
<intersection>-1760 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-1767.5,34.5,-1767.5</points>
<connection>
<GID>2524</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-1760,32.5,-1760</points>
<connection>
<GID>2523</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49.5,-1761,350,-1761</points>
<connection>
<GID>2537</GID>
<name>OUT</name></connection>
<intersection>-24 107</intersection>
<intersection>-15.5 4</intersection>
<intersection>25.5 108</intersection>
<intersection>33 16</intersection>
<intersection>73.5 109</intersection>
<intersection>80.5 23</intersection>
<intersection>123 110</intersection>
<intersection>131 31</intersection>
<intersection>171 111</intersection>
<intersection>179.5 55</intersection>
<intersection>228.5 112</intersection>
<intersection>238 56</intersection>
<intersection>283.5 113</intersection>
<intersection>292 66</intersection>
<intersection>340.5 114</intersection>
<intersection>350 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-15.5,-1768.5,-15.5,-1761</points>
<intersection>-1768.5 5</intersection>
<intersection>-1761 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-15.5,-1768.5,-14,-1768.5</points>
<connection>
<GID>2522</GID>
<name>IN_1</name></connection>
<intersection>-15.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>33,-1769.5,33,-1761</points>
<intersection>-1769.5 21</intersection>
<intersection>-1761 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>33,-1769.5,34.5,-1769.5</points>
<connection>
<GID>2524</GID>
<name>IN_1</name></connection>
<intersection>33 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>80.5,-1768.5,80.5,-1761</points>
<intersection>-1768.5 53</intersection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>131,-1768.5,131,-1761</points>
<intersection>-1768.5 115</intersection>
<intersection>-1761 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>80.5,-1768.5,81,-1768.5</points>
<connection>
<GID>2526</GID>
<name>IN_1</name></connection>
<intersection>80.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>179.5,-1768,179.5,-1761</points>
<connection>
<GID>2530</GID>
<name>IN_1</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>238,-1770,238,-1761</points>
<connection>
<GID>2532</GID>
<name>IN_1</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>292,-1769,292,-1761</points>
<intersection>-1769 118</intersection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>350,-1769.5,350,-1761</points>
<connection>
<GID>2536</GID>
<name>IN_1</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-24,-1763,-24,-1761</points>
<connection>
<GID>2521</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>25.5,-1763,25.5,-1761</points>
<connection>
<GID>2523</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>73.5,-1763,73.5,-1761</points>
<connection>
<GID>2525</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>123,-1763,123,-1761</points>
<connection>
<GID>2527</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>171,-1763,171,-1761</points>
<connection>
<GID>2529</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>228.5,-1763,228.5,-1761</points>
<connection>
<GID>2531</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>283.5,-1763,283.5,-1761</points>
<connection>
<GID>2533</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>340.5,-1763,340.5,-1761</points>
<connection>
<GID>2535</GID>
<name>clock</name></connection>
<intersection>-1761 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>131,-1768.5,131.5,-1768.5</points>
<connection>
<GID>2528</GID>
<name>IN_1</name></connection>
<intersection>131 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>291.5,-1769,292,-1769</points>
<connection>
<GID>2534</GID>
<name>IN_1</name></connection>
<intersection>292 66</intersection></hsegment></shape></wire>
<wire>
<ID>1422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-1766.5,81,-1760</points>
<connection>
<GID>2526</GID>
<name>IN_0</name></connection>
<intersection>-1760 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79.5,-1760,81,-1760</points>
<connection>
<GID>2525</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>1423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-1766.5,130.5,-1760</points>
<intersection>-1766.5 1</intersection>
<intersection>-1760 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-1766.5,131.5,-1766.5</points>
<connection>
<GID>2528</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129,-1760,130.5,-1760</points>
<connection>
<GID>2527</GID>
<name>OUT_0</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-1766,179,-1760</points>
<intersection>-1766 5</intersection>
<intersection>-1760 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177,-1760,179,-1760</points>
<connection>
<GID>2529</GID>
<name>OUT_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>179,-1766,179.5,-1766</points>
<connection>
<GID>2530</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment></shape></wire>
<wire>
<ID>1425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-1768,237.5,-1760</points>
<intersection>-1768 1</intersection>
<intersection>-1760 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>237.5,-1768,238,-1768</points>
<connection>
<GID>2532</GID>
<name>IN_0</name></connection>
<intersection>237.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234.5,-1760,237.5,-1760</points>
<connection>
<GID>2531</GID>
<name>OUT_0</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-1767,291,-1760</points>
<intersection>-1767 4</intersection>
<intersection>-1760 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289.5,-1760,291,-1760</points>
<connection>
<GID>2533</GID>
<name>OUT_0</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>291,-1767,291.5,-1767</points>
<connection>
<GID>2534</GID>
<name>IN_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>1427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-1767.5,349.5,-1760</points>
<intersection>-1767.5 1</intersection>
<intersection>-1760 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349.5,-1767.5,350,-1767.5</points>
<connection>
<GID>2536</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346.5,-1760,349.5,-1760</points>
<connection>
<GID>2535</GID>
<name>OUT_0</name></connection>
<intersection>349.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-1779.5,-17,-1773</points>
<intersection>-1779.5 1</intersection>
<intersection>-1773 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-1779.5,-14.5,-1779.5</points>
<connection>
<GID>2539</GID>
<name>IN_0</name></connection>
<intersection>-17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-18.5,-1773,-17,-1773</points>
<connection>
<GID>2538</GID>
<name>OUT_0</name></connection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>1429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-1780.5,32,-1773</points>
<intersection>-1780.5 1</intersection>
<intersection>-1773 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-1780.5,34,-1780.5</points>
<connection>
<GID>2541</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-1773,32,-1773</points>
<connection>
<GID>2540</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>1430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50,-1774,349.5,-1774</points>
<connection>
<GID>2554</GID>
<name>OUT</name></connection>
<intersection>-24.5 107</intersection>
<intersection>-16 4</intersection>
<intersection>25 108</intersection>
<intersection>32.5 16</intersection>
<intersection>73 109</intersection>
<intersection>80 23</intersection>
<intersection>122.5 110</intersection>
<intersection>130.5 31</intersection>
<intersection>170.5 111</intersection>
<intersection>179 55</intersection>
<intersection>228 112</intersection>
<intersection>237.5 56</intersection>
<intersection>283 113</intersection>
<intersection>291.5 66</intersection>
<intersection>340 114</intersection>
<intersection>349.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-16,-1781.5,-16,-1774</points>
<intersection>-1781.5 5</intersection>
<intersection>-1774 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-16,-1781.5,-14.5,-1781.5</points>
<connection>
<GID>2539</GID>
<name>IN_1</name></connection>
<intersection>-16 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>32.5,-1782.5,32.5,-1774</points>
<intersection>-1782.5 21</intersection>
<intersection>-1774 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>32.5,-1782.5,34,-1782.5</points>
<connection>
<GID>2541</GID>
<name>IN_1</name></connection>
<intersection>32.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>80,-1781.5,80,-1774</points>
<intersection>-1781.5 53</intersection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>130.5,-1781.5,130.5,-1774</points>
<intersection>-1781.5 115</intersection>
<intersection>-1774 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>80,-1781.5,80.5,-1781.5</points>
<connection>
<GID>2543</GID>
<name>IN_1</name></connection>
<intersection>80 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>179,-1781,179,-1774</points>
<connection>
<GID>2547</GID>
<name>IN_1</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>237.5,-1783,237.5,-1774</points>
<connection>
<GID>2549</GID>
<name>IN_1</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>291.5,-1782,291.5,-1774</points>
<intersection>-1782 118</intersection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>349.5,-1782.5,349.5,-1774</points>
<connection>
<GID>2553</GID>
<name>IN_1</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-24.5,-1776,-24.5,-1774</points>
<connection>
<GID>2538</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>25,-1776,25,-1774</points>
<connection>
<GID>2540</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>73,-1776,73,-1774</points>
<connection>
<GID>2542</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>122.5,-1776,122.5,-1774</points>
<connection>
<GID>2544</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>170.5,-1776,170.5,-1774</points>
<connection>
<GID>2546</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>228,-1776,228,-1774</points>
<connection>
<GID>2548</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>283,-1776,283,-1774</points>
<connection>
<GID>2550</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>340,-1776,340,-1774</points>
<connection>
<GID>2552</GID>
<name>clock</name></connection>
<intersection>-1774 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>130.5,-1781.5,131,-1781.5</points>
<connection>
<GID>2545</GID>
<name>IN_1</name></connection>
<intersection>130.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>291,-1782,291.5,-1782</points>
<connection>
<GID>2551</GID>
<name>IN_1</name></connection>
<intersection>291.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-1779.5,80.5,-1773</points>
<connection>
<GID>2543</GID>
<name>IN_0</name></connection>
<intersection>-1773 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1773,80.5,-1773</points>
<connection>
<GID>2542</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-1779.5,130,-1773</points>
<intersection>-1779.5 1</intersection>
<intersection>-1773 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-1779.5,131,-1779.5</points>
<connection>
<GID>2545</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>128.5,-1773,130,-1773</points>
<connection>
<GID>2544</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>1433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-1779,178.5,-1773</points>
<intersection>-1779 5</intersection>
<intersection>-1773 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>176.5,-1773,178.5,-1773</points>
<connection>
<GID>2546</GID>
<name>OUT_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>178.5,-1779,179,-1779</points>
<connection>
<GID>2547</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-1781,237,-1773</points>
<intersection>-1781 1</intersection>
<intersection>-1773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>237,-1781,237.5,-1781</points>
<connection>
<GID>2549</GID>
<name>IN_0</name></connection>
<intersection>237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,-1773,237,-1773</points>
<connection>
<GID>2548</GID>
<name>OUT_0</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>1435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-1780,290.5,-1773</points>
<intersection>-1780 4</intersection>
<intersection>-1773 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-1773,290.5,-1773</points>
<connection>
<GID>2550</GID>
<name>OUT_0</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>290.5,-1780,291,-1780</points>
<connection>
<GID>2551</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,-1780.5,349,-1773</points>
<intersection>-1780.5 1</intersection>
<intersection>-1773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349,-1780.5,349.5,-1780.5</points>
<connection>
<GID>2553</GID>
<name>IN_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346,-1773,349,-1773</points>
<connection>
<GID>2552</GID>
<name>OUT_0</name></connection>
<intersection>349 0</intersection></hsegment></shape></wire>
<wire>
<ID>1437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-1794.5,-17,-1788</points>
<intersection>-1794.5 1</intersection>
<intersection>-1788 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-1794.5,-14.5,-1794.5</points>
<connection>
<GID>2420</GID>
<name>IN_0</name></connection>
<intersection>-17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-18.5,-1788,-17,-1788</points>
<connection>
<GID>2419</GID>
<name>OUT_0</name></connection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>1438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-1795.5,32,-1788</points>
<intersection>-1795.5 1</intersection>
<intersection>-1788 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-1795.5,34,-1795.5</points>
<connection>
<GID>2422</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-1788,32,-1788</points>
<connection>
<GID>2421</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>1439</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50,-1789,349.5,-1789</points>
<connection>
<GID>2435</GID>
<name>OUT</name></connection>
<intersection>-24.5 107</intersection>
<intersection>-16 4</intersection>
<intersection>25 108</intersection>
<intersection>32.5 16</intersection>
<intersection>73 109</intersection>
<intersection>80 23</intersection>
<intersection>122.5 110</intersection>
<intersection>130.5 31</intersection>
<intersection>170.5 111</intersection>
<intersection>179 55</intersection>
<intersection>228 112</intersection>
<intersection>237.5 56</intersection>
<intersection>283 113</intersection>
<intersection>291.5 66</intersection>
<intersection>340 114</intersection>
<intersection>349.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-16,-1796.5,-16,-1789</points>
<intersection>-1796.5 5</intersection>
<intersection>-1789 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-16,-1796.5,-14.5,-1796.5</points>
<connection>
<GID>2420</GID>
<name>IN_1</name></connection>
<intersection>-16 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>32.5,-1797.5,32.5,-1789</points>
<intersection>-1797.5 21</intersection>
<intersection>-1789 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>32.5,-1797.5,34,-1797.5</points>
<connection>
<GID>2422</GID>
<name>IN_1</name></connection>
<intersection>32.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>80,-1796.5,80,-1789</points>
<intersection>-1796.5 53</intersection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>130.5,-1796.5,130.5,-1789</points>
<intersection>-1796.5 115</intersection>
<intersection>-1789 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>80,-1796.5,80.5,-1796.5</points>
<connection>
<GID>2424</GID>
<name>IN_1</name></connection>
<intersection>80 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>179,-1796,179,-1789</points>
<connection>
<GID>2428</GID>
<name>IN_1</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>237.5,-1798,237.5,-1789</points>
<connection>
<GID>2430</GID>
<name>IN_1</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>291.5,-1797,291.5,-1789</points>
<intersection>-1797 118</intersection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>349.5,-1797.5,349.5,-1789</points>
<connection>
<GID>2434</GID>
<name>IN_1</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-24.5,-1791,-24.5,-1789</points>
<connection>
<GID>2419</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>25,-1791,25,-1789</points>
<connection>
<GID>2421</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>73,-1791,73,-1789</points>
<connection>
<GID>2423</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>122.5,-1791,122.5,-1789</points>
<connection>
<GID>2425</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>170.5,-1791,170.5,-1789</points>
<connection>
<GID>2427</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>228,-1791,228,-1789</points>
<connection>
<GID>2429</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>283,-1791,283,-1789</points>
<connection>
<GID>2431</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>340,-1791,340,-1789</points>
<connection>
<GID>2433</GID>
<name>clock</name></connection>
<intersection>-1789 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>130.5,-1796.5,131,-1796.5</points>
<connection>
<GID>2426</GID>
<name>IN_1</name></connection>
<intersection>130.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>291,-1797,291.5,-1797</points>
<connection>
<GID>2432</GID>
<name>IN_1</name></connection>
<intersection>291.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-1794.5,80.5,-1788</points>
<connection>
<GID>2424</GID>
<name>IN_0</name></connection>
<intersection>-1788 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1788,80.5,-1788</points>
<connection>
<GID>2423</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-266,-1329,-94,-1329</points>
<connection>
<GID>1152</GID>
<name>OUT_0</name></connection>
<intersection>-204 23</intersection>
<intersection>-94 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-94,-2068.5,-94,-328</points>
<intersection>-2068.5 20</intersection>
<intersection>-1770.5 25</intersection>
<intersection>-1476 18</intersection>
<intersection>-1329 1</intersection>
<intersection>-1239.5 16</intersection>
<intersection>-922 15</intersection>
<intersection>-623 13</intersection>
<intersection>-328 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-94,-328,-84.5,-328</points>
<connection>
<GID>195</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-94,-623,-92,-623</points>
<connection>
<GID>332</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-94,-922,-85,-922</points>
<connection>
<GID>469</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-94,-1239.5,-92,-1239.5</points>
<connection>
<GID>606</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-94,-1476,-88.5,-1476</points>
<connection>
<GID>743</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-94,-2068.5,-89.5,-2068.5</points>
<connection>
<GID>1017</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-204,-1329,-204,-89.5</points>
<intersection>-1329 1</intersection>
<intersection>-89.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-204,-89.5,-88,-89.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>-204 23</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-94,-1770.5,-92.5,-1770.5</points>
<connection>
<GID>880</GID>
<name>IN_2</name></connection>
<intersection>-94 9</intersection></hsegment></shape></wire>
<wire>
<ID>1441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-1794.5,130,-1788</points>
<intersection>-1794.5 1</intersection>
<intersection>-1788 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-1794.5,131,-1794.5</points>
<connection>
<GID>2426</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>128.5,-1788,130,-1788</points>
<connection>
<GID>2425</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>1442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-1794,178.5,-1788</points>
<intersection>-1794 5</intersection>
<intersection>-1788 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>176.5,-1788,178.5,-1788</points>
<connection>
<GID>2427</GID>
<name>OUT_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>178.5,-1794,179,-1794</points>
<connection>
<GID>2428</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-266,-1322.5,-202,-1322.5</points>
<connection>
<GID>1154</GID>
<name>OUT_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-202,-2070.5,-202,-91.5</points>
<intersection>-2070.5 17</intersection>
<intersection>-1772.5 15</intersection>
<intersection>-1478 13</intersection>
<intersection>-1322.5 1</intersection>
<intersection>-1241.5 11</intersection>
<intersection>-924 9</intersection>
<intersection>-625 7</intersection>
<intersection>-330 5</intersection>
<intersection>-91.5 18</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-202,-330,-84.5,-330</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-202,-625,-92,-625</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-202,-924,-85,-924</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-202,-1241.5,-92,-1241.5</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-202,-1478,-88.5,-1478</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-202,-1772.5,-92.5,-1772.5</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-202,-2070.5,-89.5,-2070.5</points>
<connection>
<GID>1017</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-202,-91.5,-88,-91.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-202 3</intersection></hsegment></shape></wire>
<wire>
<ID>1443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-1796,237,-1788</points>
<intersection>-1796 1</intersection>
<intersection>-1788 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>237,-1796,237.5,-1796</points>
<connection>
<GID>2430</GID>
<name>IN_0</name></connection>
<intersection>237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,-1788,237,-1788</points>
<connection>
<GID>2429</GID>
<name>OUT_0</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-203,-2069.5,-203,-90.5</points>
<intersection>-2069.5 16</intersection>
<intersection>-1771.5 14</intersection>
<intersection>-1477 12</intersection>
<intersection>-1325.5 2</intersection>
<intersection>-1240.5 10</intersection>
<intersection>-923 8</intersection>
<intersection>-624 6</intersection>
<intersection>-329 1</intersection>
<intersection>-90.5 18</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-203,-329,-84.5,-329</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-266,-1325.5,-203,-1325.5</points>
<connection>
<GID>1153</GID>
<name>OUT_0</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-203,-624,-92,-624</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-203,-923,-85,-923</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-203,-1240.5,-92,-1240.5</points>
<connection>
<GID>606</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-203,-1477,-88.5,-1477</points>
<connection>
<GID>743</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-203,-1771.5,-92.5,-1771.5</points>
<connection>
<GID>880</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-203,-2069.5,-89.5,-2069.5</points>
<connection>
<GID>1017</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-203,-90.5,-88,-90.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment></shape></wire>
<wire>
<ID>1444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-1795,290.5,-1788</points>
<intersection>-1795 4</intersection>
<intersection>-1788 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-1788,290.5,-1788</points>
<connection>
<GID>2431</GID>
<name>OUT_0</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>290.5,-1795,291,-1795</points>
<connection>
<GID>2432</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,-1795.5,349,-1788</points>
<intersection>-1795.5 1</intersection>
<intersection>-1788 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349,-1795.5,349.5,-1795.5</points>
<connection>
<GID>2434</GID>
<name>IN_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346,-1788,349,-1788</points>
<connection>
<GID>2433</GID>
<name>OUT_0</name></connection>
<intersection>349 0</intersection></hsegment></shape></wire>
<wire>
<ID>1446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-1808.5,-17,-1802</points>
<intersection>-1808.5 1</intersection>
<intersection>-1802 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-1808.5,-14.5,-1808.5</points>
<connection>
<GID>2437</GID>
<name>IN_0</name></connection>
<intersection>-17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-18.5,-1802,-17,-1802</points>
<connection>
<GID>2436</GID>
<name>OUT_0</name></connection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>1447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-1809.5,32,-1802</points>
<intersection>-1809.5 1</intersection>
<intersection>-1802 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-1809.5,34,-1809.5</points>
<connection>
<GID>2439</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-1802,32,-1802</points>
<connection>
<GID>2438</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>1448</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50,-1803,349.5,-1803</points>
<connection>
<GID>2452</GID>
<name>OUT</name></connection>
<intersection>-24.5 107</intersection>
<intersection>-16 4</intersection>
<intersection>25 108</intersection>
<intersection>32.5 16</intersection>
<intersection>73 109</intersection>
<intersection>80 23</intersection>
<intersection>122.5 110</intersection>
<intersection>130.5 31</intersection>
<intersection>170.5 111</intersection>
<intersection>179 55</intersection>
<intersection>228 112</intersection>
<intersection>237.5 56</intersection>
<intersection>283 113</intersection>
<intersection>291.5 66</intersection>
<intersection>340 114</intersection>
<intersection>349.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-16,-1810.5,-16,-1803</points>
<intersection>-1810.5 5</intersection>
<intersection>-1803 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-16,-1810.5,-14.5,-1810.5</points>
<connection>
<GID>2437</GID>
<name>IN_1</name></connection>
<intersection>-16 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>32.5,-1811.5,32.5,-1803</points>
<intersection>-1811.5 21</intersection>
<intersection>-1803 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>32.5,-1811.5,34,-1811.5</points>
<connection>
<GID>2439</GID>
<name>IN_1</name></connection>
<intersection>32.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>80,-1810.5,80,-1803</points>
<intersection>-1810.5 53</intersection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>130.5,-1810.5,130.5,-1803</points>
<intersection>-1810.5 115</intersection>
<intersection>-1803 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>80,-1810.5,80.5,-1810.5</points>
<connection>
<GID>2441</GID>
<name>IN_1</name></connection>
<intersection>80 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>179,-1810,179,-1803</points>
<connection>
<GID>2445</GID>
<name>IN_1</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>237.5,-1812,237.5,-1803</points>
<connection>
<GID>2447</GID>
<name>IN_1</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>291.5,-1811,291.5,-1803</points>
<intersection>-1811 118</intersection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>349.5,-1811.5,349.5,-1803</points>
<connection>
<GID>2451</GID>
<name>IN_1</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-24.5,-1805,-24.5,-1803</points>
<connection>
<GID>2436</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>25,-1805,25,-1803</points>
<connection>
<GID>2438</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>73,-1805,73,-1803</points>
<connection>
<GID>2440</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>122.5,-1805,122.5,-1803</points>
<connection>
<GID>2442</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>170.5,-1805,170.5,-1803</points>
<connection>
<GID>2444</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>228,-1805,228,-1803</points>
<connection>
<GID>2446</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>283,-1805,283,-1803</points>
<connection>
<GID>2448</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>340,-1805,340,-1803</points>
<connection>
<GID>2450</GID>
<name>clock</name></connection>
<intersection>-1803 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>130.5,-1810.5,131,-1810.5</points>
<connection>
<GID>2443</GID>
<name>IN_1</name></connection>
<intersection>130.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>291,-1811,291.5,-1811</points>
<connection>
<GID>2449</GID>
<name>IN_1</name></connection>
<intersection>291.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-1808.5,80.5,-1802</points>
<connection>
<GID>2441</GID>
<name>IN_0</name></connection>
<intersection>-1802 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-1802,80.5,-1802</points>
<connection>
<GID>2440</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-1808.5,130,-1802</points>
<intersection>-1808.5 1</intersection>
<intersection>-1802 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-1808.5,131,-1808.5</points>
<connection>
<GID>2443</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>128.5,-1802,130,-1802</points>
<connection>
<GID>2442</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>1451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-1808,178.5,-1802</points>
<intersection>-1808 5</intersection>
<intersection>-1802 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>176.5,-1802,178.5,-1802</points>
<connection>
<GID>2444</GID>
<name>OUT_0</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>178.5,-1808,179,-1808</points>
<connection>
<GID>2445</GID>
<name>IN_0</name></connection>
<intersection>178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-1810,237,-1802</points>
<intersection>-1810 1</intersection>
<intersection>-1802 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>237,-1810,237.5,-1810</points>
<connection>
<GID>2447</GID>
<name>IN_0</name></connection>
<intersection>237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,-1802,237,-1802</points>
<connection>
<GID>2446</GID>
<name>OUT_0</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>1453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-1809,290.5,-1802</points>
<intersection>-1809 4</intersection>
<intersection>-1802 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,-1802,290.5,-1802</points>
<connection>
<GID>2448</GID>
<name>OUT_0</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>290.5,-1809,291,-1809</points>
<connection>
<GID>2449</GID>
<name>IN_0</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,-1809.5,349,-1802</points>
<intersection>-1809.5 1</intersection>
<intersection>-1802 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349,-1809.5,349.5,-1809.5</points>
<connection>
<GID>2451</GID>
<name>IN_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346,-1802,349,-1802</points>
<connection>
<GID>2450</GID>
<name>OUT_0</name></connection>
<intersection>349 0</intersection></hsegment></shape></wire>
<wire>
<ID>1455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-1826,-17.5,-1819.5</points>
<intersection>-1826 1</intersection>
<intersection>-1819.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-1826,-15,-1826</points>
<connection>
<GID>2454</GID>
<name>IN_0</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19,-1819.5,-17.5,-1819.5</points>
<connection>
<GID>2453</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-1827,31.5,-1819.5</points>
<intersection>-1827 1</intersection>
<intersection>-1819.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-1827,33.5,-1827</points>
<connection>
<GID>2456</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-1819.5,31.5,-1819.5</points>
<connection>
<GID>2455</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1457</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50.5,-1820.5,349,-1820.5</points>
<connection>
<GID>2469</GID>
<name>OUT</name></connection>
<intersection>-25 107</intersection>
<intersection>-16.5 4</intersection>
<intersection>24.5 108</intersection>
<intersection>32 16</intersection>
<intersection>72.5 109</intersection>
<intersection>79.5 23</intersection>
<intersection>122 110</intersection>
<intersection>130 31</intersection>
<intersection>170 111</intersection>
<intersection>178.5 55</intersection>
<intersection>227.5 112</intersection>
<intersection>237 56</intersection>
<intersection>282.5 113</intersection>
<intersection>291 66</intersection>
<intersection>339.5 114</intersection>
<intersection>349 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-16.5,-1828,-16.5,-1820.5</points>
<intersection>-1828 5</intersection>
<intersection>-1820.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-16.5,-1828,-15,-1828</points>
<connection>
<GID>2454</GID>
<name>IN_1</name></connection>
<intersection>-16.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>32,-1829,32,-1820.5</points>
<intersection>-1829 21</intersection>
<intersection>-1820.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>32,-1829,33.5,-1829</points>
<connection>
<GID>2456</GID>
<name>IN_1</name></connection>
<intersection>32 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>79.5,-1828,79.5,-1820.5</points>
<intersection>-1828 53</intersection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>130,-1828,130,-1820.5</points>
<intersection>-1828 115</intersection>
<intersection>-1820.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>79.5,-1828,80,-1828</points>
<connection>
<GID>2458</GID>
<name>IN_1</name></connection>
<intersection>79.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>178.5,-1827.5,178.5,-1820.5</points>
<connection>
<GID>2462</GID>
<name>IN_1</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>237,-1829.5,237,-1820.5</points>
<connection>
<GID>2464</GID>
<name>IN_1</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>291,-1828.5,291,-1820.5</points>
<intersection>-1828.5 118</intersection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>349,-1829,349,-1820.5</points>
<connection>
<GID>2468</GID>
<name>IN_1</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-25,-1822.5,-25,-1820.5</points>
<connection>
<GID>2453</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>24.5,-1822.5,24.5,-1820.5</points>
<connection>
<GID>2455</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>72.5,-1822.5,72.5,-1820.5</points>
<connection>
<GID>2457</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>122,-1822.5,122,-1820.5</points>
<connection>
<GID>2459</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>170,-1822.5,170,-1820.5</points>
<connection>
<GID>2461</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>227.5,-1822.5,227.5,-1820.5</points>
<connection>
<GID>2463</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>282.5,-1822.5,282.5,-1820.5</points>
<connection>
<GID>2465</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>339.5,-1822.5,339.5,-1820.5</points>
<connection>
<GID>2467</GID>
<name>clock</name></connection>
<intersection>-1820.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>130,-1828,130.5,-1828</points>
<connection>
<GID>2460</GID>
<name>IN_1</name></connection>
<intersection>130 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>290.5,-1828.5,291,-1828.5</points>
<connection>
<GID>2466</GID>
<name>IN_1</name></connection>
<intersection>291 66</intersection></hsegment></shape></wire>
<wire>
<ID>1458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-1826,80,-1819.5</points>
<connection>
<GID>2458</GID>
<name>IN_0</name></connection>
<intersection>-1819.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>78.5,-1819.5,80,-1819.5</points>
<connection>
<GID>2457</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>1459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-1826,129.5,-1819.5</points>
<intersection>-1826 1</intersection>
<intersection>-1819.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-1826,130.5,-1826</points>
<connection>
<GID>2460</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>128,-1819.5,129.5,-1819.5</points>
<connection>
<GID>2459</GID>
<name>OUT_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-1825.5,178,-1819.5</points>
<intersection>-1825.5 5</intersection>
<intersection>-1819.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>176,-1819.5,178,-1819.5</points>
<connection>
<GID>2461</GID>
<name>OUT_0</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>178,-1825.5,178.5,-1825.5</points>
<connection>
<GID>2462</GID>
<name>IN_0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>1461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,-1827.5,236.5,-1819.5</points>
<intersection>-1827.5 1</intersection>
<intersection>-1819.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,-1827.5,237,-1827.5</points>
<connection>
<GID>2464</GID>
<name>IN_0</name></connection>
<intersection>236.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233.5,-1819.5,236.5,-1819.5</points>
<connection>
<GID>2463</GID>
<name>OUT_0</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-1826.5,290,-1819.5</points>
<intersection>-1826.5 4</intersection>
<intersection>-1819.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>288.5,-1819.5,290,-1819.5</points>
<connection>
<GID>2465</GID>
<name>OUT_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>290,-1826.5,290.5,-1826.5</points>
<connection>
<GID>2466</GID>
<name>IN_0</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>1463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>348.5,-1827,348.5,-1819.5</points>
<intersection>-1827 1</intersection>
<intersection>-1819.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>348.5,-1827,349,-1827</points>
<connection>
<GID>2468</GID>
<name>IN_0</name></connection>
<intersection>348.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>345.5,-1819.5,348.5,-1819.5</points>
<connection>
<GID>2467</GID>
<name>OUT_0</name></connection>
<intersection>348.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,-1765.5,-72,-1720</points>
<intersection>-1765.5 2</intersection>
<intersection>-1720 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,-1720,-55,-1720</points>
<connection>
<GID>2486</GID>
<name>IN_0</name></connection>
<intersection>-72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1765.5,-72,-1765.5</points>
<connection>
<GID>880</GID>
<name>OUT_7</name></connection>
<intersection>-72 0</intersection></hsegment></shape></wire>
<wire>
<ID>1465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,-1766.5,-70.5,-1733</points>
<intersection>-1766.5 2</intersection>
<intersection>-1733 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70.5,-1733,-55,-1733</points>
<connection>
<GID>2503</GID>
<name>IN_0</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1766.5,-70.5,-1766.5</points>
<connection>
<GID>880</GID>
<name>OUT_6</name></connection>
<intersection>-70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-1767.5,-69,-1747.5</points>
<intersection>-1767.5 2</intersection>
<intersection>-1747.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-1747.5,-55,-1747.5</points>
<connection>
<GID>2520</GID>
<name>IN_0</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1767.5,-69,-1767.5</points>
<connection>
<GID>880</GID>
<name>OUT_5</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>1467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-1768.5,-67.5,-1760</points>
<intersection>-1768.5 2</intersection>
<intersection>-1760 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-1760,-55.5,-1760</points>
<connection>
<GID>2537</GID>
<name>IN_0</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1768.5,-67.5,-1768.5</points>
<connection>
<GID>880</GID>
<name>OUT_4</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-1773,-67.5,-1769.5</points>
<intersection>-1773 1</intersection>
<intersection>-1769.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-1773,-56,-1773</points>
<connection>
<GID>2554</GID>
<name>IN_0</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1769.5,-67.5,-1769.5</points>
<connection>
<GID>880</GID>
<name>OUT_3</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-1788,-69,-1770.5</points>
<intersection>-1788 1</intersection>
<intersection>-1770.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-1788,-56,-1788</points>
<connection>
<GID>2435</GID>
<name>IN_0</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1770.5,-69,-1770.5</points>
<connection>
<GID>880</GID>
<name>OUT_2</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>1470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,-1802,-71,-1771.5</points>
<intersection>-1802 1</intersection>
<intersection>-1771.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,-1802,-56,-1802</points>
<connection>
<GID>2452</GID>
<name>IN_0</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1771.5,-71,-1771.5</points>
<connection>
<GID>880</GID>
<name>OUT_1</name></connection>
<intersection>-71 0</intersection></hsegment></shape></wire>
<wire>
<ID>1471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,-1819.5,-72.5,-1772.5</points>
<intersection>-1819.5 1</intersection>
<intersection>-1772.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72.5,-1819.5,-56.5,-1819.5</points>
<connection>
<GID>2469</GID>
<name>IN_0</name></connection>
<intersection>-72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-1772.5,-72.5,-1772.5</points>
<connection>
<GID>880</GID>
<name>OUT_0</name></connection>
<intersection>-72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-2020,-11,-2013.5</points>
<intersection>-2020 1</intersection>
<intersection>-2013.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-2020,-8.5,-2020</points>
<connection>
<GID>2607</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12.5,-2013.5,-11,-2013.5</points>
<connection>
<GID>2606</GID>
<name>OUT_0</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>1473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-2021,38,-2013.5</points>
<intersection>-2021 1</intersection>
<intersection>-2013.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-2021,40,-2021</points>
<connection>
<GID>2609</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>37,-2013.5,38,-2013.5</points>
<connection>
<GID>2608</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>1474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44,-2014.5,355.5,-2014.5</points>
<connection>
<GID>2622</GID>
<name>OUT</name></connection>
<intersection>-18.5 107</intersection>
<intersection>-10 4</intersection>
<intersection>31 108</intersection>
<intersection>38.5 16</intersection>
<intersection>79 109</intersection>
<intersection>86 23</intersection>
<intersection>128.5 110</intersection>
<intersection>136.5 31</intersection>
<intersection>176.5 111</intersection>
<intersection>185 55</intersection>
<intersection>234 112</intersection>
<intersection>243.5 56</intersection>
<intersection>289 113</intersection>
<intersection>297.5 66</intersection>
<intersection>346 114</intersection>
<intersection>355.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-10,-2022,-10,-2014.5</points>
<intersection>-2022 5</intersection>
<intersection>-2014.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-10,-2022,-8.5,-2022</points>
<connection>
<GID>2607</GID>
<name>IN_1</name></connection>
<intersection>-10 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>38.5,-2023,38.5,-2014.5</points>
<intersection>-2023 21</intersection>
<intersection>-2014.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>38.5,-2023,40,-2023</points>
<connection>
<GID>2609</GID>
<name>IN_1</name></connection>
<intersection>38.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>86,-2022,86,-2014.5</points>
<intersection>-2022 53</intersection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>136.5,-2022,136.5,-2014.5</points>
<intersection>-2022 115</intersection>
<intersection>-2014.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>86,-2022,86.5,-2022</points>
<connection>
<GID>2611</GID>
<name>IN_1</name></connection>
<intersection>86 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>185,-2021.5,185,-2014.5</points>
<connection>
<GID>2615</GID>
<name>IN_1</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>243.5,-2023.5,243.5,-2014.5</points>
<connection>
<GID>2617</GID>
<name>IN_1</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>297.5,-2022.5,297.5,-2014.5</points>
<intersection>-2022.5 118</intersection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>355.5,-2023,355.5,-2014.5</points>
<connection>
<GID>2621</GID>
<name>IN_1</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-18.5,-2016.5,-18.5,-2014.5</points>
<connection>
<GID>2606</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>31,-2016.5,31,-2014.5</points>
<connection>
<GID>2608</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>79,-2016.5,79,-2014.5</points>
<connection>
<GID>2610</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>128.5,-2016.5,128.5,-2014.5</points>
<connection>
<GID>2612</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>176.5,-2016.5,176.5,-2014.5</points>
<connection>
<GID>2614</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>234,-2016.5,234,-2014.5</points>
<connection>
<GID>2616</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>289,-2016.5,289,-2014.5</points>
<connection>
<GID>2618</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>346,-2016.5,346,-2014.5</points>
<connection>
<GID>2620</GID>
<name>clock</name></connection>
<intersection>-2014.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>136.5,-2022,137,-2022</points>
<connection>
<GID>2613</GID>
<name>IN_1</name></connection>
<intersection>136.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>297,-2022.5,297.5,-2022.5</points>
<connection>
<GID>2619</GID>
<name>IN_1</name></connection>
<intersection>297.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-2020,86.5,-2013.5</points>
<connection>
<GID>2611</GID>
<name>IN_0</name></connection>
<intersection>-2013.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>85,-2013.5,86.5,-2013.5</points>
<connection>
<GID>2610</GID>
<name>OUT_0</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-2020,136,-2013.5</points>
<intersection>-2020 1</intersection>
<intersection>-2013.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-2020,137,-2020</points>
<connection>
<GID>2613</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>134.5,-2013.5,136,-2013.5</points>
<connection>
<GID>2612</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>1477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-2019.5,184.5,-2013.5</points>
<intersection>-2019.5 5</intersection>
<intersection>-2013.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>182.5,-2013.5,184.5,-2013.5</points>
<connection>
<GID>2614</GID>
<name>OUT_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>184.5,-2019.5,185,-2019.5</points>
<connection>
<GID>2615</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-2021.5,243,-2013.5</points>
<intersection>-2021.5 1</intersection>
<intersection>-2013.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-2021.5,243.5,-2021.5</points>
<connection>
<GID>2617</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>240,-2013.5,243,-2013.5</points>
<connection>
<GID>2616</GID>
<name>OUT_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>1479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-2020.5,296.5,-2013.5</points>
<intersection>-2020.5 4</intersection>
<intersection>-2013.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>295,-2013.5,296.5,-2013.5</points>
<connection>
<GID>2618</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>296.5,-2020.5,297,-2020.5</points>
<connection>
<GID>2619</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-2021,355,-2013.5</points>
<intersection>-2021 1</intersection>
<intersection>-2013.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-2021,355.5,-2021</points>
<connection>
<GID>2621</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-2013.5,355,-2013.5</points>
<connection>
<GID>2620</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>1481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-2033,-11,-2026.5</points>
<intersection>-2033 1</intersection>
<intersection>-2026.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-2033,-8.5,-2033</points>
<connection>
<GID>2624</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12.5,-2026.5,-11,-2026.5</points>
<connection>
<GID>2623</GID>
<name>OUT_0</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>1482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-2034,38,-2026.5</points>
<intersection>-2034 1</intersection>
<intersection>-2026.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-2034,40,-2034</points>
<connection>
<GID>2626</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>37,-2026.5,38,-2026.5</points>
<connection>
<GID>2625</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>1483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44,-2027.5,355.5,-2027.5</points>
<connection>
<GID>2639</GID>
<name>OUT</name></connection>
<intersection>-18.5 107</intersection>
<intersection>-10 4</intersection>
<intersection>31 108</intersection>
<intersection>38.5 16</intersection>
<intersection>79 109</intersection>
<intersection>86 23</intersection>
<intersection>128.5 110</intersection>
<intersection>136.5 31</intersection>
<intersection>176.5 111</intersection>
<intersection>185 55</intersection>
<intersection>234 112</intersection>
<intersection>243.5 56</intersection>
<intersection>289 113</intersection>
<intersection>297.5 66</intersection>
<intersection>346 114</intersection>
<intersection>355.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-10,-2035,-10,-2027.5</points>
<intersection>-2035 5</intersection>
<intersection>-2027.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-10,-2035,-8.5,-2035</points>
<connection>
<GID>2624</GID>
<name>IN_1</name></connection>
<intersection>-10 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>38.5,-2036,38.5,-2027.5</points>
<intersection>-2036 21</intersection>
<intersection>-2027.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>38.5,-2036,40,-2036</points>
<connection>
<GID>2626</GID>
<name>IN_1</name></connection>
<intersection>38.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>86,-2035,86,-2027.5</points>
<intersection>-2035 53</intersection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>136.5,-2035,136.5,-2027.5</points>
<intersection>-2035 115</intersection>
<intersection>-2027.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>86,-2035,86.5,-2035</points>
<connection>
<GID>2628</GID>
<name>IN_1</name></connection>
<intersection>86 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>185,-2034.5,185,-2027.5</points>
<connection>
<GID>2632</GID>
<name>IN_1</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>243.5,-2036.5,243.5,-2027.5</points>
<connection>
<GID>2634</GID>
<name>IN_1</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>297.5,-2035.5,297.5,-2027.5</points>
<intersection>-2035.5 118</intersection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>355.5,-2036,355.5,-2027.5</points>
<connection>
<GID>2638</GID>
<name>IN_1</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-18.5,-2029.5,-18.5,-2027.5</points>
<connection>
<GID>2623</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>31,-2029.5,31,-2027.5</points>
<connection>
<GID>2625</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>79,-2029.5,79,-2027.5</points>
<connection>
<GID>2627</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>128.5,-2029.5,128.5,-2027.5</points>
<connection>
<GID>2629</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>176.5,-2029.5,176.5,-2027.5</points>
<connection>
<GID>2631</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>234,-2029.5,234,-2027.5</points>
<connection>
<GID>2633</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>289,-2029.5,289,-2027.5</points>
<connection>
<GID>2635</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>346,-2029.5,346,-2027.5</points>
<connection>
<GID>2637</GID>
<name>clock</name></connection>
<intersection>-2027.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>136.5,-2035,137,-2035</points>
<connection>
<GID>2630</GID>
<name>IN_1</name></connection>
<intersection>136.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>297,-2035.5,297.5,-2035.5</points>
<connection>
<GID>2636</GID>
<name>IN_1</name></connection>
<intersection>297.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-2033,86.5,-2026.5</points>
<connection>
<GID>2628</GID>
<name>IN_0</name></connection>
<intersection>-2026.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>85,-2026.5,86.5,-2026.5</points>
<connection>
<GID>2627</GID>
<name>OUT_0</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-2033,136,-2026.5</points>
<intersection>-2033 1</intersection>
<intersection>-2026.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-2033,137,-2033</points>
<connection>
<GID>2630</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>134.5,-2026.5,136,-2026.5</points>
<connection>
<GID>2629</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>1486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-2032.5,184.5,-2026.5</points>
<intersection>-2032.5 5</intersection>
<intersection>-2026.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>182.5,-2026.5,184.5,-2026.5</points>
<connection>
<GID>2631</GID>
<name>OUT_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>184.5,-2032.5,185,-2032.5</points>
<connection>
<GID>2632</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-2034.5,243,-2026.5</points>
<intersection>-2034.5 1</intersection>
<intersection>-2026.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-2034.5,243.5,-2034.5</points>
<connection>
<GID>2634</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>240,-2026.5,243,-2026.5</points>
<connection>
<GID>2633</GID>
<name>OUT_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>1488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-2033.5,296.5,-2026.5</points>
<intersection>-2033.5 4</intersection>
<intersection>-2026.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>295,-2026.5,296.5,-2026.5</points>
<connection>
<GID>2635</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>296.5,-2033.5,297,-2033.5</points>
<connection>
<GID>2636</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-2034,355,-2026.5</points>
<intersection>-2034 1</intersection>
<intersection>-2026.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-2034,355.5,-2034</points>
<connection>
<GID>2638</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-2026.5,355,-2026.5</points>
<connection>
<GID>2637</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>1490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-2047.5,-11,-2041</points>
<intersection>-2047.5 1</intersection>
<intersection>-2041 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-2047.5,-8.5,-2047.5</points>
<connection>
<GID>2641</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12.5,-2041,-11,-2041</points>
<connection>
<GID>2640</GID>
<name>OUT_0</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>1491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-2048.5,38,-2041</points>
<intersection>-2048.5 1</intersection>
<intersection>-2041 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-2048.5,40,-2048.5</points>
<connection>
<GID>2643</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>37,-2041,38,-2041</points>
<connection>
<GID>2642</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>1492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44,-2042,355.5,-2042</points>
<connection>
<GID>2656</GID>
<name>OUT</name></connection>
<intersection>-18.5 107</intersection>
<intersection>-10 4</intersection>
<intersection>31 108</intersection>
<intersection>38.5 16</intersection>
<intersection>79 109</intersection>
<intersection>86 23</intersection>
<intersection>128.5 110</intersection>
<intersection>136.5 31</intersection>
<intersection>176.5 111</intersection>
<intersection>185 55</intersection>
<intersection>234 112</intersection>
<intersection>243.5 56</intersection>
<intersection>289 113</intersection>
<intersection>297.5 66</intersection>
<intersection>346 114</intersection>
<intersection>355.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-10,-2049.5,-10,-2042</points>
<intersection>-2049.5 5</intersection>
<intersection>-2042 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-10,-2049.5,-8.5,-2049.5</points>
<connection>
<GID>2641</GID>
<name>IN_1</name></connection>
<intersection>-10 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>38.5,-2050.5,38.5,-2042</points>
<intersection>-2050.5 21</intersection>
<intersection>-2042 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>38.5,-2050.5,40,-2050.5</points>
<connection>
<GID>2643</GID>
<name>IN_1</name></connection>
<intersection>38.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>86,-2049.5,86,-2042</points>
<intersection>-2049.5 53</intersection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>136.5,-2049.5,136.5,-2042</points>
<intersection>-2049.5 115</intersection>
<intersection>-2042 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>86,-2049.5,86.5,-2049.5</points>
<connection>
<GID>2645</GID>
<name>IN_1</name></connection>
<intersection>86 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>185,-2049,185,-2042</points>
<connection>
<GID>2649</GID>
<name>IN_1</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>243.5,-2051,243.5,-2042</points>
<connection>
<GID>2651</GID>
<name>IN_1</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>297.5,-2050,297.5,-2042</points>
<intersection>-2050 118</intersection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>355.5,-2050.5,355.5,-2042</points>
<connection>
<GID>2655</GID>
<name>IN_1</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-18.5,-2044,-18.5,-2042</points>
<connection>
<GID>2640</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>31,-2044,31,-2042</points>
<connection>
<GID>2642</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>79,-2044,79,-2042</points>
<connection>
<GID>2644</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>128.5,-2044,128.5,-2042</points>
<connection>
<GID>2646</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>176.5,-2044,176.5,-2042</points>
<connection>
<GID>2648</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>234,-2044,234,-2042</points>
<connection>
<GID>2650</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>289,-2044,289,-2042</points>
<connection>
<GID>2652</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>346,-2044,346,-2042</points>
<connection>
<GID>2654</GID>
<name>clock</name></connection>
<intersection>-2042 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>136.5,-2049.5,137,-2049.5</points>
<connection>
<GID>2647</GID>
<name>IN_1</name></connection>
<intersection>136.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>297,-2050,297.5,-2050</points>
<connection>
<GID>2653</GID>
<name>IN_1</name></connection>
<intersection>297.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-2047.5,86.5,-2041</points>
<connection>
<GID>2645</GID>
<name>IN_0</name></connection>
<intersection>-2041 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>85,-2041,86.5,-2041</points>
<connection>
<GID>2644</GID>
<name>OUT_0</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-2047.5,136,-2041</points>
<intersection>-2047.5 1</intersection>
<intersection>-2041 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-2047.5,137,-2047.5</points>
<connection>
<GID>2647</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>134.5,-2041,136,-2041</points>
<connection>
<GID>2646</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>1495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-2047,184.5,-2041</points>
<intersection>-2047 5</intersection>
<intersection>-2041 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>182.5,-2041,184.5,-2041</points>
<connection>
<GID>2648</GID>
<name>OUT_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>184.5,-2047,185,-2047</points>
<connection>
<GID>2649</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-2049,243,-2041</points>
<intersection>-2049 1</intersection>
<intersection>-2041 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-2049,243.5,-2049</points>
<connection>
<GID>2651</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>240,-2041,243,-2041</points>
<connection>
<GID>2650</GID>
<name>OUT_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>1497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-2048,296.5,-2041</points>
<intersection>-2048 4</intersection>
<intersection>-2041 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>295,-2041,296.5,-2041</points>
<connection>
<GID>2652</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>296.5,-2048,297,-2048</points>
<connection>
<GID>2653</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-2048.5,355,-2041</points>
<intersection>-2048.5 1</intersection>
<intersection>-2041 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-2048.5,355.5,-2048.5</points>
<connection>
<GID>2655</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-2041,355,-2041</points>
<connection>
<GID>2654</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>1499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-2060,-11.5,-2053.5</points>
<intersection>-2060 1</intersection>
<intersection>-2053.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-2060,-9,-2060</points>
<connection>
<GID>2658</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-13,-2053.5,-11.5,-2053.5</points>
<connection>
<GID>2657</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-2061,37.5,-2053.5</points>
<intersection>-2061 1</intersection>
<intersection>-2053.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-2061,39.5,-2061</points>
<connection>
<GID>2660</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-2053.5,37.5,-2053.5</points>
<connection>
<GID>2659</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44.5,-2054.5,355,-2054.5</points>
<connection>
<GID>2673</GID>
<name>OUT</name></connection>
<intersection>-19 107</intersection>
<intersection>-10.5 4</intersection>
<intersection>30.5 108</intersection>
<intersection>38 16</intersection>
<intersection>78.5 109</intersection>
<intersection>85.5 23</intersection>
<intersection>128 110</intersection>
<intersection>136 31</intersection>
<intersection>176 111</intersection>
<intersection>184.5 55</intersection>
<intersection>233.5 112</intersection>
<intersection>243 56</intersection>
<intersection>288.5 113</intersection>
<intersection>297 66</intersection>
<intersection>345.5 114</intersection>
<intersection>355 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-10.5,-2062,-10.5,-2054.5</points>
<intersection>-2062 5</intersection>
<intersection>-2054.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-10.5,-2062,-9,-2062</points>
<connection>
<GID>2658</GID>
<name>IN_1</name></connection>
<intersection>-10.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>38,-2063,38,-2054.5</points>
<intersection>-2063 21</intersection>
<intersection>-2054.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>38,-2063,39.5,-2063</points>
<connection>
<GID>2660</GID>
<name>IN_1</name></connection>
<intersection>38 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>85.5,-2062,85.5,-2054.5</points>
<intersection>-2062 53</intersection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>136,-2062,136,-2054.5</points>
<intersection>-2062 115</intersection>
<intersection>-2054.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>85.5,-2062,86,-2062</points>
<connection>
<GID>2662</GID>
<name>IN_1</name></connection>
<intersection>85.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>184.5,-2061.5,184.5,-2054.5</points>
<connection>
<GID>2666</GID>
<name>IN_1</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>243,-2063.5,243,-2054.5</points>
<connection>
<GID>2668</GID>
<name>IN_1</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>297,-2062.5,297,-2054.5</points>
<intersection>-2062.5 118</intersection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>355,-2063,355,-2054.5</points>
<connection>
<GID>2672</GID>
<name>IN_1</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-19,-2056.5,-19,-2054.5</points>
<connection>
<GID>2657</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>30.5,-2056.5,30.5,-2054.5</points>
<connection>
<GID>2659</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>78.5,-2056.5,78.5,-2054.5</points>
<connection>
<GID>2661</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>128,-2056.5,128,-2054.5</points>
<connection>
<GID>2663</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>176,-2056.5,176,-2054.5</points>
<connection>
<GID>2665</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>233.5,-2056.5,233.5,-2054.5</points>
<connection>
<GID>2667</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>288.5,-2056.5,288.5,-2054.5</points>
<connection>
<GID>2669</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>345.5,-2056.5,345.5,-2054.5</points>
<connection>
<GID>2671</GID>
<name>clock</name></connection>
<intersection>-2054.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>136,-2062,136.5,-2062</points>
<connection>
<GID>2664</GID>
<name>IN_1</name></connection>
<intersection>136 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>296.5,-2062.5,297,-2062.5</points>
<connection>
<GID>2670</GID>
<name>IN_1</name></connection>
<intersection>297 66</intersection></hsegment></shape></wire>
<wire>
<ID>1502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-2060,86,-2053.5</points>
<connection>
<GID>2662</GID>
<name>IN_0</name></connection>
<intersection>-2053.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-2053.5,86,-2053.5</points>
<connection>
<GID>2661</GID>
<name>OUT_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>1503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-2060,135.5,-2053.5</points>
<intersection>-2060 1</intersection>
<intersection>-2053.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-2060,136.5,-2060</points>
<connection>
<GID>2664</GID>
<name>IN_0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>134,-2053.5,135.5,-2053.5</points>
<connection>
<GID>2663</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-2059.5,184,-2053.5</points>
<intersection>-2059.5 5</intersection>
<intersection>-2053.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>182,-2053.5,184,-2053.5</points>
<connection>
<GID>2665</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>184,-2059.5,184.5,-2059.5</points>
<connection>
<GID>2666</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>1505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-2061.5,242.5,-2053.5</points>
<intersection>-2061.5 1</intersection>
<intersection>-2053.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242.5,-2061.5,243,-2061.5</points>
<connection>
<GID>2668</GID>
<name>IN_0</name></connection>
<intersection>242.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239.5,-2053.5,242.5,-2053.5</points>
<connection>
<GID>2667</GID>
<name>OUT_0</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-2060.5,296,-2053.5</points>
<intersection>-2060.5 4</intersection>
<intersection>-2053.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>294.5,-2053.5,296,-2053.5</points>
<connection>
<GID>2669</GID>
<name>OUT_0</name></connection>
<intersection>296 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>296,-2060.5,296.5,-2060.5</points>
<connection>
<GID>2670</GID>
<name>IN_0</name></connection>
<intersection>296 0</intersection></hsegment></shape></wire>
<wire>
<ID>1507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-2061,354.5,-2053.5</points>
<intersection>-2061 1</intersection>
<intersection>-2053.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354.5,-2061,355,-2061</points>
<connection>
<GID>2672</GID>
<name>IN_0</name></connection>
<intersection>354.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351.5,-2053.5,354.5,-2053.5</points>
<connection>
<GID>2671</GID>
<name>OUT_0</name></connection>
<intersection>354.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-2073,-12,-2066.5</points>
<intersection>-2073 1</intersection>
<intersection>-2066.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-2073,-9.5,-2073</points>
<connection>
<GID>2675</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-13.5,-2066.5,-12,-2066.5</points>
<connection>
<GID>2674</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>1509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-2074,37,-2066.5</points>
<intersection>-2074 1</intersection>
<intersection>-2066.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-2074,39,-2074</points>
<connection>
<GID>2677</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-2066.5,37,-2066.5</points>
<connection>
<GID>2676</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>1510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-2067.5,354.5,-2067.5</points>
<connection>
<GID>2690</GID>
<name>OUT</name></connection>
<intersection>-19.5 107</intersection>
<intersection>-11 4</intersection>
<intersection>30 108</intersection>
<intersection>37.5 16</intersection>
<intersection>78 109</intersection>
<intersection>85 23</intersection>
<intersection>127.5 110</intersection>
<intersection>135.5 31</intersection>
<intersection>175.5 111</intersection>
<intersection>184 55</intersection>
<intersection>233 112</intersection>
<intersection>242.5 56</intersection>
<intersection>288 113</intersection>
<intersection>296.5 66</intersection>
<intersection>345 114</intersection>
<intersection>354.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11,-2075,-11,-2067.5</points>
<intersection>-2075 5</intersection>
<intersection>-2067.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-11,-2075,-9.5,-2075</points>
<connection>
<GID>2675</GID>
<name>IN_1</name></connection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>37.5,-2076,37.5,-2067.5</points>
<intersection>-2076 21</intersection>
<intersection>-2067.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>37.5,-2076,39,-2076</points>
<connection>
<GID>2677</GID>
<name>IN_1</name></connection>
<intersection>37.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>85,-2075,85,-2067.5</points>
<intersection>-2075 53</intersection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>135.5,-2075,135.5,-2067.5</points>
<intersection>-2075 115</intersection>
<intersection>-2067.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>85,-2075,85.5,-2075</points>
<connection>
<GID>2679</GID>
<name>IN_1</name></connection>
<intersection>85 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>184,-2074.5,184,-2067.5</points>
<connection>
<GID>2683</GID>
<name>IN_1</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>242.5,-2076.5,242.5,-2067.5</points>
<connection>
<GID>2685</GID>
<name>IN_1</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>296.5,-2075.5,296.5,-2067.5</points>
<intersection>-2075.5 118</intersection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>354.5,-2076,354.5,-2067.5</points>
<connection>
<GID>2689</GID>
<name>IN_1</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-19.5,-2069.5,-19.5,-2067.5</points>
<connection>
<GID>2674</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>30,-2069.5,30,-2067.5</points>
<connection>
<GID>2676</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>78,-2069.5,78,-2067.5</points>
<connection>
<GID>2678</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>127.5,-2069.5,127.5,-2067.5</points>
<connection>
<GID>2680</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>175.5,-2069.5,175.5,-2067.5</points>
<connection>
<GID>2682</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>233,-2069.5,233,-2067.5</points>
<connection>
<GID>2684</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>288,-2069.5,288,-2067.5</points>
<connection>
<GID>2686</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>345,-2069.5,345,-2067.5</points>
<connection>
<GID>2688</GID>
<name>clock</name></connection>
<intersection>-2067.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>135.5,-2075,136,-2075</points>
<connection>
<GID>2681</GID>
<name>IN_1</name></connection>
<intersection>135.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>296,-2075.5,296.5,-2075.5</points>
<connection>
<GID>2687</GID>
<name>IN_1</name></connection>
<intersection>296.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-2073,85.5,-2066.5</points>
<connection>
<GID>2679</GID>
<name>IN_0</name></connection>
<intersection>-2066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-2066.5,85.5,-2066.5</points>
<connection>
<GID>2678</GID>
<name>OUT_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-2073,135,-2066.5</points>
<intersection>-2073 1</intersection>
<intersection>-2066.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-2073,136,-2073</points>
<connection>
<GID>2681</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133.5,-2066.5,135,-2066.5</points>
<connection>
<GID>2680</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>1513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2072.5,183.5,-2066.5</points>
<intersection>-2072.5 5</intersection>
<intersection>-2066.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>181.5,-2066.5,183.5,-2066.5</points>
<connection>
<GID>2682</GID>
<name>OUT_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>183.5,-2072.5,184,-2072.5</points>
<connection>
<GID>2683</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-2074.5,242,-2066.5</points>
<intersection>-2074.5 1</intersection>
<intersection>-2066.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-2074.5,242.5,-2074.5</points>
<connection>
<GID>2685</GID>
<name>IN_0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-2066.5,242,-2066.5</points>
<connection>
<GID>2684</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>1515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-2073.5,295.5,-2066.5</points>
<intersection>-2073.5 4</intersection>
<intersection>-2066.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>294,-2066.5,295.5,-2066.5</points>
<connection>
<GID>2686</GID>
<name>OUT_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>295.5,-2073.5,296,-2073.5</points>
<connection>
<GID>2687</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-2074,354,-2066.5</points>
<intersection>-2074 1</intersection>
<intersection>-2066.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-2074,354.5,-2074</points>
<connection>
<GID>2689</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-2066.5,354,-2066.5</points>
<connection>
<GID>2688</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment></shape></wire>
<wire>
<ID>1517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-2088,-12,-2081.5</points>
<intersection>-2088 1</intersection>
<intersection>-2081.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-2088,-9.5,-2088</points>
<connection>
<GID>2556</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-13.5,-2081.5,-12,-2081.5</points>
<connection>
<GID>2555</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>1518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-2089,37,-2081.5</points>
<intersection>-2089 1</intersection>
<intersection>-2081.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-2089,39,-2089</points>
<connection>
<GID>2558</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-2081.5,37,-2081.5</points>
<connection>
<GID>2557</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>1519</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-2082.5,354.5,-2082.5</points>
<connection>
<GID>2571</GID>
<name>OUT</name></connection>
<intersection>-19.5 107</intersection>
<intersection>-11 4</intersection>
<intersection>30 108</intersection>
<intersection>37.5 16</intersection>
<intersection>78 109</intersection>
<intersection>85 23</intersection>
<intersection>127.5 110</intersection>
<intersection>135.5 31</intersection>
<intersection>175.5 111</intersection>
<intersection>184 55</intersection>
<intersection>233 112</intersection>
<intersection>242.5 56</intersection>
<intersection>288 113</intersection>
<intersection>296.5 66</intersection>
<intersection>345 114</intersection>
<intersection>354.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11,-2090,-11,-2082.5</points>
<intersection>-2090 5</intersection>
<intersection>-2082.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-11,-2090,-9.5,-2090</points>
<connection>
<GID>2556</GID>
<name>IN_1</name></connection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>37.5,-2091,37.5,-2082.5</points>
<intersection>-2091 21</intersection>
<intersection>-2082.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>37.5,-2091,39,-2091</points>
<connection>
<GID>2558</GID>
<name>IN_1</name></connection>
<intersection>37.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>85,-2090,85,-2082.5</points>
<intersection>-2090 53</intersection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>135.5,-2090,135.5,-2082.5</points>
<intersection>-2090 115</intersection>
<intersection>-2082.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>85,-2090,85.5,-2090</points>
<connection>
<GID>2560</GID>
<name>IN_1</name></connection>
<intersection>85 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>184,-2089.5,184,-2082.5</points>
<connection>
<GID>2564</GID>
<name>IN_1</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>242.5,-2091.5,242.5,-2082.5</points>
<connection>
<GID>2566</GID>
<name>IN_1</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>296.5,-2090.5,296.5,-2082.5</points>
<intersection>-2090.5 118</intersection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>354.5,-2091,354.5,-2082.5</points>
<connection>
<GID>2570</GID>
<name>IN_1</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-19.5,-2084.5,-19.5,-2082.5</points>
<connection>
<GID>2555</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>30,-2084.5,30,-2082.5</points>
<connection>
<GID>2557</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>78,-2084.5,78,-2082.5</points>
<connection>
<GID>2559</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>127.5,-2084.5,127.5,-2082.5</points>
<connection>
<GID>2561</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>175.5,-2084.5,175.5,-2082.5</points>
<connection>
<GID>2563</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>233,-2084.5,233,-2082.5</points>
<connection>
<GID>2565</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>288,-2084.5,288,-2082.5</points>
<connection>
<GID>2567</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>345,-2084.5,345,-2082.5</points>
<connection>
<GID>2569</GID>
<name>clock</name></connection>
<intersection>-2082.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>135.5,-2090,136,-2090</points>
<connection>
<GID>2562</GID>
<name>IN_1</name></connection>
<intersection>135.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>296,-2090.5,296.5,-2090.5</points>
<connection>
<GID>2568</GID>
<name>IN_1</name></connection>
<intersection>296.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-2088,85.5,-2081.5</points>
<connection>
<GID>2560</GID>
<name>IN_0</name></connection>
<intersection>-2081.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-2081.5,85.5,-2081.5</points>
<connection>
<GID>2559</GID>
<name>OUT_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-2088,135,-2081.5</points>
<intersection>-2088 1</intersection>
<intersection>-2081.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-2088,136,-2088</points>
<connection>
<GID>2562</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133.5,-2081.5,135,-2081.5</points>
<connection>
<GID>2561</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>1522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2087.5,183.5,-2081.5</points>
<intersection>-2087.5 5</intersection>
<intersection>-2081.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>181.5,-2081.5,183.5,-2081.5</points>
<connection>
<GID>2563</GID>
<name>OUT_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>183.5,-2087.5,184,-2087.5</points>
<connection>
<GID>2564</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-2089.5,242,-2081.5</points>
<intersection>-2089.5 1</intersection>
<intersection>-2081.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-2089.5,242.5,-2089.5</points>
<connection>
<GID>2566</GID>
<name>IN_0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-2081.5,242,-2081.5</points>
<connection>
<GID>2565</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>1524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-2088.5,295.5,-2081.5</points>
<intersection>-2088.5 4</intersection>
<intersection>-2081.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>294,-2081.5,295.5,-2081.5</points>
<connection>
<GID>2567</GID>
<name>OUT_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>295.5,-2088.5,296,-2088.5</points>
<connection>
<GID>2568</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-2089,354,-2081.5</points>
<intersection>-2089 1</intersection>
<intersection>-2081.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-2089,354.5,-2089</points>
<connection>
<GID>2570</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-2081.5,354,-2081.5</points>
<connection>
<GID>2569</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment></shape></wire>
<wire>
<ID>1526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-2102,-12,-2095.5</points>
<intersection>-2102 1</intersection>
<intersection>-2095.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-2102,-9.5,-2102</points>
<connection>
<GID>2573</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-13.5,-2095.5,-12,-2095.5</points>
<connection>
<GID>2572</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>1527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-2103,37,-2095.5</points>
<intersection>-2103 1</intersection>
<intersection>-2095.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-2103,39,-2103</points>
<connection>
<GID>2575</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-2095.5,37,-2095.5</points>
<connection>
<GID>2574</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>1528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-2096.5,354.5,-2096.5</points>
<connection>
<GID>2588</GID>
<name>OUT</name></connection>
<intersection>-19.5 107</intersection>
<intersection>-11 4</intersection>
<intersection>30 108</intersection>
<intersection>37.5 16</intersection>
<intersection>78 109</intersection>
<intersection>85 23</intersection>
<intersection>127.5 110</intersection>
<intersection>135.5 31</intersection>
<intersection>175.5 111</intersection>
<intersection>184 55</intersection>
<intersection>233 112</intersection>
<intersection>242.5 56</intersection>
<intersection>288 113</intersection>
<intersection>296.5 66</intersection>
<intersection>345 114</intersection>
<intersection>354.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11,-2104,-11,-2096.5</points>
<intersection>-2104 5</intersection>
<intersection>-2096.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-11,-2104,-9.5,-2104</points>
<connection>
<GID>2573</GID>
<name>IN_1</name></connection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>37.5,-2105,37.5,-2096.5</points>
<intersection>-2105 21</intersection>
<intersection>-2096.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>37.5,-2105,39,-2105</points>
<connection>
<GID>2575</GID>
<name>IN_1</name></connection>
<intersection>37.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>85,-2104,85,-2096.5</points>
<intersection>-2104 53</intersection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>135.5,-2104,135.5,-2096.5</points>
<intersection>-2104 115</intersection>
<intersection>-2096.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>85,-2104,85.5,-2104</points>
<connection>
<GID>2577</GID>
<name>IN_1</name></connection>
<intersection>85 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>184,-2103.5,184,-2096.5</points>
<connection>
<GID>2581</GID>
<name>IN_1</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>242.5,-2105.5,242.5,-2096.5</points>
<connection>
<GID>2583</GID>
<name>IN_1</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>296.5,-2104.5,296.5,-2096.5</points>
<intersection>-2104.5 118</intersection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>354.5,-2105,354.5,-2096.5</points>
<connection>
<GID>2587</GID>
<name>IN_1</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-19.5,-2098.5,-19.5,-2096.5</points>
<connection>
<GID>2572</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>30,-2098.5,30,-2096.5</points>
<connection>
<GID>2574</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>78,-2098.5,78,-2096.5</points>
<connection>
<GID>2576</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>127.5,-2098.5,127.5,-2096.5</points>
<connection>
<GID>2578</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>175.5,-2098.5,175.5,-2096.5</points>
<connection>
<GID>2580</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>233,-2098.5,233,-2096.5</points>
<connection>
<GID>2582</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>288,-2098.5,288,-2096.5</points>
<connection>
<GID>2584</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>345,-2098.5,345,-2096.5</points>
<connection>
<GID>2586</GID>
<name>clock</name></connection>
<intersection>-2096.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>135.5,-2104,136,-2104</points>
<connection>
<GID>2579</GID>
<name>IN_1</name></connection>
<intersection>135.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>296,-2104.5,296.5,-2104.5</points>
<connection>
<GID>2585</GID>
<name>IN_1</name></connection>
<intersection>296.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>1529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-2102,85.5,-2095.5</points>
<connection>
<GID>2577</GID>
<name>IN_0</name></connection>
<intersection>-2095.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84,-2095.5,85.5,-2095.5</points>
<connection>
<GID>2576</GID>
<name>OUT_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-2102,135,-2095.5</points>
<intersection>-2102 1</intersection>
<intersection>-2095.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-2102,136,-2102</points>
<connection>
<GID>2579</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133.5,-2095.5,135,-2095.5</points>
<connection>
<GID>2578</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>1531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-2101.5,183.5,-2095.5</points>
<intersection>-2101.5 5</intersection>
<intersection>-2095.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>181.5,-2095.5,183.5,-2095.5</points>
<connection>
<GID>2580</GID>
<name>OUT_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>183.5,-2101.5,184,-2101.5</points>
<connection>
<GID>2581</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-2103.5,242,-2095.5</points>
<intersection>-2103.5 1</intersection>
<intersection>-2095.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,-2103.5,242.5,-2103.5</points>
<connection>
<GID>2583</GID>
<name>IN_0</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>239,-2095.5,242,-2095.5</points>
<connection>
<GID>2582</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>1533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-2102.5,295.5,-2095.5</points>
<intersection>-2102.5 4</intersection>
<intersection>-2095.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>294,-2095.5,295.5,-2095.5</points>
<connection>
<GID>2584</GID>
<name>OUT_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>295.5,-2102.5,296,-2102.5</points>
<connection>
<GID>2585</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-2103,354,-2095.5</points>
<intersection>-2103 1</intersection>
<intersection>-2095.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-2103,354.5,-2103</points>
<connection>
<GID>2587</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-2095.5,354,-2095.5</points>
<connection>
<GID>2586</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment></shape></wire>
<wire>
<ID>1535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-2119.5,-12.5,-2113</points>
<intersection>-2119.5 1</intersection>
<intersection>-2113 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-2119.5,-10,-2119.5</points>
<connection>
<GID>2590</GID>
<name>IN_0</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-14,-2113,-12.5,-2113</points>
<connection>
<GID>2589</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-2120.5,36.5,-2113</points>
<intersection>-2120.5 1</intersection>
<intersection>-2113 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-2120.5,38.5,-2120.5</points>
<connection>
<GID>2592</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35.5,-2113,36.5,-2113</points>
<connection>
<GID>2591</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45.5,-2114,354,-2114</points>
<connection>
<GID>2605</GID>
<name>OUT</name></connection>
<intersection>-20 107</intersection>
<intersection>-11.5 4</intersection>
<intersection>29.5 108</intersection>
<intersection>37 16</intersection>
<intersection>77.5 109</intersection>
<intersection>84.5 23</intersection>
<intersection>127 110</intersection>
<intersection>135 31</intersection>
<intersection>175 111</intersection>
<intersection>183.5 55</intersection>
<intersection>232.5 112</intersection>
<intersection>242 56</intersection>
<intersection>287.5 113</intersection>
<intersection>296 66</intersection>
<intersection>344.5 114</intersection>
<intersection>354 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11.5,-2121.5,-11.5,-2114</points>
<intersection>-2121.5 5</intersection>
<intersection>-2114 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-11.5,-2121.5,-10,-2121.5</points>
<connection>
<GID>2590</GID>
<name>IN_1</name></connection>
<intersection>-11.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>37,-2122.5,37,-2114</points>
<intersection>-2122.5 21</intersection>
<intersection>-2114 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>37,-2122.5,38.5,-2122.5</points>
<connection>
<GID>2592</GID>
<name>IN_1</name></connection>
<intersection>37 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>84.5,-2121.5,84.5,-2114</points>
<intersection>-2121.5 53</intersection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>135,-2121.5,135,-2114</points>
<intersection>-2121.5 115</intersection>
<intersection>-2114 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>84.5,-2121.5,85,-2121.5</points>
<connection>
<GID>2594</GID>
<name>IN_1</name></connection>
<intersection>84.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>183.5,-2121,183.5,-2114</points>
<connection>
<GID>2598</GID>
<name>IN_1</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>242,-2123,242,-2114</points>
<connection>
<GID>2600</GID>
<name>IN_1</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>296,-2122,296,-2114</points>
<intersection>-2122 118</intersection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>354,-2122.5,354,-2114</points>
<connection>
<GID>2604</GID>
<name>IN_1</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-20,-2116,-20,-2114</points>
<connection>
<GID>2589</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>29.5,-2116,29.5,-2114</points>
<connection>
<GID>2591</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>77.5,-2116,77.5,-2114</points>
<connection>
<GID>2593</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>127,-2116,127,-2114</points>
<connection>
<GID>2595</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>175,-2116,175,-2114</points>
<connection>
<GID>2597</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>232.5,-2116,232.5,-2114</points>
<connection>
<GID>2599</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>287.5,-2116,287.5,-2114</points>
<connection>
<GID>2601</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>344.5,-2116,344.5,-2114</points>
<connection>
<GID>2603</GID>
<name>clock</name></connection>
<intersection>-2114 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>135,-2121.5,135.5,-2121.5</points>
<connection>
<GID>2596</GID>
<name>IN_1</name></connection>
<intersection>135 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>295.5,-2122,296,-2122</points>
<connection>
<GID>2602</GID>
<name>IN_1</name></connection>
<intersection>296 66</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-261.415,807.218,962.585,202.218</PageViewport>
<gate>
<ID>1159</ID>
<type>AA_AND2</type>
<position>114.5,-17.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1161</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-11.5</position>
<output>
<ID>OUT_0</ID>682 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1162</ID>
<type>AA_AND2</type>
<position>173,-18</position>
<input>
<ID>IN_0</ID>682 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>-232.5,26.5</position>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1163</ID>
<type>AA_AND2</type>
<position>-232.5,-10.5</position>
<output>
<ID>OUT</ID>676 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_DFF_LOW</type>
<position>-201,25.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1164</ID>
<type>AE_DFF_LOW</type>
<position>-201,-29</position>
<output>
<ID>OUT_0</ID>683 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>-191,20</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1165</ID>
<type>AA_AND2</type>
<position>-191,-34.5</position>
<input>
<ID>IN_0</ID>683 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,25.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1166</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,-29</position>
<output>
<ID>OUT_0</ID>684 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1167</ID>
<type>AA_AND2</type>
<position>-142.5,-35.5</position>
<input>
<ID>IN_0</ID>684 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>-142.5,19</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1168</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,-29</position>
<output>
<ID>OUT_0</ID>686 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,25.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1169</ID>
<type>AA_AND2</type>
<position>-96,-34.5</position>
<input>
<ID>IN_0</ID>686 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>-96,20</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1170</ID>
<type>AE_DFF_LOW</type>
<position>-54,-29</position>
<output>
<ID>OUT_0</ID>687 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_DFF_LOW</type>
<position>-54,25.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1171</ID>
<type>AA_AND2</type>
<position>-45.5,-34.5</position>
<input>
<ID>IN_0</ID>687 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>-46.5,20.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1172</ID>
<type>AE_DFF_LOW</type>
<position>-6,-29</position>
<output>
<ID>OUT_0</ID>688 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_DFF_LOW</type>
<position>-6,25.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1173</ID>
<type>AA_AND2</type>
<position>2.5,-34</position>
<input>
<ID>IN_0</ID>688 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>2.5,20.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1174</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-29</position>
<output>
<ID>OUT_0</ID>689 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_DFF_LOW</type>
<position>51.5,25.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1175</ID>
<type>AA_AND2</type>
<position>61,-36</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>61,18.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1176</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-29</position>
<output>
<ID>OUT_0</ID>690 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_DFF_LOW</type>
<position>106.5,25.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1177</ID>
<type>AA_AND2</type>
<position>114.5,-35</position>
<input>
<ID>IN_0</ID>690 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND2</type>
<position>113,19</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1178</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-29</position>
<output>
<ID>OUT_0</ID>691 </output>
<input>
<ID>clock</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_DFF_LOW</type>
<position>163.5,25.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1179</ID>
<type>AA_AND2</type>
<position>173,-35.5</position>
<input>
<ID>IN_0</ID>691 </input>
<input>
<ID>IN_1</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>173,19</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1180</ID>
<type>AA_AND2</type>
<position>-232.5,-28</position>
<output>
<ID>OUT</ID>685 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_DFF_LOW</type>
<position>-201,7.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1181</ID>
<type>AE_DFF_LOW</type>
<position>-201,-45</position>
<output>
<ID>OUT_0</ID>692 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>-191,2</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1182</ID>
<type>AA_AND2</type>
<position>-191,-50.5</position>
<input>
<ID>IN_0</ID>692 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,7.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1183</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,-45</position>
<output>
<ID>OUT_0</ID>693 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>-142.5,1</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1184</ID>
<type>AA_AND2</type>
<position>-142.5,-51.5</position>
<input>
<ID>IN_0</ID>693 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,7.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1185</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,-45</position>
<output>
<ID>OUT_0</ID>695 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW_NT</type>
<position>58.5,-26.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUTINV_0</ID>21 </output>
<output>
<ID>OUT_0</ID>11 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1186</ID>
<type>AA_AND2</type>
<position>-96,-50.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>40,-35</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1187</ID>
<type>AE_DFF_LOW</type>
<position>-54,-45</position>
<output>
<ID>OUT_0</ID>696 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND3</type>
<position>67,-37.5</position>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>11 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1188</ID>
<type>AA_AND2</type>
<position>-45.5,-50.5</position>
<input>
<ID>IN_0</ID>696 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>31.5,-24</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1189</ID>
<type>AE_DFF_LOW</type>
<position>-6,-45</position>
<output>
<ID>OUT_0</ID>697 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>23.5,-36</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1190</ID>
<type>AA_AND2</type>
<position>2.5,-50</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>-96,2</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1191</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-45</position>
<output>
<ID>OUT_0</ID>698 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>-54,7.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1192</ID>
<type>AA_AND2</type>
<position>61,-52</position>
<input>
<ID>IN_0</ID>698 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>67,-44.5</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1193</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-45</position>
<output>
<ID>OUT_0</ID>699 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>-45.5,2</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1194</ID>
<type>AA_AND2</type>
<position>114.5,-51</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>21,-29.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1195</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-45</position>
<output>
<ID>OUT_0</ID>700 </output>
<input>
<ID>clock</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_DFF_LOW</type>
<position>-6,7.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1196</ID>
<type>AA_AND2</type>
<position>173,-51.5</position>
<input>
<ID>IN_0</ID>700 </input>
<input>
<ID>IN_1</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>2.5,2.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1197</ID>
<type>AA_AND2</type>
<position>-232.5,-44</position>
<output>
<ID>OUT</ID>694 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>51.5,7.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1198</ID>
<type>AE_DFF_LOW</type>
<position>-201,-61.5</position>
<output>
<ID>OUT_0</ID>701 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>61,0.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1199</ID>
<type>AA_AND2</type>
<position>-191,-67</position>
<input>
<ID>IN_0</ID>701 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_DFF_LOW</type>
<position>106.5,7.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1200</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,-61.5</position>
<output>
<ID>OUT_0</ID>702 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1201</ID>
<type>AA_AND2</type>
<position>-142.5,-68</position>
<input>
<ID>IN_0</ID>702 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>114.5,1.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1202</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,-61.5</position>
<output>
<ID>OUT_0</ID>704 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1203</ID>
<type>AA_AND2</type>
<position>-96,-67</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>163.5,7.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1204</ID>
<type>AE_DFF_LOW</type>
<position>-54,-61.5</position>
<output>
<ID>OUT_0</ID>705 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>173,1</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1205</ID>
<type>AA_AND2</type>
<position>-45.5,-67</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>-232.5,8.5</position>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1206</ID>
<type>AE_DFF_LOW</type>
<position>-6,-61.5</position>
<output>
<ID>OUT_0</ID>706 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW</type>
<position>-201,-11.5</position>
<output>
<ID>OUT_0</ID>672 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1207</ID>
<type>AA_AND2</type>
<position>2.5,-66.5</position>
<input>
<ID>IN_0</ID>706 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>-191,-17</position>
<input>
<ID>IN_0</ID>672 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1208</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-61.5</position>
<output>
<ID>OUT_0</ID>707 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1209</ID>
<type>AA_AND2</type>
<position>61,-68.5</position>
<input>
<ID>IN_0</ID>707 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1210</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-61.5</position>
<output>
<ID>OUT_0</ID>708 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,-11.5</position>
<output>
<ID>OUT_0</ID>675 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1211</ID>
<type>AA_AND2</type>
<position>114.5,-67.5</position>
<input>
<ID>IN_0</ID>708 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>-142.5,-18</position>
<input>
<ID>IN_0</ID>675 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1212</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-61.5</position>
<output>
<ID>OUT_0</ID>709 </output>
<input>
<ID>clock</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,-11.5</position>
<output>
<ID>OUT_0</ID>677 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1213</ID>
<type>AA_AND2</type>
<position>173,-68</position>
<input>
<ID>IN_0</ID>709 </input>
<input>
<ID>IN_1</ID>703 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>-96,-17</position>
<input>
<ID>IN_0</ID>677 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1214</ID>
<type>AA_AND2</type>
<position>-232.5,-60.5</position>
<output>
<ID>OUT</ID>703 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_DFF_LOW</type>
<position>-54,-11.5</position>
<output>
<ID>OUT_0</ID>678 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1215</ID>
<type>AE_DFF_LOW</type>
<position>-201,-79.5</position>
<output>
<ID>OUT_0</ID>710 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1216</ID>
<type>AA_AND2</type>
<position>-191,-85</position>
<input>
<ID>IN_0</ID>710 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1217</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,-79.5</position>
<output>
<ID>OUT_0</ID>711 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1218</ID>
<type>AA_AND2</type>
<position>-142.5,-86</position>
<input>
<ID>IN_0</ID>711 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1219</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,-79.5</position>
<output>
<ID>OUT_0</ID>713 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1220</ID>
<type>AA_AND2</type>
<position>-96,-85</position>
<input>
<ID>IN_0</ID>713 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1221</ID>
<type>AE_DFF_LOW</type>
<position>-54,-79.5</position>
<output>
<ID>OUT_0</ID>714 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1222</ID>
<type>AA_AND2</type>
<position>-45.5,-85</position>
<input>
<ID>IN_0</ID>714 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1223</ID>
<type>AE_DFF_LOW</type>
<position>-6,-79.5</position>
<output>
<ID>OUT_0</ID>715 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1224</ID>
<type>AA_AND2</type>
<position>2.5,-84.5</position>
<input>
<ID>IN_0</ID>715 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1225</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-79.5</position>
<output>
<ID>OUT_0</ID>716 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1226</ID>
<type>AA_AND2</type>
<position>61,-86.5</position>
<input>
<ID>IN_0</ID>716 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1227</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-79.5</position>
<output>
<ID>OUT_0</ID>717 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1228</ID>
<type>AA_AND2</type>
<position>114.5,-85.5</position>
<input>
<ID>IN_0</ID>717 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1229</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-79.5</position>
<output>
<ID>OUT_0</ID>718 </output>
<input>
<ID>clock</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1230</ID>
<type>AA_AND2</type>
<position>173,-86</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1231</ID>
<type>AA_AND2</type>
<position>-232.5,-78.5</position>
<output>
<ID>OUT</ID>712 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1232</ID>
<type>AE_DFF_LOW</type>
<position>-201,-101.5</position>
<output>
<ID>OUT_0</ID>719 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1233</ID>
<type>AA_AND2</type>
<position>-191,-107</position>
<input>
<ID>IN_0</ID>719 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1234</ID>
<type>AE_DFF_LOW</type>
<position>-151.5,-101.5</position>
<output>
<ID>OUT_0</ID>720 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1235</ID>
<type>AA_AND2</type>
<position>-142.5,-108</position>
<input>
<ID>IN_0</ID>720 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1236</ID>
<type>AE_DFF_LOW</type>
<position>-103.5,-101.5</position>
<output>
<ID>OUT_0</ID>722 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1237</ID>
<type>AA_AND2</type>
<position>-96,-107</position>
<input>
<ID>IN_0</ID>722 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1238</ID>
<type>AE_DFF_LOW</type>
<position>-54,-101.5</position>
<output>
<ID>OUT_0</ID>723 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1239</ID>
<type>AA_AND2</type>
<position>-45.5,-107</position>
<input>
<ID>IN_0</ID>723 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1240</ID>
<type>AE_DFF_LOW</type>
<position>-6,-101.5</position>
<output>
<ID>OUT_0</ID>724 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1241</ID>
<type>AA_AND2</type>
<position>2.5,-106.5</position>
<input>
<ID>IN_0</ID>724 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1242</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-101.5</position>
<output>
<ID>OUT_0</ID>725 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1243</ID>
<type>AA_AND2</type>
<position>61,-108.5</position>
<input>
<ID>IN_0</ID>725 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1244</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-101.5</position>
<output>
<ID>OUT_0</ID>726 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>-45.5,-17</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1245</ID>
<type>AA_AND2</type>
<position>114.5,-107.5</position>
<input>
<ID>IN_0</ID>726 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1246</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-101.5</position>
<output>
<ID>OUT_0</ID>727 </output>
<input>
<ID>clock</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1247</ID>
<type>AA_AND2</type>
<position>173,-108</position>
<input>
<ID>IN_0</ID>727 </input>
<input>
<ID>IN_1</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1248</ID>
<type>AA_AND2</type>
<position>-232.5,-100.5</position>
<output>
<ID>OUT</ID>721 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1149</ID>
<type>AE_DFF_LOW</type>
<position>-6,-11.5</position>
<output>
<ID>OUT_0</ID>679 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1150</ID>
<type>AA_AND2</type>
<position>2.5,-16.5</position>
<input>
<ID>IN_0</ID>679 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1151</ID>
<type>AE_DFF_LOW</type>
<position>51.5,-11.5</position>
<output>
<ID>OUT_0</ID>680 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1155</ID>
<type>AA_AND2</type>
<position>61,-18.5</position>
<input>
<ID>IN_0</ID>680 </input>
<input>
<ID>IN_1</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1157</ID>
<type>AE_DFF_LOW</type>
<position>106.5,-11.5</position>
<output>
<ID>OUT_0</ID>681 </output>
<input>
<ID>clock</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,21,-196.5,27.5</points>
<intersection>21 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,21,-194,21</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-198,27.5,-196.5,27.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,20,-147.5,27.5</points>
<intersection>20 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,20,-145.5,20</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-148.5,27.5,-147.5,27.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,26.5,170,26.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-204 82</intersection>
<intersection>-196 4</intersection>
<intersection>-154.5 80</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 81</intersection>
<intersection>-98.5 23</intersection>
<intersection>-57 79</intersection>
<intersection>-49.5 31</intersection>
<intersection>-9 83</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 84</intersection>
<intersection>58 56</intersection>
<intersection>103.5 78</intersection>
<intersection>110 66</intersection>
<intersection>160.5 85</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-196,19,-196,26.5</points>
<intersection>19 5</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-196,19,-194,19</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-196 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,18,-147,26.5</points>
<intersection>18 21</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,18,-145.5,18</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-98.5,19,-98.5,26.5</points>
<intersection>19 53</intersection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49.5,19.5,-49.5,26.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99,19,-98.5,19</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-98.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,19.5,-0.5,26.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,17.5,58,26.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>110,18,110,26.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,18,170,26.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>103.5,24.5,103.5,26.5</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>79</ID>
<points>-57,24.5,-57,26.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>80</ID>
<points>-154.5,24.5,-154.5,26.5</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>81</ID>
<points>-106.5,24.5,-106.5,26.5</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>82</ID>
<points>-204,24.5,-204,26.5</points>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>83</ID>
<points>-9,24.5,-9,26.5</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>84</ID>
<points>48.5,24.5,48.5,26.5</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment>
<vsegment>
<ID>85</ID>
<points>160.5,24.5,160.5,26.5</points>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<intersection>26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,21,-99,27.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-100.5,27.5,-99,27.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,21.5,-50,27.5</points>
<intersection>21.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,21.5,-49.5,21.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-51,27.5,-50,27.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-50 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-34.5,65,-24.5</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-24.5,65,-24.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,21.5,-1,27.5</points>
<intersection>21.5 5</intersection>
<intersection>27.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,27.5,-1,27.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,21.5,-0.5,21.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-36,37,-36</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,19.5,57.5,27.5</points>
<intersection>19.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,19.5,58,19.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,27.5,57.5,27.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,20,109.5,27.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,20,110,20</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-43.5,67,-40.5</points>
<connection>
<GID>34</GID>
<name>N_in3</name></connection>
<connection>
<GID>29</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-24,55.5,-24</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>55.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55.5,-24.5,55.5,-24</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-34,30,-29.5</points>
<intersection>-34 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-34,37,-34</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-29.5,30,-29.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,20,169.5,27.5</points>
<intersection>20 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,20,170,20</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,27.5,169.5,27.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-35,49,-27.5</points>
<intersection>-35 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-27.5,55.5,-27.5</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-35,49,-35</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-34.5,67,-27.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-27.5,67,-27.5</points>
<connection>
<GID>27</GID>
<name>OUTINV_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,3,-196.5,9.5</points>
<intersection>3 1</intersection>
<intersection>9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,3,-194,3</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,9.5,-196.5,9.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,2,-147.5,9.5</points>
<intersection>2 1</intersection>
<intersection>9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,2,-145.5,2</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,9.5,-147.5,9.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,8.5,170,8.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,1,-195.5,8.5</points>
<intersection>1 5</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,1,-194,1</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,0,-147,8.5</points>
<intersection>0 21</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,0,-145.5,0</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,1,-99.5,8.5</points>
<intersection>1 53</intersection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,1,-49,8.5</points>
<intersection>1 115</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,1,-99,1</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,1.5,-0.5,8.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-0.5,58,8.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,0.5,112,8.5</points>
<intersection>0.5 118</intersection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,0,170,8.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,6.5,-204,8.5</points>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,6.5,-154.5,8.5</points>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,6.5,-106.5,8.5</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,6.5,-57,8.5</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,6.5,-9,8.5</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,6.5,48.5,8.5</points>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,6.5,103.5,8.5</points>
<connection>
<GID>41</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,6.5,160.5,8.5</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,1,-48.5,1</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,0.5,112,0.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,3,-99,9.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,9.5,-99,9.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,3,-49.5,9.5</points>
<intersection>3 1</intersection>
<intersection>9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,3,-48.5,3</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,9.5,-49.5,9.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,3.5,-1,9.5</points>
<intersection>3.5 5</intersection>
<intersection>9.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,9.5,-1,9.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,3.5,-0.5,3.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,1.5,57.5,9.5</points>
<intersection>1.5 1</intersection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,1.5,58,1.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,9.5,57.5,9.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,2.5,111,9.5</points>
<intersection>2.5 4</intersection>
<intersection>9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,9.5,111,9.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,2.5,111.5,2.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,2,169.5,9.5</points>
<intersection>2 1</intersection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,2,170,2</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,9.5,169.5,9.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,-16,-196.5,-9.5</points>
<intersection>-16 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,-16,-194,-16</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,-9.5,-196.5,-9.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,-17,-147.5,-9.5</points>
<intersection>-17 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,-17,-145.5,-17</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-9.5,-147.5,-9.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,-10.5,170,-10.5</points>
<connection>
<GID>1163</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-18,-195.5,-10.5</points>
<intersection>-18 5</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,-18,-194,-18</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,-19,-147,-10.5</points>
<intersection>-19 21</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,-19,-145.5,-19</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,-18,-99.5,-10.5</points>
<intersection>-18 53</intersection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,-18,-49,-10.5</points>
<intersection>-18 115</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,-18,-99,-18</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,-17.5,-0.5,-10.5</points>
<connection>
<GID>1150</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-19.5,58,-10.5</points>
<connection>
<GID>1155</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,-18.5,112,-10.5</points>
<intersection>-18.5 118</intersection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,-19,170,-10.5</points>
<connection>
<GID>1162</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,-12.5,-204,-10.5</points>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,-12.5,-154.5,-10.5</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,-12.5,-106.5,-10.5</points>
<connection>
<GID>54</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,-12.5,-57,-10.5</points>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,-12.5,-9,-10.5</points>
<connection>
<GID>1149</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,-12.5,48.5,-10.5</points>
<connection>
<GID>1151</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,-12.5,103.5,-10.5</points>
<connection>
<GID>1157</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,-12.5,160.5,-10.5</points>
<connection>
<GID>1161</GID>
<name>clock</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,-18,-48.5,-18</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,-18.5,112,-18.5</points>
<connection>
<GID>1159</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,-16,-99,-9.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,-9.5,-99,-9.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,-16,-49.5,-9.5</points>
<intersection>-16 1</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-16,-48.5,-16</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,-9.5,-49.5,-9.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-15.5,-1,-9.5</points>
<intersection>-15.5 5</intersection>
<intersection>-9.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,-9.5,-1,-9.5</points>
<connection>
<GID>1149</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,-15.5,-0.5,-15.5</points>
<connection>
<GID>1150</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-17.5,57.5,-9.5</points>
<intersection>-17.5 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-17.5,58,-17.5</points>
<connection>
<GID>1155</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-9.5,57.5,-9.5</points>
<connection>
<GID>1151</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-16.5,111,-9.5</points>
<intersection>-16.5 4</intersection>
<intersection>-9.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-9.5,111,-9.5</points>
<connection>
<GID>1157</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-16.5,111.5,-16.5</points>
<connection>
<GID>1159</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-17,169.5,-9.5</points>
<intersection>-17 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-17,170,-17</points>
<connection>
<GID>1162</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-9.5,169.5,-9.5</points>
<connection>
<GID>1161</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,-33.5,-196.5,-27</points>
<intersection>-33.5 1</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,-33.5,-194,-33.5</points>
<connection>
<GID>1165</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,-27,-196.5,-27</points>
<connection>
<GID>1164</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,-34.5,-147.5,-27</points>
<intersection>-34.5 1</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,-34.5,-145.5,-34.5</points>
<connection>
<GID>1167</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-27,-147.5,-27</points>
<connection>
<GID>1166</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,-28,170,-28</points>
<connection>
<GID>1180</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-35.5,-195.5,-28</points>
<intersection>-35.5 5</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,-35.5,-194,-35.5</points>
<connection>
<GID>1165</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,-36.5,-147,-28</points>
<intersection>-36.5 21</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,-36.5,-145.5,-36.5</points>
<connection>
<GID>1167</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,-35.5,-99.5,-28</points>
<intersection>-35.5 53</intersection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,-35.5,-49,-28</points>
<intersection>-35.5 115</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,-35.5,-99,-35.5</points>
<connection>
<GID>1169</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,-35,-0.5,-28</points>
<connection>
<GID>1173</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-37,58,-28</points>
<connection>
<GID>1175</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,-36,112,-28</points>
<intersection>-36 118</intersection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,-36.5,170,-28</points>
<connection>
<GID>1179</GID>
<name>IN_1</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,-30,-204,-28</points>
<connection>
<GID>1164</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,-30,-154.5,-28</points>
<connection>
<GID>1166</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,-30,-106.5,-28</points>
<connection>
<GID>1168</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,-30,-57,-28</points>
<connection>
<GID>1170</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,-30,-9,-28</points>
<connection>
<GID>1172</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,-30,48.5,-28</points>
<connection>
<GID>1174</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,-30,103.5,-28</points>
<connection>
<GID>1176</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,-30,160.5,-28</points>
<connection>
<GID>1178</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,-35.5,-48.5,-35.5</points>
<connection>
<GID>1171</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,-36,112,-36</points>
<connection>
<GID>1177</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,-33.5,-99,-27</points>
<connection>
<GID>1169</GID>
<name>IN_0</name></connection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,-27,-99,-27</points>
<connection>
<GID>1168</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,-33.5,-49.5,-27</points>
<intersection>-33.5 1</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-33.5,-48.5,-33.5</points>
<connection>
<GID>1171</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,-27,-49.5,-27</points>
<connection>
<GID>1170</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-33,-1,-27</points>
<intersection>-33 5</intersection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,-27,-1,-27</points>
<connection>
<GID>1172</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,-33,-0.5,-33</points>
<connection>
<GID>1173</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-35,57.5,-27</points>
<intersection>-35 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-35,58,-35</points>
<connection>
<GID>1175</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-27,57.5,-27</points>
<connection>
<GID>1174</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-34,111,-27</points>
<intersection>-34 4</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-27,111,-27</points>
<connection>
<GID>1176</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-34,111.5,-34</points>
<connection>
<GID>1177</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-34.5,169.5,-27</points>
<intersection>-34.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-34.5,170,-34.5</points>
<connection>
<GID>1179</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-27,169.5,-27</points>
<connection>
<GID>1178</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,-49.5,-196.5,-43</points>
<intersection>-49.5 1</intersection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,-49.5,-194,-49.5</points>
<connection>
<GID>1182</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,-43,-196.5,-43</points>
<connection>
<GID>1181</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,-50.5,-147.5,-43</points>
<intersection>-50.5 1</intersection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,-50.5,-145.5,-50.5</points>
<connection>
<GID>1184</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-43,-147.5,-43</points>
<connection>
<GID>1183</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,-44,170,-44</points>
<connection>
<GID>1197</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-51.5,-195.5,-44</points>
<intersection>-51.5 5</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,-51.5,-194,-51.5</points>
<connection>
<GID>1182</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,-52.5,-147,-44</points>
<intersection>-52.5 21</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,-52.5,-145.5,-52.5</points>
<connection>
<GID>1184</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,-51.5,-99.5,-44</points>
<intersection>-51.5 53</intersection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,-51.5,-49,-44</points>
<intersection>-51.5 115</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,-51.5,-99,-51.5</points>
<connection>
<GID>1186</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,-51,-0.5,-44</points>
<connection>
<GID>1190</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-53,58,-44</points>
<connection>
<GID>1192</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,-52,112,-44</points>
<intersection>-52 118</intersection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,-52.5,170,-44</points>
<connection>
<GID>1196</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,-46,-204,-44</points>
<connection>
<GID>1181</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,-46,-154.5,-44</points>
<connection>
<GID>1183</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,-46,-106.5,-44</points>
<connection>
<GID>1185</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,-46,-57,-44</points>
<connection>
<GID>1187</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,-46,-9,-44</points>
<connection>
<GID>1189</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,-46,48.5,-44</points>
<connection>
<GID>1191</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,-46,103.5,-44</points>
<connection>
<GID>1193</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,-46,160.5,-44</points>
<connection>
<GID>1195</GID>
<name>clock</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,-51.5,-48.5,-51.5</points>
<connection>
<GID>1188</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,-52,112,-52</points>
<connection>
<GID>1194</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,-49.5,-99,-43</points>
<connection>
<GID>1186</GID>
<name>IN_0</name></connection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,-43,-99,-43</points>
<connection>
<GID>1185</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,-49.5,-49.5,-43</points>
<intersection>-49.5 1</intersection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-49.5,-48.5,-49.5</points>
<connection>
<GID>1188</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,-43,-49.5,-43</points>
<connection>
<GID>1187</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-49,-1,-43</points>
<intersection>-49 5</intersection>
<intersection>-43 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,-43,-1,-43</points>
<connection>
<GID>1189</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,-49,-0.5,-49</points>
<connection>
<GID>1190</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-51,57.5,-43</points>
<intersection>-51 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-51,58,-51</points>
<connection>
<GID>1192</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-43,57.5,-43</points>
<connection>
<GID>1191</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-50,111,-43</points>
<intersection>-50 4</intersection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-43,111,-43</points>
<connection>
<GID>1193</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-50,111.5,-50</points>
<connection>
<GID>1194</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-50.5,169.5,-43</points>
<intersection>-50.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-50.5,170,-50.5</points>
<connection>
<GID>1196</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-43,169.5,-43</points>
<connection>
<GID>1195</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,-66,-196.5,-59.5</points>
<intersection>-66 1</intersection>
<intersection>-59.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,-66,-194,-66</points>
<connection>
<GID>1199</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,-59.5,-196.5,-59.5</points>
<connection>
<GID>1198</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,-67,-147.5,-59.5</points>
<intersection>-67 1</intersection>
<intersection>-59.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,-67,-145.5,-67</points>
<connection>
<GID>1201</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-59.5,-147.5,-59.5</points>
<connection>
<GID>1200</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,-60.5,170,-60.5</points>
<connection>
<GID>1214</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-68,-195.5,-60.5</points>
<intersection>-68 5</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,-68,-194,-68</points>
<connection>
<GID>1199</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,-69,-147,-60.5</points>
<intersection>-69 21</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,-69,-145.5,-69</points>
<connection>
<GID>1201</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,-68,-99.5,-60.5</points>
<intersection>-68 53</intersection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,-68,-49,-60.5</points>
<intersection>-68 115</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,-68,-99,-68</points>
<connection>
<GID>1203</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,-67.5,-0.5,-60.5</points>
<connection>
<GID>1207</GID>
<name>IN_1</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-69.5,58,-60.5</points>
<connection>
<GID>1209</GID>
<name>IN_1</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,-68.5,112,-60.5</points>
<intersection>-68.5 118</intersection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,-69,170,-60.5</points>
<connection>
<GID>1213</GID>
<name>IN_1</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,-62.5,-204,-60.5</points>
<connection>
<GID>1198</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,-62.5,-154.5,-60.5</points>
<connection>
<GID>1200</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,-62.5,-106.5,-60.5</points>
<connection>
<GID>1202</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,-62.5,-57,-60.5</points>
<connection>
<GID>1204</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,-62.5,-9,-60.5</points>
<connection>
<GID>1206</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,-62.5,48.5,-60.5</points>
<connection>
<GID>1208</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,-62.5,103.5,-60.5</points>
<connection>
<GID>1210</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,-62.5,160.5,-60.5</points>
<connection>
<GID>1212</GID>
<name>clock</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,-68,-48.5,-68</points>
<connection>
<GID>1205</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,-68.5,112,-68.5</points>
<connection>
<GID>1211</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,-66,-99,-59.5</points>
<connection>
<GID>1203</GID>
<name>IN_0</name></connection>
<intersection>-59.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,-59.5,-99,-59.5</points>
<connection>
<GID>1202</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,-66,-49.5,-59.5</points>
<intersection>-66 1</intersection>
<intersection>-59.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-66,-48.5,-66</points>
<connection>
<GID>1205</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,-59.5,-49.5,-59.5</points>
<connection>
<GID>1204</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-65.5,-1,-59.5</points>
<intersection>-65.5 5</intersection>
<intersection>-59.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,-59.5,-1,-59.5</points>
<connection>
<GID>1206</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,-65.5,-0.5,-65.5</points>
<connection>
<GID>1207</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-67.5,57.5,-59.5</points>
<intersection>-67.5 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-67.5,58,-67.5</points>
<connection>
<GID>1209</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-59.5,57.5,-59.5</points>
<connection>
<GID>1208</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-66.5,111,-59.5</points>
<intersection>-66.5 4</intersection>
<intersection>-59.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-59.5,111,-59.5</points>
<connection>
<GID>1210</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-66.5,111.5,-66.5</points>
<connection>
<GID>1211</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-67,169.5,-59.5</points>
<intersection>-67 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-67,170,-67</points>
<connection>
<GID>1213</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-59.5,169.5,-59.5</points>
<connection>
<GID>1212</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,-84,-196.5,-77.5</points>
<intersection>-84 1</intersection>
<intersection>-77.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,-84,-194,-84</points>
<connection>
<GID>1216</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,-77.5,-196.5,-77.5</points>
<connection>
<GID>1215</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,-85,-147.5,-77.5</points>
<intersection>-85 1</intersection>
<intersection>-77.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,-85,-145.5,-85</points>
<connection>
<GID>1218</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-77.5,-147.5,-77.5</points>
<connection>
<GID>1217</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,-78.5,170,-78.5</points>
<connection>
<GID>1231</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-86,-195.5,-78.5</points>
<intersection>-86 5</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,-86,-194,-86</points>
<connection>
<GID>1216</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,-87,-147,-78.5</points>
<intersection>-87 21</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,-87,-145.5,-87</points>
<connection>
<GID>1218</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,-86,-99.5,-78.5</points>
<intersection>-86 53</intersection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,-86,-49,-78.5</points>
<intersection>-86 115</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,-86,-99,-86</points>
<connection>
<GID>1220</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,-85.5,-0.5,-78.5</points>
<connection>
<GID>1224</GID>
<name>IN_1</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-87.5,58,-78.5</points>
<connection>
<GID>1226</GID>
<name>IN_1</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,-86.5,112,-78.5</points>
<intersection>-86.5 118</intersection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,-87,170,-78.5</points>
<connection>
<GID>1230</GID>
<name>IN_1</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,-80.5,-204,-78.5</points>
<connection>
<GID>1215</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,-80.5,-154.5,-78.5</points>
<connection>
<GID>1217</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,-80.5,-106.5,-78.5</points>
<connection>
<GID>1219</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,-80.5,-57,-78.5</points>
<connection>
<GID>1221</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,-80.5,-9,-78.5</points>
<connection>
<GID>1223</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,-80.5,48.5,-78.5</points>
<connection>
<GID>1225</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,-80.5,103.5,-78.5</points>
<connection>
<GID>1227</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,-80.5,160.5,-78.5</points>
<connection>
<GID>1229</GID>
<name>clock</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,-86,-48.5,-86</points>
<connection>
<GID>1222</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,-86.5,112,-86.5</points>
<connection>
<GID>1228</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,-84,-99,-77.5</points>
<connection>
<GID>1220</GID>
<name>IN_0</name></connection>
<intersection>-77.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,-77.5,-99,-77.5</points>
<connection>
<GID>1219</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,-84,-49.5,-77.5</points>
<intersection>-84 1</intersection>
<intersection>-77.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-84,-48.5,-84</points>
<connection>
<GID>1222</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,-77.5,-49.5,-77.5</points>
<connection>
<GID>1221</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-83.5,-1,-77.5</points>
<intersection>-83.5 5</intersection>
<intersection>-77.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,-77.5,-1,-77.5</points>
<connection>
<GID>1223</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,-83.5,-0.5,-83.5</points>
<connection>
<GID>1224</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-85.5,57.5,-77.5</points>
<intersection>-85.5 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-85.5,58,-85.5</points>
<connection>
<GID>1226</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-77.5,57.5,-77.5</points>
<connection>
<GID>1225</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-84.5,111,-77.5</points>
<intersection>-84.5 4</intersection>
<intersection>-77.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-77.5,111,-77.5</points>
<connection>
<GID>1227</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-84.5,111.5,-84.5</points>
<connection>
<GID>1228</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-85,169.5,-77.5</points>
<intersection>-85 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-85,170,-85</points>
<connection>
<GID>1230</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-77.5,169.5,-77.5</points>
<connection>
<GID>1229</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196.5,-106,-196.5,-99.5</points>
<intersection>-106 1</intersection>
<intersection>-99.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196.5,-106,-194,-106</points>
<connection>
<GID>1233</GID>
<name>IN_0</name></connection>
<intersection>-196.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-198,-99.5,-196.5,-99.5</points>
<connection>
<GID>1232</GID>
<name>OUT_0</name></connection>
<intersection>-196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147.5,-107,-147.5,-99.5</points>
<intersection>-107 1</intersection>
<intersection>-99.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147.5,-107,-145.5,-107</points>
<connection>
<GID>1235</GID>
<name>IN_0</name></connection>
<intersection>-147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-99.5,-147.5,-99.5</points>
<connection>
<GID>1234</GID>
<name>OUT_0</name></connection>
<intersection>-147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-229.5,-100.5,170,-100.5</points>
<connection>
<GID>1248</GID>
<name>OUT</name></connection>
<intersection>-204 107</intersection>
<intersection>-195.5 4</intersection>
<intersection>-154.5 108</intersection>
<intersection>-147 16</intersection>
<intersection>-106.5 109</intersection>
<intersection>-99.5 23</intersection>
<intersection>-57 110</intersection>
<intersection>-49 31</intersection>
<intersection>-9 111</intersection>
<intersection>-0.5 55</intersection>
<intersection>48.5 112</intersection>
<intersection>58 56</intersection>
<intersection>103.5 113</intersection>
<intersection>112 66</intersection>
<intersection>160.5 114</intersection>
<intersection>170 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-108,-195.5,-100.5</points>
<intersection>-108 5</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-195.5,-108,-194,-108</points>
<connection>
<GID>1233</GID>
<name>IN_1</name></connection>
<intersection>-195.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-147,-109,-147,-100.5</points>
<intersection>-109 21</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-147,-109,-145.5,-109</points>
<connection>
<GID>1235</GID>
<name>IN_1</name></connection>
<intersection>-147 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-99.5,-108,-99.5,-100.5</points>
<intersection>-108 53</intersection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-49,-108,-49,-100.5</points>
<intersection>-108 115</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>-99.5,-108,-99,-108</points>
<connection>
<GID>1237</GID>
<name>IN_1</name></connection>
<intersection>-99.5 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>-0.5,-107.5,-0.5,-100.5</points>
<connection>
<GID>1241</GID>
<name>IN_1</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>58,-109.5,58,-100.5</points>
<connection>
<GID>1243</GID>
<name>IN_1</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>112,-108.5,112,-100.5</points>
<intersection>-108.5 118</intersection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>170,-109,170,-100.5</points>
<connection>
<GID>1247</GID>
<name>IN_1</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-204,-102.5,-204,-100.5</points>
<connection>
<GID>1232</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-154.5,-102.5,-154.5,-100.5</points>
<connection>
<GID>1234</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-106.5,-102.5,-106.5,-100.5</points>
<connection>
<GID>1236</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-57,-102.5,-57,-100.5</points>
<connection>
<GID>1238</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-9,-102.5,-9,-100.5</points>
<connection>
<GID>1240</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>48.5,-102.5,48.5,-100.5</points>
<connection>
<GID>1242</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>103.5,-102.5,103.5,-100.5</points>
<connection>
<GID>1244</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>160.5,-102.5,160.5,-100.5</points>
<connection>
<GID>1246</GID>
<name>clock</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>-49,-108,-48.5,-108</points>
<connection>
<GID>1239</GID>
<name>IN_1</name></connection>
<intersection>-49 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>111.5,-108.5,112,-108.5</points>
<connection>
<GID>1245</GID>
<name>IN_1</name></connection>
<intersection>112 66</intersection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99,-106,-99,-99.5</points>
<connection>
<GID>1237</GID>
<name>IN_0</name></connection>
<intersection>-99.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100.5,-99.5,-99,-99.5</points>
<connection>
<GID>1236</GID>
<name>OUT_0</name></connection>
<intersection>-99 0</intersection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49.5,-106,-49.5,-99.5</points>
<intersection>-106 1</intersection>
<intersection>-99.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-106,-48.5,-106</points>
<connection>
<GID>1239</GID>
<name>IN_0</name></connection>
<intersection>-49.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-51,-99.5,-49.5,-99.5</points>
<connection>
<GID>1238</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-105.5,-1,-99.5</points>
<intersection>-105.5 5</intersection>
<intersection>-99.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-3,-99.5,-1,-99.5</points>
<connection>
<GID>1240</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1,-105.5,-0.5,-105.5</points>
<connection>
<GID>1241</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-107.5,57.5,-99.5</points>
<intersection>-107.5 1</intersection>
<intersection>-99.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-107.5,58,-107.5</points>
<connection>
<GID>1243</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-99.5,57.5,-99.5</points>
<connection>
<GID>1242</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-106.5,111,-99.5</points>
<intersection>-106.5 4</intersection>
<intersection>-99.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-99.5,111,-99.5</points>
<connection>
<GID>1244</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-106.5,111.5,-106.5</points>
<connection>
<GID>1245</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-107,169.5,-99.5</points>
<intersection>-107 1</intersection>
<intersection>-99.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-107,170,-107</points>
<connection>
<GID>1247</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,-99.5,169.5,-99.5</points>
<connection>
<GID>1246</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-307.385,556.518,916.615,-48.4823</PageViewport>
<gate>
<ID>1351</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-79</position>
<output>
<ID>OUT_0</ID>782 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1352</ID>
<type>AA_AND2</type>
<position>106.5,-84.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1353</ID>
<type>AE_DFF_LOW</type>
<position>146,-79</position>
<output>
<ID>OUT_0</ID>783 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1354</ID>
<type>AA_AND2</type>
<position>155,-85.5</position>
<input>
<ID>IN_0</ID>783 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1355</ID>
<type>AE_DFF_LOW</type>
<position>194,-79</position>
<output>
<ID>OUT_0</ID>785 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1356</ID>
<type>AA_AND2</type>
<position>201.5,-84.5</position>
<input>
<ID>IN_0</ID>785 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1357</ID>
<type>AE_DFF_LOW</type>
<position>243.5,-79</position>
<output>
<ID>OUT_0</ID>786 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1358</ID>
<type>AA_AND2</type>
<position>252,-84.5</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1359</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-79</position>
<output>
<ID>OUT_0</ID>787 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1360</ID>
<type>AA_AND2</type>
<position>300,-84</position>
<input>
<ID>IN_0</ID>787 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1361</ID>
<type>AE_DFF_LOW</type>
<position>349,-79</position>
<output>
<ID>OUT_0</ID>788 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1362</ID>
<type>AA_AND2</type>
<position>358.5,-86</position>
<input>
<ID>IN_0</ID>788 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1363</ID>
<type>AE_DFF_LOW</type>
<position>404,-79</position>
<output>
<ID>OUT_0</ID>789 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1364</ID>
<type>AA_AND2</type>
<position>412,-85</position>
<input>
<ID>IN_0</ID>789 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1365</ID>
<type>AE_DFF_LOW</type>
<position>461,-79</position>
<output>
<ID>OUT_0</ID>790 </output>
<input>
<ID>clock</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1366</ID>
<type>AA_AND2</type>
<position>470.5,-85.5</position>
<input>
<ID>IN_0</ID>790 </input>
<input>
<ID>IN_1</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1367</ID>
<type>AA_AND2</type>
<position>65,-78</position>
<output>
<ID>OUT</ID>784 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1368</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-101</position>
<output>
<ID>OUT_0</ID>791 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1369</ID>
<type>AA_AND2</type>
<position>106.5,-106.5</position>
<input>
<ID>IN_0</ID>791 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1370</ID>
<type>AE_DFF_LOW</type>
<position>146,-101</position>
<output>
<ID>OUT_0</ID>792 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1371</ID>
<type>AA_AND2</type>
<position>155,-107.5</position>
<input>
<ID>IN_0</ID>792 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1372</ID>
<type>AE_DFF_LOW</type>
<position>194,-101</position>
<output>
<ID>OUT_0</ID>794 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1373</ID>
<type>AA_AND2</type>
<position>201.5,-106.5</position>
<input>
<ID>IN_0</ID>794 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1374</ID>
<type>AE_DFF_LOW</type>
<position>243.5,-101</position>
<output>
<ID>OUT_0</ID>795 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1375</ID>
<type>AA_AND2</type>
<position>252,-106.5</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1376</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-101</position>
<output>
<ID>OUT_0</ID>796 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1377</ID>
<type>AA_AND2</type>
<position>300,-106</position>
<input>
<ID>IN_0</ID>796 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1378</ID>
<type>AE_DFF_LOW</type>
<position>349,-101</position>
<output>
<ID>OUT_0</ID>797 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1379</ID>
<type>AA_AND2</type>
<position>358.5,-108</position>
<input>
<ID>IN_0</ID>797 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1380</ID>
<type>AE_DFF_LOW</type>
<position>404,-101</position>
<output>
<ID>OUT_0</ID>798 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1381</ID>
<type>AA_AND2</type>
<position>412,-107</position>
<input>
<ID>IN_0</ID>798 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1382</ID>
<type>AE_DFF_LOW</type>
<position>461,-101</position>
<output>
<ID>OUT_0</ID>799 </output>
<input>
<ID>clock</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1383</ID>
<type>AA_AND2</type>
<position>470.5,-107.5</position>
<input>
<ID>IN_0</ID>799 </input>
<input>
<ID>IN_1</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1384</ID>
<type>AA_AND2</type>
<position>65,-100</position>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1249</ID>
<type>AA_AND2</type>
<position>65,27</position>
<output>
<ID>OUT</ID>730 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1250</ID>
<type>AE_DFF_LOW</type>
<position>96.5,26</position>
<output>
<ID>OUT_0</ID>728 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1251</ID>
<type>AA_AND2</type>
<position>106.5,20.5</position>
<input>
<ID>IN_0</ID>728 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1252</ID>
<type>AE_DFF_LOW</type>
<position>146,26</position>
<output>
<ID>OUT_0</ID>729 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1253</ID>
<type>AA_AND2</type>
<position>155,19.5</position>
<input>
<ID>IN_0</ID>729 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1254</ID>
<type>AE_DFF_LOW</type>
<position>194,26</position>
<output>
<ID>OUT_0</ID>731 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1255</ID>
<type>AA_AND2</type>
<position>201.5,20.5</position>
<input>
<ID>IN_0</ID>731 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1256</ID>
<type>AE_DFF_LOW</type>
<position>243.5,26</position>
<output>
<ID>OUT_0</ID>732 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1257</ID>
<type>AA_AND2</type>
<position>251,21</position>
<input>
<ID>IN_0</ID>732 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1258</ID>
<type>AE_DFF_LOW</type>
<position>291.5,26</position>
<output>
<ID>OUT_0</ID>733 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1259</ID>
<type>AA_AND2</type>
<position>300,21</position>
<input>
<ID>IN_0</ID>733 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1260</ID>
<type>AE_DFF_LOW</type>
<position>349,26</position>
<output>
<ID>OUT_0</ID>734 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1261</ID>
<type>AA_AND2</type>
<position>358.5,19</position>
<input>
<ID>IN_0</ID>734 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1262</ID>
<type>AE_DFF_LOW</type>
<position>404,26</position>
<output>
<ID>OUT_0</ID>735 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1263</ID>
<type>AA_AND2</type>
<position>410.5,19.5</position>
<input>
<ID>IN_0</ID>735 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1264</ID>
<type>AE_DFF_LOW</type>
<position>461,26</position>
<output>
<ID>OUT_0</ID>736 </output>
<input>
<ID>clock</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1265</ID>
<type>AA_AND2</type>
<position>470.5,19.5</position>
<input>
<ID>IN_0</ID>736 </input>
<input>
<ID>IN_1</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1266</ID>
<type>AE_DFF_LOW</type>
<position>96.5,8</position>
<output>
<ID>OUT_0</ID>737 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1267</ID>
<type>AA_AND2</type>
<position>106.5,2.5</position>
<input>
<ID>IN_0</ID>737 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1268</ID>
<type>AE_DFF_LOW</type>
<position>146,8</position>
<output>
<ID>OUT_0</ID>738 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1269</ID>
<type>AA_AND2</type>
<position>155,1.5</position>
<input>
<ID>IN_0</ID>738 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1270</ID>
<type>AE_DFF_LOW</type>
<position>194,8</position>
<output>
<ID>OUT_0</ID>740 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1271</ID>
<type>AA_AND2</type>
<position>201.5,2.5</position>
<input>
<ID>IN_0</ID>740 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1272</ID>
<type>AE_DFF_LOW</type>
<position>243.5,8</position>
<output>
<ID>OUT_0</ID>741 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1273</ID>
<type>AA_AND2</type>
<position>252,2.5</position>
<input>
<ID>IN_0</ID>741 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1274</ID>
<type>AE_DFF_LOW</type>
<position>291.5,8</position>
<output>
<ID>OUT_0</ID>742 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1275</ID>
<type>AA_AND2</type>
<position>300,3</position>
<input>
<ID>IN_0</ID>742 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1276</ID>
<type>AE_DFF_LOW</type>
<position>349,8</position>
<output>
<ID>OUT_0</ID>743 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1277</ID>
<type>AA_AND2</type>
<position>358.5,1</position>
<input>
<ID>IN_0</ID>743 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1278</ID>
<type>AE_DFF_LOW</type>
<position>404,8</position>
<output>
<ID>OUT_0</ID>744 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1279</ID>
<type>AA_AND2</type>
<position>412,2</position>
<input>
<ID>IN_0</ID>744 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1280</ID>
<type>AE_DFF_LOW</type>
<position>461,8</position>
<output>
<ID>OUT_0</ID>745 </output>
<input>
<ID>clock</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1281</ID>
<type>AA_AND2</type>
<position>470.5,1.5</position>
<input>
<ID>IN_0</ID>745 </input>
<input>
<ID>IN_1</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1282</ID>
<type>AA_AND2</type>
<position>65,9</position>
<output>
<ID>OUT</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1283</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-11</position>
<output>
<ID>OUT_0</ID>746 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1284</ID>
<type>AA_AND2</type>
<position>106.5,-16.5</position>
<input>
<ID>IN_0</ID>746 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1285</ID>
<type>AE_DFF_LOW</type>
<position>146,-11</position>
<output>
<ID>OUT_0</ID>747 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1286</ID>
<type>AA_AND2</type>
<position>155,-17.5</position>
<input>
<ID>IN_0</ID>747 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1287</ID>
<type>AE_DFF_LOW</type>
<position>194,-11</position>
<output>
<ID>OUT_0</ID>749 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1288</ID>
<type>AA_AND2</type>
<position>201.5,-16.5</position>
<input>
<ID>IN_0</ID>749 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1289</ID>
<type>AE_DFF_LOW</type>
<position>243.5,-11</position>
<output>
<ID>OUT_0</ID>750 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1290</ID>
<type>AA_AND2</type>
<position>252,-16.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1291</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-11</position>
<output>
<ID>OUT_0</ID>751 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1292</ID>
<type>AA_AND2</type>
<position>300,-16</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1293</ID>
<type>AE_DFF_LOW</type>
<position>349,-11</position>
<output>
<ID>OUT_0</ID>752 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1294</ID>
<type>AA_AND2</type>
<position>358.5,-18</position>
<input>
<ID>IN_0</ID>752 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1295</ID>
<type>AE_DFF_LOW</type>
<position>404,-11</position>
<output>
<ID>OUT_0</ID>753 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1296</ID>
<type>AA_AND2</type>
<position>412,-17</position>
<input>
<ID>IN_0</ID>753 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1297</ID>
<type>AE_DFF_LOW</type>
<position>461,-11</position>
<output>
<ID>OUT_0</ID>754 </output>
<input>
<ID>clock</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1298</ID>
<type>AA_AND2</type>
<position>470.5,-17.5</position>
<input>
<ID>IN_0</ID>754 </input>
<input>
<ID>IN_1</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1299</ID>
<type>AA_AND2</type>
<position>65,-10</position>
<output>
<ID>OUT</ID>748 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1300</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-28.5</position>
<output>
<ID>OUT_0</ID>755 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1301</ID>
<type>AA_AND2</type>
<position>106.5,-34</position>
<input>
<ID>IN_0</ID>755 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1302</ID>
<type>AE_DFF_LOW</type>
<position>146,-28.5</position>
<output>
<ID>OUT_0</ID>756 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1303</ID>
<type>AA_AND2</type>
<position>155,-35</position>
<input>
<ID>IN_0</ID>756 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1304</ID>
<type>AE_DFF_LOW</type>
<position>194,-28.5</position>
<output>
<ID>OUT_0</ID>758 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1305</ID>
<type>AA_AND2</type>
<position>201.5,-34</position>
<input>
<ID>IN_0</ID>758 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1306</ID>
<type>AE_DFF_LOW</type>
<position>243.5,-28.5</position>
<output>
<ID>OUT_0</ID>759 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1307</ID>
<type>AA_AND2</type>
<position>252,-34</position>
<input>
<ID>IN_0</ID>759 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1308</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-28.5</position>
<output>
<ID>OUT_0</ID>760 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1309</ID>
<type>AA_AND2</type>
<position>300,-33.5</position>
<input>
<ID>IN_0</ID>760 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1310</ID>
<type>AE_DFF_LOW</type>
<position>349,-28.5</position>
<output>
<ID>OUT_0</ID>761 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1311</ID>
<type>AA_AND2</type>
<position>358.5,-35.5</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1312</ID>
<type>AE_DFF_LOW</type>
<position>404,-28.5</position>
<output>
<ID>OUT_0</ID>762 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1313</ID>
<type>AA_AND2</type>
<position>412,-34.5</position>
<input>
<ID>IN_0</ID>762 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1314</ID>
<type>AE_DFF_LOW</type>
<position>461,-28.5</position>
<output>
<ID>OUT_0</ID>763 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1315</ID>
<type>AA_AND2</type>
<position>470.5,-35</position>
<input>
<ID>IN_0</ID>763 </input>
<input>
<ID>IN_1</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1316</ID>
<type>AA_AND2</type>
<position>65,-27.5</position>
<output>
<ID>OUT</ID>757 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1317</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-44.5</position>
<output>
<ID>OUT_0</ID>764 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1318</ID>
<type>AA_AND2</type>
<position>106.5,-50</position>
<input>
<ID>IN_0</ID>764 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1319</ID>
<type>AE_DFF_LOW</type>
<position>146,-44.5</position>
<output>
<ID>OUT_0</ID>765 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1320</ID>
<type>AA_AND2</type>
<position>155,-51</position>
<input>
<ID>IN_0</ID>765 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1321</ID>
<type>AE_DFF_LOW</type>
<position>194,-44.5</position>
<output>
<ID>OUT_0</ID>767 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1322</ID>
<type>AA_AND2</type>
<position>201.5,-50</position>
<input>
<ID>IN_0</ID>767 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1323</ID>
<type>AE_DFF_LOW</type>
<position>243.5,-44.5</position>
<output>
<ID>OUT_0</ID>768 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1324</ID>
<type>AA_AND2</type>
<position>252,-50</position>
<input>
<ID>IN_0</ID>768 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1325</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-44.5</position>
<output>
<ID>OUT_0</ID>769 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1326</ID>
<type>AA_AND2</type>
<position>300,-49.5</position>
<input>
<ID>IN_0</ID>769 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1327</ID>
<type>AE_DFF_LOW</type>
<position>349,-44.5</position>
<output>
<ID>OUT_0</ID>770 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1328</ID>
<type>AA_AND2</type>
<position>358.5,-51.5</position>
<input>
<ID>IN_0</ID>770 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1329</ID>
<type>AE_DFF_LOW</type>
<position>404,-44.5</position>
<output>
<ID>OUT_0</ID>771 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1330</ID>
<type>AA_AND2</type>
<position>412,-50.5</position>
<input>
<ID>IN_0</ID>771 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1331</ID>
<type>AE_DFF_LOW</type>
<position>461,-44.5</position>
<output>
<ID>OUT_0</ID>772 </output>
<input>
<ID>clock</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1332</ID>
<type>AA_AND2</type>
<position>470.5,-51</position>
<input>
<ID>IN_0</ID>772 </input>
<input>
<ID>IN_1</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1333</ID>
<type>AA_AND2</type>
<position>65,-43.5</position>
<output>
<ID>OUT</ID>766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1334</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-61</position>
<output>
<ID>OUT_0</ID>773 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1335</ID>
<type>AA_AND2</type>
<position>106.5,-66.5</position>
<input>
<ID>IN_0</ID>773 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1336</ID>
<type>AE_DFF_LOW</type>
<position>146,-61</position>
<output>
<ID>OUT_0</ID>774 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1337</ID>
<type>AA_AND2</type>
<position>155,-67.5</position>
<input>
<ID>IN_0</ID>774 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1338</ID>
<type>AE_DFF_LOW</type>
<position>194,-61</position>
<output>
<ID>OUT_0</ID>776 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1339</ID>
<type>AA_AND2</type>
<position>201.5,-66.5</position>
<input>
<ID>IN_0</ID>776 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1340</ID>
<type>AE_DFF_LOW</type>
<position>243.5,-61</position>
<output>
<ID>OUT_0</ID>777 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1341</ID>
<type>AA_AND2</type>
<position>252,-66.5</position>
<input>
<ID>IN_0</ID>777 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1342</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-61</position>
<output>
<ID>OUT_0</ID>778 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1343</ID>
<type>AA_AND2</type>
<position>300,-66</position>
<input>
<ID>IN_0</ID>778 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1344</ID>
<type>AE_DFF_LOW</type>
<position>349,-61</position>
<output>
<ID>OUT_0</ID>779 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1345</ID>
<type>AA_AND2</type>
<position>358.5,-68</position>
<input>
<ID>IN_0</ID>779 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1346</ID>
<type>AE_DFF_LOW</type>
<position>404,-61</position>
<output>
<ID>OUT_0</ID>780 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1347</ID>
<type>AA_AND2</type>
<position>412,-67</position>
<input>
<ID>IN_0</ID>780 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1348</ID>
<type>AE_DFF_LOW</type>
<position>461,-61</position>
<output>
<ID>OUT_0</ID>781 </output>
<input>
<ID>clock</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1349</ID>
<type>AA_AND2</type>
<position>470.5,-67.5</position>
<input>
<ID>IN_0</ID>781 </input>
<input>
<ID>IN_1</ID>775 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1350</ID>
<type>AA_AND2</type>
<position>65,-60</position>
<output>
<ID>OUT</ID>775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-50,467,-42.5</points>
<intersection>-50 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-50,467.5,-50</points>
<connection>
<GID>1332</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-42.5,467,-42.5</points>
<connection>
<GID>1331</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-65.5,101,-59</points>
<intersection>-65.5 1</intersection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-65.5,103.5,-65.5</points>
<connection>
<GID>1335</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-59,101,-59</points>
<connection>
<GID>1334</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-66.5,150,-59</points>
<intersection>-66.5 1</intersection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-66.5,152,-66.5</points>
<connection>
<GID>1337</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-59,150,-59</points>
<connection>
<GID>1336</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-60,467.5,-60</points>
<connection>
<GID>1350</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-67.5,102,-60</points>
<intersection>-67.5 5</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-67.5,103.5,-67.5</points>
<connection>
<GID>1335</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,-68.5,150.5,-60</points>
<intersection>-68.5 21</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,-68.5,152,-68.5</points>
<connection>
<GID>1337</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,-67.5,198,-60</points>
<intersection>-67.5 53</intersection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,-67.5,248.5,-60</points>
<intersection>-67.5 115</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,-67.5,198.5,-67.5</points>
<connection>
<GID>1339</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,-67,297,-60</points>
<connection>
<GID>1343</GID>
<name>IN_1</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,-69,355.5,-60</points>
<connection>
<GID>1345</GID>
<name>IN_1</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,-68,409.5,-60</points>
<intersection>-68 118</intersection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,-68.5,467.5,-60</points>
<connection>
<GID>1349</GID>
<name>IN_1</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,-62,93.5,-60</points>
<connection>
<GID>1334</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,-62,143,-60</points>
<connection>
<GID>1336</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,-62,191,-60</points>
<connection>
<GID>1338</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,-62,240.5,-60</points>
<connection>
<GID>1340</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,-62,288.5,-60</points>
<connection>
<GID>1342</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,-62,346,-60</points>
<connection>
<GID>1344</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,-62,401,-60</points>
<connection>
<GID>1346</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,-62,458,-60</points>
<connection>
<GID>1348</GID>
<name>clock</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,-67.5,249,-67.5</points>
<connection>
<GID>1341</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,-68,409.5,-68</points>
<connection>
<GID>1347</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-65.5,198.5,-59</points>
<connection>
<GID>1339</GID>
<name>IN_0</name></connection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-59,198.5,-59</points>
<connection>
<GID>1338</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-65.5,248,-59</points>
<intersection>-65.5 1</intersection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-65.5,249,-65.5</points>
<connection>
<GID>1341</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-59,248,-59</points>
<connection>
<GID>1340</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-65,296.5,-59</points>
<intersection>-65 5</intersection>
<intersection>-59 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-59,296.5,-59</points>
<connection>
<GID>1342</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,-65,297,-65</points>
<connection>
<GID>1343</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-67,355,-59</points>
<intersection>-67 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-67,355.5,-67</points>
<connection>
<GID>1345</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-59,355,-59</points>
<connection>
<GID>1344</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-66,408.5,-59</points>
<intersection>-66 4</intersection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,-59,408.5,-59</points>
<connection>
<GID>1346</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,-66,409,-66</points>
<connection>
<GID>1347</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-66.5,467,-59</points>
<intersection>-66.5 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-66.5,467.5,-66.5</points>
<connection>
<GID>1349</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-59,467,-59</points>
<connection>
<GID>1348</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-83.5,101,-77</points>
<intersection>-83.5 1</intersection>
<intersection>-77 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-83.5,103.5,-83.5</points>
<connection>
<GID>1352</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-77,101,-77</points>
<connection>
<GID>1351</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-84.5,150,-77</points>
<intersection>-84.5 1</intersection>
<intersection>-77 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-84.5,152,-84.5</points>
<connection>
<GID>1354</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-77,150,-77</points>
<connection>
<GID>1353</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-78,467.5,-78</points>
<connection>
<GID>1367</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-85.5,102,-78</points>
<intersection>-85.5 5</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-85.5,103.5,-85.5</points>
<connection>
<GID>1352</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,-86.5,150.5,-78</points>
<intersection>-86.5 21</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,-86.5,152,-86.5</points>
<connection>
<GID>1354</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,-85.5,198,-78</points>
<intersection>-85.5 53</intersection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,-85.5,248.5,-78</points>
<intersection>-85.5 115</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,-85.5,198.5,-85.5</points>
<connection>
<GID>1356</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,-85,297,-78</points>
<connection>
<GID>1360</GID>
<name>IN_1</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,-87,355.5,-78</points>
<connection>
<GID>1362</GID>
<name>IN_1</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,-86,409.5,-78</points>
<intersection>-86 118</intersection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,-86.5,467.5,-78</points>
<connection>
<GID>1366</GID>
<name>IN_1</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,-80,93.5,-78</points>
<connection>
<GID>1351</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,-80,143,-78</points>
<connection>
<GID>1353</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,-80,191,-78</points>
<connection>
<GID>1355</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,-80,240.5,-78</points>
<connection>
<GID>1357</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,-80,288.5,-78</points>
<connection>
<GID>1359</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,-80,346,-78</points>
<connection>
<GID>1361</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,-80,401,-78</points>
<connection>
<GID>1363</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,-80,458,-78</points>
<connection>
<GID>1365</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,-85.5,249,-85.5</points>
<connection>
<GID>1358</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,-86,409.5,-86</points>
<connection>
<GID>1364</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-83.5,198.5,-77</points>
<connection>
<GID>1356</GID>
<name>IN_0</name></connection>
<intersection>-77 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-77,198.5,-77</points>
<connection>
<GID>1355</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-83.5,248,-77</points>
<intersection>-83.5 1</intersection>
<intersection>-77 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-83.5,249,-83.5</points>
<connection>
<GID>1358</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-77,248,-77</points>
<connection>
<GID>1357</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-83,296.5,-77</points>
<intersection>-83 5</intersection>
<intersection>-77 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-77,296.5,-77</points>
<connection>
<GID>1359</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,-83,297,-83</points>
<connection>
<GID>1360</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-85,355,-77</points>
<intersection>-85 1</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-85,355.5,-85</points>
<connection>
<GID>1362</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-77,355,-77</points>
<connection>
<GID>1361</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-84,408.5,-77</points>
<intersection>-84 4</intersection>
<intersection>-77 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,-77,408.5,-77</points>
<connection>
<GID>1363</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,-84,409,-84</points>
<connection>
<GID>1364</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-84.5,467,-77</points>
<intersection>-84.5 1</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-84.5,467.5,-84.5</points>
<connection>
<GID>1366</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-77,467,-77</points>
<connection>
<GID>1365</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-105.5,101,-99</points>
<intersection>-105.5 1</intersection>
<intersection>-99 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-105.5,103.5,-105.5</points>
<connection>
<GID>1369</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-99,101,-99</points>
<connection>
<GID>1368</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-106.5,150,-99</points>
<intersection>-106.5 1</intersection>
<intersection>-99 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-106.5,152,-106.5</points>
<connection>
<GID>1371</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-99,150,-99</points>
<connection>
<GID>1370</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-100,467.5,-100</points>
<connection>
<GID>1384</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-107.5,102,-100</points>
<intersection>-107.5 5</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-107.5,103.5,-107.5</points>
<connection>
<GID>1369</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,-108.5,150.5,-100</points>
<intersection>-108.5 21</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,-108.5,152,-108.5</points>
<connection>
<GID>1371</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,-107.5,198,-100</points>
<intersection>-107.5 53</intersection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,-107.5,248.5,-100</points>
<intersection>-107.5 115</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,-107.5,198.5,-107.5</points>
<connection>
<GID>1373</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,-107,297,-100</points>
<connection>
<GID>1377</GID>
<name>IN_1</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,-109,355.5,-100</points>
<connection>
<GID>1379</GID>
<name>IN_1</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,-108,409.5,-100</points>
<intersection>-108 118</intersection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,-108.5,467.5,-100</points>
<connection>
<GID>1383</GID>
<name>IN_1</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,-102,93.5,-100</points>
<connection>
<GID>1368</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,-102,143,-100</points>
<connection>
<GID>1370</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,-102,191,-100</points>
<connection>
<GID>1372</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,-102,240.5,-100</points>
<connection>
<GID>1374</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,-102,288.5,-100</points>
<connection>
<GID>1376</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,-102,346,-100</points>
<connection>
<GID>1378</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,-102,401,-100</points>
<connection>
<GID>1380</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,-102,458,-100</points>
<connection>
<GID>1382</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,-107.5,249,-107.5</points>
<connection>
<GID>1375</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,-108,409.5,-108</points>
<connection>
<GID>1381</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-105.5,198.5,-99</points>
<connection>
<GID>1373</GID>
<name>IN_0</name></connection>
<intersection>-99 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-99,198.5,-99</points>
<connection>
<GID>1372</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-105.5,248,-99</points>
<intersection>-105.5 1</intersection>
<intersection>-99 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-105.5,249,-105.5</points>
<connection>
<GID>1375</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-99,248,-99</points>
<connection>
<GID>1374</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-105,296.5,-99</points>
<intersection>-105 5</intersection>
<intersection>-99 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-99,296.5,-99</points>
<connection>
<GID>1376</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,-105,297,-105</points>
<connection>
<GID>1377</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-107,355,-99</points>
<intersection>-107 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-107,355.5,-107</points>
<connection>
<GID>1379</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-99,355,-99</points>
<connection>
<GID>1378</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-106,408.5,-99</points>
<intersection>-106 4</intersection>
<intersection>-99 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,-99,408.5,-99</points>
<connection>
<GID>1380</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,-106,409,-106</points>
<connection>
<GID>1381</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-106.5,467,-99</points>
<intersection>-106.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-106.5,467.5,-106.5</points>
<connection>
<GID>1383</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-99,467,-99</points>
<connection>
<GID>1382</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,21.5,101,28</points>
<intersection>21.5 1</intersection>
<intersection>28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,21.5,103.5,21.5</points>
<connection>
<GID>1251</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,28,101,28</points>
<connection>
<GID>1250</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,20.5,150,28</points>
<intersection>20.5 1</intersection>
<intersection>28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,20.5,152,20.5</points>
<connection>
<GID>1253</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149,28,150,28</points>
<connection>
<GID>1252</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,27,467.5,27</points>
<connection>
<GID>1249</GID>
<name>OUT</name></connection>
<intersection>93.5 82</intersection>
<intersection>101.5 4</intersection>
<intersection>143 80</intersection>
<intersection>150.5 16</intersection>
<intersection>191 81</intersection>
<intersection>199 23</intersection>
<intersection>240.5 79</intersection>
<intersection>248 31</intersection>
<intersection>288.5 83</intersection>
<intersection>297 55</intersection>
<intersection>346 84</intersection>
<intersection>355.5 56</intersection>
<intersection>401 78</intersection>
<intersection>407.5 66</intersection>
<intersection>458 85</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>101.5,19.5,101.5,27</points>
<intersection>19.5 5</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>101.5,19.5,103.5,19.5</points>
<connection>
<GID>1251</GID>
<name>IN_1</name></connection>
<intersection>101.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,18.5,150.5,27</points>
<intersection>18.5 21</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,18.5,152,18.5</points>
<connection>
<GID>1253</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>199,19.5,199,27</points>
<intersection>19.5 53</intersection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248,20,248,27</points>
<connection>
<GID>1257</GID>
<name>IN_1</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198.5,19.5,199,19.5</points>
<connection>
<GID>1255</GID>
<name>IN_1</name></connection>
<intersection>199 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,20,297,27</points>
<connection>
<GID>1259</GID>
<name>IN_1</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,18,355.5,27</points>
<connection>
<GID>1261</GID>
<name>IN_1</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>407.5,18.5,407.5,27</points>
<connection>
<GID>1263</GID>
<name>IN_1</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,18.5,467.5,27</points>
<connection>
<GID>1265</GID>
<name>IN_1</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>401,25,401,27</points>
<connection>
<GID>1262</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>79</ID>
<points>240.5,25,240.5,27</points>
<connection>
<GID>1256</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>80</ID>
<points>143,25,143,27</points>
<connection>
<GID>1252</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>81</ID>
<points>191,25,191,27</points>
<connection>
<GID>1254</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>82</ID>
<points>93.5,25,93.5,27</points>
<connection>
<GID>1250</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>83</ID>
<points>288.5,25,288.5,27</points>
<connection>
<GID>1258</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>84</ID>
<points>346,25,346,27</points>
<connection>
<GID>1260</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment>
<vsegment>
<ID>85</ID>
<points>458,25,458,27</points>
<connection>
<GID>1264</GID>
<name>clock</name></connection>
<intersection>27 1</intersection></vsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,21.5,198.5,28</points>
<connection>
<GID>1255</GID>
<name>IN_0</name></connection>
<intersection>28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197,28,198.5,28</points>
<connection>
<GID>1254</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,22,247.5,28</points>
<intersection>22 1</intersection>
<intersection>28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247.5,22,248,22</points>
<connection>
<GID>1257</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>246.5,28,247.5,28</points>
<connection>
<GID>1256</GID>
<name>OUT_0</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,22,296.5,28</points>
<intersection>22 5</intersection>
<intersection>28 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,28,296.5,28</points>
<connection>
<GID>1258</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,22,297,22</points>
<connection>
<GID>1259</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,20,355,28</points>
<intersection>20 1</intersection>
<intersection>28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,20,355.5,20</points>
<connection>
<GID>1261</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,28,355,28</points>
<connection>
<GID>1260</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407,20.5,407,28</points>
<connection>
<GID>1262</GID>
<name>OUT_0</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>407,20.5,407.5,20.5</points>
<connection>
<GID>1263</GID>
<name>IN_0</name></connection>
<intersection>407 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,20.5,467,28</points>
<intersection>20.5 1</intersection>
<intersection>28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,20.5,467.5,20.5</points>
<connection>
<GID>1265</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,28,467,28</points>
<connection>
<GID>1264</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,3.5,101,10</points>
<intersection>3.5 1</intersection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,3.5,103.5,3.5</points>
<connection>
<GID>1267</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,10,101,10</points>
<connection>
<GID>1266</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,2.5,150,10</points>
<intersection>2.5 1</intersection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,2.5,152,2.5</points>
<connection>
<GID>1269</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,10,150,10</points>
<connection>
<GID>1268</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,9,467.5,9</points>
<connection>
<GID>1282</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,1.5,102,9</points>
<intersection>1.5 5</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,1.5,103.5,1.5</points>
<connection>
<GID>1267</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,0.5,150.5,9</points>
<intersection>0.5 21</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,0.5,152,0.5</points>
<connection>
<GID>1269</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,1.5,198,9</points>
<intersection>1.5 53</intersection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,1.5,248.5,9</points>
<intersection>1.5 115</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,1.5,198.5,1.5</points>
<connection>
<GID>1271</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,2,297,9</points>
<connection>
<GID>1275</GID>
<name>IN_1</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,0,355.5,9</points>
<connection>
<GID>1277</GID>
<name>IN_1</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,1,409.5,9</points>
<intersection>1 118</intersection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,0.5,467.5,9</points>
<connection>
<GID>1281</GID>
<name>IN_1</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,7,93.5,9</points>
<connection>
<GID>1266</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,7,143,9</points>
<connection>
<GID>1268</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,7,191,9</points>
<connection>
<GID>1270</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,7,240.5,9</points>
<connection>
<GID>1272</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,7,288.5,9</points>
<connection>
<GID>1274</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,7,346,9</points>
<connection>
<GID>1276</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,7,401,9</points>
<connection>
<GID>1278</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,7,458,9</points>
<connection>
<GID>1280</GID>
<name>clock</name></connection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,1.5,249,1.5</points>
<connection>
<GID>1273</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,1,409.5,1</points>
<connection>
<GID>1279</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,3.5,198.5,10</points>
<connection>
<GID>1271</GID>
<name>IN_0</name></connection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,10,198.5,10</points>
<connection>
<GID>1270</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,3.5,248,10</points>
<intersection>3.5 1</intersection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,3.5,249,3.5</points>
<connection>
<GID>1273</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,10,248,10</points>
<connection>
<GID>1272</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,4,296.5,10</points>
<intersection>4 5</intersection>
<intersection>10 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,10,296.5,10</points>
<connection>
<GID>1274</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,4,297,4</points>
<connection>
<GID>1275</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,2,355,10</points>
<intersection>2 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,2,355.5,2</points>
<connection>
<GID>1277</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,10,355,10</points>
<connection>
<GID>1276</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,3,408.5,10</points>
<intersection>3 4</intersection>
<intersection>10 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,10,408.5,10</points>
<connection>
<GID>1278</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,3,409,3</points>
<connection>
<GID>1279</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,2.5,467,10</points>
<intersection>2.5 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,2.5,467.5,2.5</points>
<connection>
<GID>1281</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,10,467,10</points>
<connection>
<GID>1280</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-15.5,101,-9</points>
<intersection>-15.5 1</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-15.5,103.5,-15.5</points>
<connection>
<GID>1284</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-9,101,-9</points>
<connection>
<GID>1283</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-16.5,150,-9</points>
<intersection>-16.5 1</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-16.5,152,-16.5</points>
<connection>
<GID>1286</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-9,150,-9</points>
<connection>
<GID>1285</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-10,467.5,-10</points>
<connection>
<GID>1299</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-17.5,102,-10</points>
<intersection>-17.5 5</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-17.5,103.5,-17.5</points>
<connection>
<GID>1284</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,-18.5,150.5,-10</points>
<intersection>-18.5 21</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,-18.5,152,-18.5</points>
<connection>
<GID>1286</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,-17.5,198,-10</points>
<intersection>-17.5 53</intersection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,-17.5,248.5,-10</points>
<intersection>-17.5 115</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,-17.5,198.5,-17.5</points>
<connection>
<GID>1288</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,-17,297,-10</points>
<connection>
<GID>1292</GID>
<name>IN_1</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,-19,355.5,-10</points>
<connection>
<GID>1294</GID>
<name>IN_1</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,-18,409.5,-10</points>
<intersection>-18 118</intersection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,-18.5,467.5,-10</points>
<connection>
<GID>1298</GID>
<name>IN_1</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,-12,93.5,-10</points>
<connection>
<GID>1283</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,-12,143,-10</points>
<connection>
<GID>1285</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,-12,191,-10</points>
<connection>
<GID>1287</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,-12,240.5,-10</points>
<connection>
<GID>1289</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,-12,288.5,-10</points>
<connection>
<GID>1291</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,-12,346,-10</points>
<connection>
<GID>1293</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,-12,401,-10</points>
<connection>
<GID>1295</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,-12,458,-10</points>
<connection>
<GID>1297</GID>
<name>clock</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,-17.5,249,-17.5</points>
<connection>
<GID>1290</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,-18,409.5,-18</points>
<connection>
<GID>1296</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-15.5,198.5,-9</points>
<connection>
<GID>1288</GID>
<name>IN_0</name></connection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-9,198.5,-9</points>
<connection>
<GID>1287</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-15.5,248,-9</points>
<intersection>-15.5 1</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-15.5,249,-15.5</points>
<connection>
<GID>1290</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-9,248,-9</points>
<connection>
<GID>1289</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-15,296.5,-9</points>
<intersection>-15 5</intersection>
<intersection>-9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-9,296.5,-9</points>
<connection>
<GID>1291</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,-15,297,-15</points>
<connection>
<GID>1292</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-17,355,-9</points>
<intersection>-17 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-17,355.5,-17</points>
<connection>
<GID>1294</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-9,355,-9</points>
<connection>
<GID>1293</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-16,408.5,-9</points>
<intersection>-16 4</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,-9,408.5,-9</points>
<connection>
<GID>1295</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,-16,409,-16</points>
<connection>
<GID>1296</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-16.5,467,-9</points>
<intersection>-16.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-16.5,467.5,-16.5</points>
<connection>
<GID>1298</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-9,467,-9</points>
<connection>
<GID>1297</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-33,101,-26.5</points>
<intersection>-33 1</intersection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-33,103.5,-33</points>
<connection>
<GID>1301</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-26.5,101,-26.5</points>
<connection>
<GID>1300</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-34,150,-26.5</points>
<intersection>-34 1</intersection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-34,152,-34</points>
<connection>
<GID>1303</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-26.5,150,-26.5</points>
<connection>
<GID>1302</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-27.5,467.5,-27.5</points>
<connection>
<GID>1316</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-35,102,-27.5</points>
<intersection>-35 5</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-35,103.5,-35</points>
<connection>
<GID>1301</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,-36,150.5,-27.5</points>
<intersection>-36 21</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,-36,152,-36</points>
<connection>
<GID>1303</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,-35,198,-27.5</points>
<intersection>-35 53</intersection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,-35,248.5,-27.5</points>
<intersection>-35 115</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,-35,198.5,-35</points>
<connection>
<GID>1305</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,-34.5,297,-27.5</points>
<connection>
<GID>1309</GID>
<name>IN_1</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,-36.5,355.5,-27.5</points>
<connection>
<GID>1311</GID>
<name>IN_1</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,-35.5,409.5,-27.5</points>
<intersection>-35.5 118</intersection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,-36,467.5,-27.5</points>
<connection>
<GID>1315</GID>
<name>IN_1</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,-29.5,93.5,-27.5</points>
<connection>
<GID>1300</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,-29.5,143,-27.5</points>
<connection>
<GID>1302</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,-29.5,191,-27.5</points>
<connection>
<GID>1304</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,-29.5,240.5,-27.5</points>
<connection>
<GID>1306</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,-29.5,288.5,-27.5</points>
<connection>
<GID>1308</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,-29.5,346,-27.5</points>
<connection>
<GID>1310</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,-29.5,401,-27.5</points>
<connection>
<GID>1312</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,-29.5,458,-27.5</points>
<connection>
<GID>1314</GID>
<name>clock</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,-35,249,-35</points>
<connection>
<GID>1307</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,-35.5,409.5,-35.5</points>
<connection>
<GID>1313</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-33,198.5,-26.5</points>
<connection>
<GID>1305</GID>
<name>IN_0</name></connection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-26.5,198.5,-26.5</points>
<connection>
<GID>1304</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-33,248,-26.5</points>
<intersection>-33 1</intersection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-33,249,-33</points>
<connection>
<GID>1307</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-26.5,248,-26.5</points>
<connection>
<GID>1306</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-32.5,296.5,-26.5</points>
<intersection>-32.5 5</intersection>
<intersection>-26.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-26.5,296.5,-26.5</points>
<connection>
<GID>1308</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,-32.5,297,-32.5</points>
<connection>
<GID>1309</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-34.5,355,-26.5</points>
<intersection>-34.5 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-34.5,355.5,-34.5</points>
<connection>
<GID>1311</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-26.5,355,-26.5</points>
<connection>
<GID>1310</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-33.5,408.5,-26.5</points>
<intersection>-33.5 4</intersection>
<intersection>-26.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,-26.5,408.5,-26.5</points>
<connection>
<GID>1312</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,-33.5,409,-33.5</points>
<connection>
<GID>1313</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-34,467,-26.5</points>
<intersection>-34 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-34,467.5,-34</points>
<connection>
<GID>1315</GID>
<name>IN_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-26.5,467,-26.5</points>
<connection>
<GID>1314</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-49,101,-42.5</points>
<intersection>-49 1</intersection>
<intersection>-42.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-49,103.5,-49</points>
<connection>
<GID>1318</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-42.5,101,-42.5</points>
<connection>
<GID>1317</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-50,150,-42.5</points>
<intersection>-50 1</intersection>
<intersection>-42.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-50,152,-50</points>
<connection>
<GID>1320</GID>
<name>IN_0</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149,-42.5,150,-42.5</points>
<connection>
<GID>1319</GID>
<name>OUT_0</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-43.5,467.5,-43.5</points>
<connection>
<GID>1333</GID>
<name>OUT</name></connection>
<intersection>93.5 107</intersection>
<intersection>102 4</intersection>
<intersection>143 108</intersection>
<intersection>150.5 16</intersection>
<intersection>191 109</intersection>
<intersection>198 23</intersection>
<intersection>240.5 110</intersection>
<intersection>248.5 31</intersection>
<intersection>288.5 111</intersection>
<intersection>297 55</intersection>
<intersection>346 112</intersection>
<intersection>355.5 56</intersection>
<intersection>401 113</intersection>
<intersection>409.5 66</intersection>
<intersection>458 114</intersection>
<intersection>467.5 77</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-51,102,-43.5</points>
<intersection>-51 5</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-51,103.5,-51</points>
<connection>
<GID>1318</GID>
<name>IN_1</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>150.5,-52,150.5,-43.5</points>
<intersection>-52 21</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>150.5,-52,152,-52</points>
<connection>
<GID>1320</GID>
<name>IN_1</name></connection>
<intersection>150.5 16</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>198,-51,198,-43.5</points>
<intersection>-51 53</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>248.5,-51,248.5,-43.5</points>
<intersection>-51 115</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>198,-51,198.5,-51</points>
<connection>
<GID>1322</GID>
<name>IN_1</name></connection>
<intersection>198 23</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>297,-50.5,297,-43.5</points>
<connection>
<GID>1326</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>355.5,-52.5,355.5,-43.5</points>
<connection>
<GID>1328</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>409.5,-51.5,409.5,-43.5</points>
<intersection>-51.5 118</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>467.5,-52,467.5,-43.5</points>
<connection>
<GID>1332</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>93.5,-45.5,93.5,-43.5</points>
<connection>
<GID>1317</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>143,-45.5,143,-43.5</points>
<connection>
<GID>1319</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>191,-45.5,191,-43.5</points>
<connection>
<GID>1321</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>240.5,-45.5,240.5,-43.5</points>
<connection>
<GID>1323</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>288.5,-45.5,288.5,-43.5</points>
<connection>
<GID>1325</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>346,-45.5,346,-43.5</points>
<connection>
<GID>1327</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>401,-45.5,401,-43.5</points>
<connection>
<GID>1329</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>458,-45.5,458,-43.5</points>
<connection>
<GID>1331</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>115</ID>
<points>248.5,-51,249,-51</points>
<connection>
<GID>1324</GID>
<name>IN_1</name></connection>
<intersection>248.5 31</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>409,-51.5,409.5,-51.5</points>
<connection>
<GID>1330</GID>
<name>IN_1</name></connection>
<intersection>409.5 66</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-49,198.5,-42.5</points>
<connection>
<GID>1322</GID>
<name>IN_0</name></connection>
<intersection>-42.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>197,-42.5,198.5,-42.5</points>
<connection>
<GID>1321</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-49,248,-42.5</points>
<intersection>-49 1</intersection>
<intersection>-42.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-49,249,-49</points>
<connection>
<GID>1324</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>246.5,-42.5,248,-42.5</points>
<connection>
<GID>1323</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-48.5,296.5,-42.5</points>
<intersection>-48.5 5</intersection>
<intersection>-42.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>294.5,-42.5,296.5,-42.5</points>
<connection>
<GID>1325</GID>
<name>OUT_0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>296.5,-48.5,297,-48.5</points>
<connection>
<GID>1326</GID>
<name>IN_0</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-50.5,355,-42.5</points>
<intersection>-50.5 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-50.5,355.5,-50.5</points>
<connection>
<GID>1328</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-42.5,355,-42.5</points>
<connection>
<GID>1327</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-49.5,408.5,-42.5</points>
<intersection>-49.5 4</intersection>
<intersection>-42.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407,-42.5,408.5,-42.5</points>
<connection>
<GID>1329</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>408.5,-49.5,409,-49.5</points>
<connection>
<GID>1330</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>186.987,362.142,404.833,254.465</PageViewport>
<gate>
<ID>193</ID>
<type>BA_TRI_STATE</type>
<position>346.5,176</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>194</ID>
<type>BA_TRI_STATE</type>
<position>394,173.5</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>BA_TRI_STATE</type>
<position>442.5,173.5</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_TRI_STATE</type>
<position>497.5,175</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>BA_TRI_STATE</type>
<position>553.5,174.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>199</ID>
<type>BA_TRI_STATE</type>
<position>615.5,173</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>228,309</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_TOGGLE</type>
<position>214,193</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>247,160.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_TOGGLE</type>
<position>299,160</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_TOGGLE</type>
<position>346,159.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_TOGGLE</type>
<position>393.5,160</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_TOGGLE</type>
<position>443,160.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>498,160.5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_TOGGLE</type>
<position>554,160</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_TOGGLE</type>
<position>615,160.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>211</ID>
<type>BA_TRI_STATE</type>
<position>238.5,212</position>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>213</ID>
<type>BA_TRI_STATE</type>
<position>240.5,240.5</position>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>BA_TRI_STATE</type>
<position>239,273</position>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>215</ID>
<type>BA_TRI_STATE</type>
<position>239.5,304.5</position>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_DFF_LOW</type>
<position>259.5,310</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>31 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>269.5,304.5</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_DFF_LOW</type>
<position>309,310</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>318,303.5</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AE_DFF_LOW</type>
<position>357,310</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_AND2</type>
<position>364.5,304.5</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_DFF_LOW</type>
<position>406.5,310</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>36 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>414,305</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_DFF_LOW</type>
<position>454.5,310</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_AND2</type>
<position>463,305</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_DFF_LOW</type>
<position>512,310</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>521.5,303</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_DFF_LOW</type>
<position>567,310</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>573.5,303.5</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_DFF_LOW</type>
<position>624,310</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>633.5,303.5</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>226.5,337.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>252,346.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>294.5,346.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>345,346.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>398.5,346.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>464,345.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>525.5,344</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>576,342.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>630,340</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>BA_TRI_STATE</type>
<position>476,305</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>91</ID>
<type>BA_TRI_STATE</type>
<position>536,303</position>
<input>
<ID>ENABLE_0</ID>117 </input>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>BA_TRI_STATE</type>
<position>595,304</position>
<input>
<ID>ENABLE_0</ID>118 </input>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>BA_TRI_STATE</type>
<position>650.5,303.5</position>
<input>
<ID>ENABLE_0</ID>125 </input>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>94</ID>
<type>BA_TRI_STATE</type>
<position>429,304.5</position>
<input>
<ID>ENABLE_0</ID>105 </input>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>97</ID>
<type>BA_TRI_STATE</type>
<position>380.5,303.5</position>
<input>
<ID>ENABLE_0</ID>101 </input>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_TRI_STATE</type>
<position>331.5,304.5</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>BA_TRI_STATE</type>
<position>285.5,304</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>100</ID>
<type>BA_TRI_STATE</type>
<position>290.5,338</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>BA_TRI_STATE</type>
<position>337.5,336.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>BA_TRI_STATE</type>
<position>384.5,337</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>BA_TRI_STATE</type>
<position>434.5,337.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>BA_TRI_STATE</type>
<position>482,337.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>BA_TRI_STATE</type>
<position>541,336</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_TRI_STATE</type>
<position>598.5,331.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>108</ID>
<type>BA_TRI_STATE</type>
<position>654.5,329.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>112</ID>
<type>BA_DECODER_2x4</type>
<position>201.5,308.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>71 </output>
<output>
<ID>OUT_3</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>227,276.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_DFF_LOW</type>
<position>258.5,277.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>268.5,272</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_DFF_LOW</type>
<position>308,277.5</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>317,271</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_DFF_LOW</type>
<position>356,277.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>363.5,272</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_DFF_LOW</type>
<position>405.5,277.5</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>413,272.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AE_DFF_LOW</type>
<position>453.5,277.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND2</type>
<position>462,273</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AE_DFF_LOW</type>
<position>511,277.5</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>520.5,270.5</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AE_DFF_LOW</type>
<position>566,277.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>572.5,271</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>AE_DFF_LOW</type>
<position>623,277.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>632.5,271</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>BA_TRI_STATE</type>
<position>475,272.5</position>
<input>
<ID>ENABLE_0</ID>111 </input>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>131</ID>
<type>BA_TRI_STATE</type>
<position>534.5,271</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>BA_TRI_STATE</type>
<position>594,270.5</position>
<input>
<ID>ENABLE_0</ID>119 </input>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>133</ID>
<type>BA_TRI_STATE</type>
<position>649,270.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_TRI_STATE</type>
<position>428,272</position>
<input>
<ID>ENABLE_0</ID>107 </input>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>135</ID>
<type>BA_TRI_STATE</type>
<position>379.5,271</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>BA_TRI_STATE</type>
<position>286,271</position>
<input>
<ID>ENABLE_0</ID>95 </input>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>BA_TRI_STATE</type>
<position>332,270</position>
<input>
<ID>ENABLE_0</ID>98 </input>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_AND2</type>
<position>226,244</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AE_DFF_LOW</type>
<position>257.5,245.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND2</type>
<position>267.5,240</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>AE_DFF_LOW</type>
<position>307,245.5</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND2</type>
<position>316,239</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_DFF_LOW</type>
<position>355,245.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>362.5,240</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_DFF_LOW</type>
<position>404.5,245.5</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>55 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND2</type>
<position>417,240</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_DFF_LOW</type>
<position>452.5,245.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>56 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND2</type>
<position>461,240.5</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AE_DFF_LOW</type>
<position>510,245.5</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>57 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>519.5,238.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_DFF_LOW</type>
<position>565,245.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_AND2</type>
<position>571.5,239</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AE_DFF_LOW</type>
<position>622,245.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND2</type>
<position>631.5,239</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>BA_TRI_STATE</type>
<position>474,240.5</position>
<input>
<ID>ENABLE_0</ID>112 </input>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>BA_TRI_STATE</type>
<position>531.5,239</position>
<input>
<ID>ENABLE_0</ID>115 </input>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>BA_TRI_STATE</type>
<position>593,238.5</position>
<input>
<ID>ENABLE_0</ID>120 </input>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>158</ID>
<type>BA_TRI_STATE</type>
<position>648.5,238.5</position>
<input>
<ID>ENABLE_0</ID>123 </input>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>BA_TRI_STATE</type>
<position>427,240</position>
<input>
<ID>ENABLE_0</ID>108 </input>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>160</ID>
<type>BA_TRI_STATE</type>
<position>378.5,239</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>161</ID>
<type>BA_TRI_STATE</type>
<position>328,239</position>
<input>
<ID>ENABLE_0</ID>99 </input>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>BA_TRI_STATE</type>
<position>286.5,239.5</position>
<input>
<ID>ENABLE_0</ID>93 </input>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_AND2</type>
<position>226,217</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_DFF_LOW</type>
<position>257.5,218</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>61 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_AND2</type>
<position>267.5,212.5</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_DFF_LOW</type>
<position>307,218</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>62 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_AND2</type>
<position>316,211.5</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_DFF_LOW</type>
<position>355,218</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>63 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND2</type>
<position>362.5,212.5</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AE_DFF_LOW</type>
<position>404.5,218</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND2</type>
<position>412,213</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AE_DFF_LOW</type>
<position>452.5,218</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>461,213</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AE_DFF_LOW</type>
<position>510,218</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>519.5,211</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_DFF_LOW</type>
<position>565,218</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND2</type>
<position>571.5,211.5</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_DFF_LOW</type>
<position>622,218</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND2</type>
<position>631.5,211.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>BA_TRI_STATE</type>
<position>474,213</position>
<input>
<ID>ENABLE_0</ID>113 </input>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>181</ID>
<type>BA_TRI_STATE</type>
<position>534,212</position>
<input>
<ID>ENABLE_0</ID>114 </input>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>BA_TRI_STATE</type>
<position>593,211.5</position>
<input>
<ID>ENABLE_0</ID>121 </input>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>183</ID>
<type>BA_TRI_STATE</type>
<position>651.5,214</position>
<input>
<ID>ENABLE_0</ID>122 </input>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>184</ID>
<type>BA_TRI_STATE</type>
<position>427,212.5</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>185</ID>
<type>BA_TRI_STATE</type>
<position>378.5,211.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>186</ID>
<type>BA_TRI_STATE</type>
<position>328,211.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>BA_TRI_STATE</type>
<position>286.5,212</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>215.5,176.5</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>191</ID>
<type>BA_TRI_STATE</type>
<position>249.5,176.5</position>
<input>
<ID>ENABLE_0</ID>75 </input>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>BA_TRI_STATE</type>
<position>298.5,176</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,300,264,312</points>
<intersection>300 1</intersection>
<intersection>305.5 5</intersection>
<intersection>312 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264,300,285.5,300</points>
<intersection>264 0</intersection>
<intersection>285.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>262.5,312,264,312</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>264 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>285.5,300,285.5,301</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>300 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>264,305.5,266.5,305.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>264 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,299.5,313,312</points>
<intersection>299.5 1</intersection>
<intersection>304.5 5</intersection>
<intersection>312 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,299.5,331.5,299.5</points>
<intersection>313 0</intersection>
<intersection>331.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>312,312,313,312</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>313 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>331.5,299.5,331.5,301.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>299.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>313,304.5,315,304.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434,215,434,274.5</points>
<intersection>215 3</intersection>
<intersection>242.5 4</intersection>
<intersection>274.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>434.5,274.5,434.5,334.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>274.5 2</intersection>
<intersection>307 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>428,274.5,434.5,274.5</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>434 0</intersection>
<intersection>434.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427,215,434,215</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>427,242.5,434,242.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>429,307,434.5,307</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>434.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359.5,300.5,359.5,312</points>
<intersection>300.5 4</intersection>
<intersection>305.5 5</intersection>
<intersection>312 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>359.5,312,360,312</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>359.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>359.5,300.5,380.5,300.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>359.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>359.5,305.5,361.5,305.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>359.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410.5,300.5,410.5,312</points>
<intersection>300.5 1</intersection>
<intersection>306 5</intersection>
<intersection>312 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>410.5,300.5,429,300.5</points>
<intersection>410.5 0</intersection>
<intersection>429 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>409.5,312,410.5,312</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>410.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>429,300.5,429,301.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>300.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>410.5,306,411,306</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>410.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,300,458,306.5</points>
<intersection>300 5</intersection>
<intersection>306 9</intersection>
<intersection>306.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>457.5,306.5,458,306.5</points>
<intersection>457.5 6</intersection>
<intersection>458 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>458,300,476,300</points>
<intersection>458 0</intersection>
<intersection>476 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>457.5,306.5,457.5,312</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>306.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>476,300,476,302</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>300 5</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>458,306,460,306</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>458 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518,304,518,312</points>
<intersection>304 1</intersection>
<intersection>312 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>518,304,536,304</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>518 0</intersection>
<intersection>536 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515,312,518,312</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>518 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>536,300,536,304</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>304 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570,304.5,570,312</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>304.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>570,304.5,595,304.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>570 0</intersection>
<intersection>595 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>595,301,595,304.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>304.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>630,304.5,630,312</points>
<intersection>304.5 1</intersection>
<intersection>312 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>630,304.5,650.5,304.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>630 0</intersection>
<intersection>650.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>627,312,630,312</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>630 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>650.5,300.5,650.5,304.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>304.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>231,309,621,309</points>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<connection>
<GID>64</GID>
<name>clock</name></connection>
<connection>
<GID>62</GID>
<name>clock</name></connection>
<connection>
<GID>60</GID>
<name>clock</name></connection>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<connection>
<GID>8</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>385.5,214,385.5,274</points>
<intersection>214 3</intersection>
<intersection>241.5 4</intersection>
<intersection>274 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>384.5,273.5,384.5,334</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>273.5 5</intersection>
<intersection>274 2</intersection>
<intersection>306 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>384.5,274,385.5,274</points>
<intersection>384.5 1</intersection>
<intersection>385.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>378.5,214,385.5,214</points>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection>
<intersection>385.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>378.5,241.5,385.5,241.5</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>385.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>379.5,273.5,384.5,273.5</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>384.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380.5,306,384.5,306</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>384.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,267,263,279.5</points>
<intersection>267 1</intersection>
<intersection>273 5</intersection>
<intersection>279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,267,286,267</points>
<intersection>263 0</intersection>
<intersection>286 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>261.5,279.5,263,279.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>263 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>286,267,286,268</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>267 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>263,273,265.5,273</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>263 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,266,312,279.5</points>
<intersection>266 1</intersection>
<intersection>279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,266,332,266</points>
<intersection>311.5 4</intersection>
<intersection>312 0</intersection>
<intersection>332 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>311,279.5,312,279.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>312 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>332,266,332,267</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>266 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>311.5,266,311.5,272</points>
<intersection>266 1</intersection>
<intersection>272 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>311.5,272,314,272</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>311.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358.5,268,358.5,279</points>
<intersection>268 7</intersection>
<intersection>273 8</intersection>
<intersection>279 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>358.5,279,359,279</points>
<intersection>358.5 0</intersection>
<intersection>359 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>359,279,359,279.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>279 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>358.5,268,379.5,268</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>358.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>358.5,273,360.5,273</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>358.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>409,268.5,409,279.5</points>
<intersection>268.5 1</intersection>
<intersection>273.5 5</intersection>
<intersection>279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>409,268.5,428,268.5</points>
<intersection>409 0</intersection>
<intersection>428 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>408.5,279.5,409,279.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>409 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>428,268.5,428,269</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>268.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>409,273.5,410,273.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>409 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>454.5,268,475,268</points>
<intersection>454.5 8</intersection>
<intersection>456.5 6</intersection>
<intersection>475 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>456.5,268,456.5,279.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>268 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>475,268,475,269.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>268 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>454.5,268,454.5,274</points>
<intersection>268 4</intersection>
<intersection>274 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>454.5,274,459,274</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>454.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,271.5,517,279.5</points>
<intersection>271.5 1</intersection>
<intersection>279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,271.5,534.5,271.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection>
<intersection>534.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,279.5,517,279.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>517 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>534.5,268,534.5,271.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>271.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569,272,569,279.5</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>272 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569,272,594,272</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>569 0</intersection>
<intersection>594 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>594,267.5,594,272</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>272 1</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>629,272,629,279.5</points>
<intersection>272 1</intersection>
<intersection>279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>629,272,649,272</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>629 0</intersection>
<intersection>649 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>626,279.5,629,279.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>629 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>649,267.5,649,272</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>272 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230,276.5,620,276.5</points>
<connection>
<GID>128</GID>
<name>clock</name></connection>
<connection>
<GID>126</GID>
<name>clock</name></connection>
<connection>
<GID>122</GID>
<name>clock</name></connection>
<connection>
<GID>120</GID>
<name>clock</name></connection>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<connection>
<GID>116</GID>
<name>clock</name></connection>
<connection>
<GID>114</GID>
<name>clock</name></connection>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<connection>
<GID>124</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,234,263,247.5</points>
<intersection>234 1</intersection>
<intersection>241 5</intersection>
<intersection>247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,234,286.5,234</points>
<intersection>263 0</intersection>
<intersection>286.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260.5,247.5,263,247.5</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>263 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>286.5,234,286.5,236.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>234 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>263,241,264.5,241</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>263 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,234,311,247.5</points>
<intersection>234 1</intersection>
<intersection>240 5</intersection>
<intersection>247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,234,328,234</points>
<intersection>311 0</intersection>
<intersection>328 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,247.5,311,247.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>311 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>328,234,328,236</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>234 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>311,240,313,240</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357.5,236,357.5,247.5</points>
<intersection>236 4</intersection>
<intersection>241 5</intersection>
<intersection>247.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>357.5,247.5,358,247.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>357.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>357.5,236,378.5,236</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>357.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>357.5,241,359.5,241</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>357.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,236,408.5,247.5</points>
<intersection>236 1</intersection>
<intersection>247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,236,427,236</points>
<intersection>408.5 0</intersection>
<intersection>409.5 4</intersection>
<intersection>427 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>407.5,247.5,408.5,247.5</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>427,236,427,237</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>236 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>409.5,236,409.5,241</points>
<intersection>236 1</intersection>
<intersection>241 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>409.5,241,414,241</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>409.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,241.5,457.5,247.5</points>
<intersection>241.5 5</intersection>
<intersection>247.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>455.5,247.5,457.5,247.5</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>457.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>457.5,241.5,474,241.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>457.5 0</intersection>
<intersection>474 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>474,237.5,474,241.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>241.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,239.5,516,247.5</points>
<intersection>239.5 1</intersection>
<intersection>247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,239.5,531.5,239.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection>
<intersection>531.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,247.5,516,247.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>516 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>531.5,236,531.5,239.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>239.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568,240,568,247.5</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>240 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>568,240,593,240</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>568 0</intersection>
<intersection>593 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>593,235.5,593,240</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>240 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>628,240,628,247.5</points>
<intersection>240 1</intersection>
<intersection>247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>628,240,648.5,240</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>628 0</intersection>
<intersection>648.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>625,247.5,628,247.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>628 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>648.5,235.5,648.5,240</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>240 1</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229,244,619,244</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>254.5 25</intersection>
<intersection>304 24</intersection>
<intersection>352 23</intersection>
<intersection>401.5 22</intersection>
<intersection>449.5 21</intersection>
<intersection>507 20</intersection>
<intersection>562 19</intersection>
<intersection>619 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>619,244,619,244.5</points>
<connection>
<GID>153</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>562,244,562,244.5</points>
<connection>
<GID>151</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>507,244,507,244.5</points>
<connection>
<GID>149</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>449.5,244,449.5,244.5</points>
<connection>
<GID>147</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>401.5,244,401.5,244.5</points>
<connection>
<GID>145</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>352,244,352,244.5</points>
<connection>
<GID>143</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>304,244,304,244.5</points>
<connection>
<GID>141</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>254.5,244,254.5,244.5</points>
<connection>
<GID>139</GID>
<name>clock</name></connection>
<intersection>244 1</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,207.5,262,220</points>
<intersection>207.5 1</intersection>
<intersection>213.5 5</intersection>
<intersection>220 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,207.5,286.5,207.5</points>
<intersection>262 0</intersection>
<intersection>286.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>260.5,220,262,220</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>262 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>286.5,207.5,286.5,209</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>207.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>262,213.5,264.5,213.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,206.5,311.5,220</points>
<intersection>206.5 1</intersection>
<intersection>212.5 5</intersection>
<intersection>220 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,206.5,328,206.5</points>
<intersection>311.5 0</intersection>
<intersection>328 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,220,311.5,220</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>311.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>328,206.5,328,208.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>206.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>311.5,212.5,313,212.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358,208.5,358,220</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<intersection>208.5 3</intersection>
<intersection>213.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>358,208.5,378.5,208.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>358,213.5,359.5,213.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>358 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,207,408.5,220</points>
<intersection>207 1</intersection>
<intersection>220 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408,207,427,207</points>
<intersection>408 4</intersection>
<intersection>408.5 0</intersection>
<intersection>427 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>407.5,220,408.5,220</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>427,207,427,209.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>207 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>408,207,408,214</points>
<intersection>207 1</intersection>
<intersection>214 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>408,214,409,214</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>408 4</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,214,457.5,220</points>
<intersection>214 5</intersection>
<intersection>220 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>455.5,220,457.5,220</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>457.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>457.5,214,474,214</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>457.5 0</intersection>
<intersection>474 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>474,210,474,214</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>214 5</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,212,516,220</points>
<intersection>212 1</intersection>
<intersection>220 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,212,534,212</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection>
<intersection>534 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,220,516,220</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>516 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>534,209,534,212</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>212 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568,212.5,568,220</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>212.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>568,212.5,593,212.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>568 0</intersection>
<intersection>593 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>593,208.5,593,212.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>212.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>628,212.5,628,220</points>
<intersection>212.5 1</intersection>
<intersection>220 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>628,212.5,651.5,212.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>628 0</intersection>
<intersection>651.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>625,220,628,220</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>628 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>651.5,211,651.5,212.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>212.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229,217,619,217</points>
<connection>
<GID>178</GID>
<name>clock</name></connection>
<connection>
<GID>176</GID>
<name>clock</name></connection>
<connection>
<GID>174</GID>
<name>clock</name></connection>
<connection>
<GID>172</GID>
<name>clock</name></connection>
<connection>
<GID>170</GID>
<name>clock</name></connection>
<connection>
<GID>168</GID>
<name>clock</name></connection>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<connection>
<GID>163</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,310,225,310</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,277.5,214,309</points>
<intersection>277.5 1</intersection>
<intersection>309 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,277.5,224,277.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,309,214,309</points>
<connection>
<GID>112</GID>
<name>OUT_2</name></connection>
<intersection>214 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,245,213.5,308</points>
<intersection>245 1</intersection>
<intersection>308 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,245,223,245</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,308,213.5,308</points>
<connection>
<GID>112</GID>
<name>OUT_1</name></connection>
<intersection>213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209.5,218,209.5,307</points>
<intersection>218 1</intersection>
<intersection>307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,218,223,218</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>209.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,307,209.5,307</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>209.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,193,219.5,216</points>
<intersection>193 1</intersection>
<intersection>216 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,193,219.5,193</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>219.5,216,223,216</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>219.5 0</intersection>
<intersection>221.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>221.5,216,221.5,243</points>
<intersection>216 2</intersection>
<intersection>243 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>218.5,243,223,243</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>218.5 6</intersection>
<intersection>221.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>218.5,243,218.5,275.5</points>
<intersection>243 4</intersection>
<intersection>275.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>218.5,275.5,224,275.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>218.5 6</intersection>
<intersection>220 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>220,275.5,220,308</points>
<intersection>275.5 7</intersection>
<intersection>308 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>220,308,225,308</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>220 8</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217.5,176.5,247.5,176.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<connection>
<GID>191</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,162.5,247,168</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>168 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>249.5,168,249.5,173.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>168 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>247,168,249.5,168</points>
<intersection>247 0</intersection>
<intersection>249.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299,162,299,167.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>167.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>298.5,167.5,298.5,173</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>167.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>298.5,167.5,299,167.5</points>
<intersection>298.5 1</intersection>
<intersection>299 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346,161.5,346,167</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>167 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>346.5,167,346.5,173</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>167 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>346,167,346.5,167</points>
<intersection>346 0</intersection>
<intersection>346.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,162,393.5,166</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<intersection>166 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>394,166,394,170.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>166 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>393.5,166,394,166</points>
<intersection>393.5 0</intersection>
<intersection>394 1</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,162.5,443,166.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>166.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>442.5,166.5,442.5,170.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>442.5,166.5,443,166.5</points>
<intersection>442.5 1</intersection>
<intersection>443 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498,162.5,498,167</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>167 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>497.5,167,497.5,172</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>167 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>497.5,167,498,167</points>
<intersection>497.5 1</intersection>
<intersection>498 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>554,162,554,166.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>166.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>553.5,166.5,553.5,171.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>553.5,166.5,554,166.5</points>
<intersection>553.5 1</intersection>
<intersection>554 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>615,162.5,615,166</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>166 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>615.5,166,615.5,170</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>166 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>615,166,615.5,166</points>
<intersection>615 0</intersection>
<intersection>615.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>615.5,175.5,615.5,312</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>220 4</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 2</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>615.5,312,621,312</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>615.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>615.5,279.5,620,279.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>615.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>615.5,247.5,619,247.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>615.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>615.5,220,619,220</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>615.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>553.5,177,553.5,312</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>220 4</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 2</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>553.5,312,564,312</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>553.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553.5,279.5,563,279.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>553.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>553.5,247.5,562,247.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>553.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>553.5,220,562,220</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>553.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497.5,177.5,497.5,312</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>220 5</intersection>
<intersection>247.5 4</intersection>
<intersection>279.5 1</intersection>
<intersection>312 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,279.5,508,279.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>497.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>497.5,312,509,312</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>497.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>497.5,247.5,507,247.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>497.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>497.5,220,507,220</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>497.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442.5,176,442.5,312</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>220 4</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 2</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,312,451.5,312</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>442.5,279.5,450.5,279.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>442.5,247.5,449.5,247.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>442.5,220,449.5,220</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,176,394,312</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>220 4</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 2</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>394,312,403.5,312</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>394 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>394,279.5,402.5,279.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>394 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>394,247.5,401.5,247.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>394 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>394,220,401.5,220</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>394 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346.5,178.5,346.5,312</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>220 4</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 2</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>346.5,312,354,312</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346.5,279.5,353,279.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>346.5,247.5,352,247.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>346.5,220,352,220</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,178.5,298.5,312</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 4</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>298.5,312,306,312</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298.5,220,304,220</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>298.5,247.5,304,247.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>298.5,279.5,305,279.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,179,249.5,312</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>220 2</intersection>
<intersection>247.5 3</intersection>
<intersection>279.5 4</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,312,256.5,312</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,220,254.5,220</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>249.5,247.5,254.5,247.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>249.5,279.5,255.5,279.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,212,277.5,212.5</points>
<intersection>212 1</intersection>
<intersection>212.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,212,284.5,212</points>
<connection>
<GID>187</GID>
<name>ENABLE_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270.5,212.5,277.5,212.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>277.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,239.5,277.5,240</points>
<intersection>239.5 1</intersection>
<intersection>240 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,239.5,284.5,239.5</points>
<connection>
<GID>162</GID>
<name>ENABLE_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>270.5,240,277.5,240</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<intersection>277.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,214,339.5,273.5</points>
<intersection>214 3</intersection>
<intersection>241.5 4</intersection>
<intersection>273.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>337.5,272.5,337.5,333.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>272.5 5</intersection>
<intersection>273.5 2</intersection>
<intersection>307 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,273.5,339.5,273.5</points>
<intersection>337.5 1</intersection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>328,214,339.5,214</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>328,241.5,339.5,241.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>332,272.5,337.5,272.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>337.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>331.5,307,337.5,307</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>337.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,271,279,272</points>
<intersection>271 1</intersection>
<intersection>272 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,271,284,271</points>
<connection>
<GID>136</GID>
<name>ENABLE_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>271.5,272,279,272</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,304,279.5,304.5</points>
<intersection>304 1</intersection>
<intersection>304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,304,283.5,304</points>
<connection>
<GID>99</GID>
<name>ENABLE_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>272.5,304.5,279.5,304.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,303.5,325,304.5</points>
<intersection>303.5 1</intersection>
<intersection>304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,303.5,325,303.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>325 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>325,304.5,329.5,304.5</points>
<connection>
<GID>98</GID>
<name>ENABLE_0</name></connection>
<intersection>325 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327,270,327,271</points>
<intersection>270 1</intersection>
<intersection>271 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327,270,330,270</points>
<connection>
<GID>137</GID>
<name>ENABLE_0</name></connection>
<intersection>327 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320,271,327,271</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>327 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>319,239,326,239</points>
<connection>
<GID>161</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>142</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>319,211.5,326,211.5</points>
<connection>
<GID>186</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>167</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,303.5,373,304.5</points>
<intersection>303.5 1</intersection>
<intersection>304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373,303.5,378.5,303.5</points>
<connection>
<GID>97</GID>
<name>ENABLE_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>367.5,304.5,373,304.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>373 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,271,372,272</points>
<intersection>271 1</intersection>
<intersection>272 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372,271,377.5,271</points>
<connection>
<GID>135</GID>
<name>ENABLE_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366.5,272,372,272</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>372 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>371,239,371,240</points>
<intersection>239 1</intersection>
<intersection>240 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>371,239,376.5,239</points>
<connection>
<GID>160</GID>
<name>ENABLE_0</name></connection>
<intersection>371 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>365.5,240,371,240</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>371 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>371,211.5,371,212.5</points>
<intersection>211.5 1</intersection>
<intersection>212.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>371,211.5,376.5,211.5</points>
<connection>
<GID>185</GID>
<name>ENABLE_0</name></connection>
<intersection>371 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>365.5,212.5,371,212.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>371 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422,304.5,422,305</points>
<intersection>304.5 1</intersection>
<intersection>305 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>422,304.5,427,304.5</points>
<connection>
<GID>94</GID>
<name>ENABLE_0</name></connection>
<intersection>422 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>417,305,422,305</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>422 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,214.5,291,274.5</points>
<intersection>214.5 3</intersection>
<intersection>242 4</intersection>
<intersection>274.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>290.5,273.5,290.5,335</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>273.5 5</intersection>
<intersection>274.5 2</intersection>
<intersection>306.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,274.5,291,274.5</points>
<intersection>290.5 1</intersection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286.5,214.5,291,214.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>286.5,242,291,242</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>286,273.5,290.5,273.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>290.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285.5,306.5,290.5,306.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>290.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421,272,421,272.5</points>
<intersection>272 1</intersection>
<intersection>272.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>421,272,426,272</points>
<connection>
<GID>134</GID>
<name>ENABLE_0</name></connection>
<intersection>421 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>416,272.5,421,272.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>421 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>420,240,425,240</points>
<connection>
<GID>159</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>146</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420,212.5,420,213</points>
<intersection>212.5 1</intersection>
<intersection>213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420,212.5,425,212.5</points>
<connection>
<GID>184</GID>
<name>ENABLE_0</name></connection>
<intersection>420 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>415,213,420,213</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>420 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>466,305,474,305</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469,272.5,469,273</points>
<intersection>272.5 1</intersection>
<intersection>273 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>469,272.5,473,272.5</points>
<connection>
<GID>130</GID>
<name>ENABLE_0</name></connection>
<intersection>469 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>465,273,469,273</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>469 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>464,240.5,472,240.5</points>
<connection>
<GID>155</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>148</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>464,213,472,213</points>
<connection>
<GID>180</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>173</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>527,211,527,212</points>
<intersection>211 1</intersection>
<intersection>212 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>522.5,211,527,211</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>527 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527,212,532,212</points>
<connection>
<GID>181</GID>
<name>ENABLE_0</name></connection>
<intersection>527 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>527,238.5,527,239</points>
<intersection>238.5 1</intersection>
<intersection>239 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>522.5,238.5,527,238.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>527 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527,239,529.5,239</points>
<connection>
<GID>156</GID>
<name>ENABLE_0</name></connection>
<intersection>527 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>528,270.5,528,271</points>
<intersection>270.5 2</intersection>
<intersection>271 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>528,271,532.5,271</points>
<connection>
<GID>131</GID>
<name>ENABLE_0</name></connection>
<intersection>528 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>523.5,270.5,528,270.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>528 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524.5,303,534,303</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<connection>
<GID>91</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,303.5,584.5,304</points>
<intersection>303.5 1</intersection>
<intersection>304 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>576.5,303.5,584.5,303.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,304,593,304</points>
<connection>
<GID>92</GID>
<name>ENABLE_0</name></connection>
<intersection>584.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,270.5,583.5,271</points>
<intersection>270.5 1</intersection>
<intersection>271 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,270.5,592,270.5</points>
<connection>
<GID>132</GID>
<name>ENABLE_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>575.5,271,583.5,271</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>583.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>582.5,238.5,582.5,239</points>
<intersection>238.5 2</intersection>
<intersection>239 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>574.5,239,582.5,239</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>582.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,238.5,591,238.5</points>
<connection>
<GID>157</GID>
<name>ENABLE_0</name></connection>
<intersection>582.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,211.5,591,211.5</points>
<connection>
<GID>182</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>177</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641,211.5,641,214</points>
<intersection>211.5 2</intersection>
<intersection>214 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641,214,649.5,214</points>
<connection>
<GID>183</GID>
<name>ENABLE_0</name></connection>
<intersection>641 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>634.5,211.5,641,211.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>641 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,238.5,640,239</points>
<intersection>238.5 1</intersection>
<intersection>239 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,238.5,646.5,238.5</points>
<connection>
<GID>158</GID>
<name>ENABLE_0</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>634.5,239,640,239</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641,270.5,641,271</points>
<intersection>270.5 1</intersection>
<intersection>271 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641,270.5,647,270.5</points>
<connection>
<GID>133</GID>
<name>ENABLE_0</name></connection>
<intersection>641 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>635.5,271,641,271</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>641 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>636.5,303.5,648.5,303.5</points>
<connection>
<GID>93</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>655.5,316,655.5,326.5</points>
<intersection>316 2</intersection>
<intersection>326.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>650.5,216.5,650.5,316</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>216.5 4</intersection>
<intersection>241 6</intersection>
<intersection>273 5</intersection>
<intersection>316 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>650.5,316,655.5,316</points>
<intersection>650.5 1</intersection>
<intersection>655.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>654.5,326.5,655.5,326.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>655.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>650.5,216.5,651.5,216.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>650.5 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>649,273,650.5,273</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>650.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>648.5,241,650.5,241</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>650.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,214,603,271</points>
<intersection>214 3</intersection>
<intersection>241 4</intersection>
<intersection>271 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>598.5,271,598.5,328.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>271 2</intersection>
<intersection>273 5</intersection>
<intersection>306.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>598.5,271,603,271</points>
<intersection>598.5 1</intersection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>593,214,603,214</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>593,241,603,241</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>594,273,598.5,273</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>598.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>595,306.5,598.5,306.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>598.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,214.5,540,273.5</points>
<intersection>214.5 3</intersection>
<intersection>241.5 4</intersection>
<intersection>273.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>541,273.5,541,333</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>273.5 2</intersection>
<intersection>305.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>534.5,273.5,541,273.5</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>540 0</intersection>
<intersection>541 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>534,214.5,540,214.5</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>540 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>531.5,241.5,540,241.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>540 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>536,305.5,541,305.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>541 1</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>481,215.5,481,275</points>
<intersection>215.5 3</intersection>
<intersection>243 4</intersection>
<intersection>275 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>482,275,482,334.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>275 2</intersection>
<intersection>307.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>475,275,482,275</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>481 0</intersection>
<intersection>482 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>474,215.5,481,215.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>481 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>474,243,481,243</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>481 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>476,307.5,482,307.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>482 1</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-3.20813e-005,719.901,1224,114.901</PageViewport></page 4>
<page 5>
<PageViewport>-3.20813e-005,719.901,1224,114.901</PageViewport></page 5>
<page 6>
<PageViewport>-3.20813e-005,719.901,1224,114.901</PageViewport></page 6>
<page 7>
<PageViewport>-3.20813e-005,719.901,1224,114.901</PageViewport></page 7>
<page 8>
<PageViewport>-3.20813e-005,719.901,1224,114.901</PageViewport></page 8>
<page 9>
<PageViewport>-3.20813e-005,719.901,1224,114.901</PageViewport></page 9></circuit>