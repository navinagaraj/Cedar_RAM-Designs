<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-62.8331,131.756,759.607,-274.76</PageViewport></page 0>
<page 1>
<PageViewport>12.4661,27.3892,359.434,-144.11</PageViewport>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>93,-14.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>100.5,-14.5</position>
<gparam>LABEL_TEXT X2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>BA_TRI_STATE</type>
<position>93,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>BA_TRI_STATE</type>
<position>100.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_FULLADDER_1BIT</type>
<position>111,-36</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_B_0</ID>100 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>carry_in</ID>115 </input>
<output>
<ID>carry_out</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>GA_LED</type>
<position>111,-43</position>
<input>
<ID>N_in3</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_TOGGLE</type>
<position>107.5,-18</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_TOGGLE</type>
<position>115,-18</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>107.5,-14.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_LABEL</type>
<position>115,-14.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>BA_TRI_STATE</type>
<position>107.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>204</ID>
<type>BA_TRI_STATE</type>
<position>115,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_FULLADDER_1BIT</type>
<position>124.5,-36</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_B_0</ID>105 </input>
<output>
<ID>OUT_0</ID>101 </output>
<output>
<ID>carry_out</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>206</ID>
<type>GA_LED</type>
<position>124.5,-43</position>
<input>
<ID>N_in3</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>121,-18</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_TOGGLE</type>
<position>128.5,-18</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>121,-14.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>128.5,-14.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>BA_TRI_STATE</type>
<position>121,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>212</ID>
<type>BA_TRI_STATE</type>
<position>128.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>133,-49</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>220</ID>
<type>GA_LED</type>
<position>19,-50.5</position>
<input>
<ID>N_in3</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>82,0.5</position>
<gparam>LABEL_TEXT X Input Data</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>133,-51.5</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>18.5,-53</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_LABEL</type>
<position>110,0.5</position>
<gparam>LABEL_TEXT 8-bit Data = 10101011</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>110,-3.5</position>
<gparam>LABEL_TEXT 8-bit Data = 11010101</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>73.5,-47.5</position>
<gparam>LABEL_TEXT SUM   = 10000000</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>82,-3.5</position>
<gparam>LABEL_TEXT Y Input Data</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>19.5,-57</position>
<gparam>LABEL_TEXT Carry = 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_FULLADDER_1BIT</type>
<position>25,-36</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_B_0</ID>70 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>carry_in</ID>109 </input>
<output>
<ID>carry_out</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>25,-43</position>
<input>
<ID>N_in3</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>21.5,-18</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>29,-18</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>21.5,-14.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>29,-14.5</position>
<gparam>LABEL_TEXT X7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>BA_TRI_STATE</type>
<position>21.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>BA_TRI_STATE</type>
<position>29,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_FULLADDER_1BIT</type>
<position>40,-36</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_B_0</ID>75 </input>
<output>
<ID>OUT_0</ID>71 </output>
<input>
<ID>carry_in</ID>110 </input>
<output>
<ID>carry_out</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>40,-43</position>
<input>
<ID>N_in3</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>36.5,-18</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_TOGGLE</type>
<position>44,-18</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>36.5,-14.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>44,-14.5</position>
<gparam>LABEL_TEXT X6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>BA_TRI_STATE</type>
<position>36.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>BA_TRI_STATE</type>
<position>44,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_FULLADDER_1BIT</type>
<position>54.5,-36</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_B_0</ID>80 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>carry_in</ID>111 </input>
<output>
<ID>carry_out</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>GA_LED</type>
<position>54.5,-43</position>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>51,-18</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>58.5,-18</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>51,-14.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>58.5,-14.5</position>
<gparam>LABEL_TEXT X5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>BA_TRI_STATE</type>
<position>51,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>172</ID>
<type>BA_TRI_STATE</type>
<position>58.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_FULLADDER_1BIT</type>
<position>68,-36</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_B_0</ID>85 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>carry_in</ID>112 </input>
<output>
<ID>carry_out</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>68,-43</position>
<input>
<ID>N_in3</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_TOGGLE</type>
<position>64.5,-18</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_TOGGLE</type>
<position>72,-18</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>64.5,-14.5</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>72,-14.5</position>
<gparam>LABEL_TEXT X4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>BA_TRI_STATE</type>
<position>64.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>BA_TRI_STATE</type>
<position>72,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_FULLADDER_1BIT</type>
<position>81.5,-36</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_B_0</ID>90 </input>
<output>
<ID>OUT_0</ID>86 </output>
<input>
<ID>carry_in</ID>113 </input>
<output>
<ID>carry_out</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>81.5,-43</position>
<input>
<ID>N_in3</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>78,-18</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_TOGGLE</type>
<position>85.5,-18</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>78,-14.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>85.5,-14.5</position>
<gparam>LABEL_TEXT X3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>BA_TRI_STATE</type>
<position>78,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>188</ID>
<type>BA_TRI_STATE</type>
<position>85.5,-29</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_FULLADDER_1BIT</type>
<position>96.5,-36</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_B_0</ID>95 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>carry_in</ID>114 </input>
<output>
<ID>carry_out</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>190</ID>
<type>GA_LED</type>
<position>96.5,-43</position>
<input>
<ID>N_in3</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>93,-18</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>100.5,-18</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-42,25,-39</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>96</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-26,21.5,-20</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-26,29,-20</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-33,26,-32</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,-32,29,-31.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26,-32,29,-32</points>
<intersection>26 0</intersection>
<intersection>29 1</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-33,24,-32</points>
<connection>
<GID>79</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>21.5,-32,21.5,-31.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-32,24,-32</points>
<intersection>21.5 1</intersection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-42,40,-39</points>
<connection>
<GID>158</GID>
<name>N_in3</name></connection>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-26,36.5,-20</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-26,44,-20</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-33,41,-32</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44,-32,44,-31.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41,-32,44,-32</points>
<intersection>41 0</intersection>
<intersection>44 1</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-33,39,-32</points>
<connection>
<GID>157</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>36.5,-32,36.5,-31.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-32,39,-32</points>
<intersection>36.5 1</intersection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-42,54.5,-39</points>
<connection>
<GID>166</GID>
<name>N_in3</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-26,51,-20</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-26,58.5,-20</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-33,55.5,-32</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58.5,-32,58.5,-31.5</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-32,58.5,-32</points>
<intersection>55.5 0</intersection>
<intersection>58.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-33,53.5,-32</points>
<connection>
<GID>165</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51,-32,51,-31.5</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51,-32,53.5,-32</points>
<intersection>51 1</intersection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-42,68,-39</points>
<connection>
<GID>174</GID>
<name>N_in3</name></connection>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-26,64.5,-20</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-26,72,-20</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-33,69,-32</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72,-32,72,-31.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-32,72,-32</points>
<intersection>69 0</intersection>
<intersection>72 1</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-33,67,-32</points>
<connection>
<GID>173</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-32,64.5,-31.5</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-32,67,-32</points>
<intersection>64.5 1</intersection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-42,81.5,-39</points>
<connection>
<GID>182</GID>
<name>N_in3</name></connection>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-26,78,-20</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-26,85.5,-20</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-33,82.5,-32</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>85.5,-32,85.5,-31.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-32,85.5,-32</points>
<intersection>82.5 0</intersection>
<intersection>85.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-33,80.5,-32</points>
<connection>
<GID>181</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78,-32,78,-31.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-32,80.5,-32</points>
<intersection>78 1</intersection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-42,96.5,-39</points>
<connection>
<GID>190</GID>
<name>N_in3</name></connection>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-26,93,-20</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-26,100.5,-20</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<connection>
<GID>196</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-33,97.5,-32</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>100.5,-32,100.5,-31.5</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-32,100.5,-32</points>
<intersection>97.5 0</intersection>
<intersection>100.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-33,95.5,-32</points>
<connection>
<GID>189</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93,-32,93,-31.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>93,-32,95.5,-32</points>
<intersection>93 1</intersection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-42,111,-39</points>
<connection>
<GID>198</GID>
<name>N_in3</name></connection>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-26,107.5,-20</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-26,115,-20</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-33,112,-32</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>115,-32,115,-31.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112,-32,115,-32</points>
<intersection>112 0</intersection>
<intersection>115 1</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-33,110,-32</points>
<connection>
<GID>197</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>107.5,-32,107.5,-31.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-32,110,-32</points>
<intersection>107.5 1</intersection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-42,124.5,-39</points>
<connection>
<GID>206</GID>
<name>N_in3</name></connection>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-26,121,-20</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-26,128.5,-20</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-33,125.5,-32</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>128.5,-32,128.5,-31.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-32,128.5,-32</points>
<intersection>125.5 0</intersection>
<intersection>128.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-33,123.5,-32</points>
<connection>
<GID>205</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>121,-32,121,-31.5</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121,-32,123.5,-32</points>
<intersection>121 1</intersection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-29,133,-29</points>
<connection>
<GID>154</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>156</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>163</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>164</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>171</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>172</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>179</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>180</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>187</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>188</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>195</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>196</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>203</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>204</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>211</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>212</GID>
<name>ENABLE_0</name></connection>
<intersection>133 66</intersection></hsegment>
<vsegment>
<ID>66</ID>
<points>133,-47,133,-29</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-49.5,19,-36</points>
<connection>
<GID>220</GID>
<name>N_in3</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-36,21,-36</points>
<connection>
<GID>79</GID>
<name>carry_out</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-36,36,-36</points>
<connection>
<GID>79</GID>
<name>carry_in</name></connection>
<connection>
<GID>157</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-36,50.5,-36</points>
<connection>
<GID>157</GID>
<name>carry_in</name></connection>
<connection>
<GID>165</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-36,64,-36</points>
<connection>
<GID>165</GID>
<name>carry_in</name></connection>
<connection>
<GID>173</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-36,77.5,-36</points>
<connection>
<GID>173</GID>
<name>carry_in</name></connection>
<connection>
<GID>181</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-36,92.5,-36</points>
<connection>
<GID>181</GID>
<name>carry_in</name></connection>
<connection>
<GID>189</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-36,107,-36</points>
<connection>
<GID>189</GID>
<name>carry_in</name></connection>
<connection>
<GID>197</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-36,120.5,-36</points>
<connection>
<GID>197</GID>
<name>carry_in</name></connection>
<connection>
<GID>205</GID>
<name>carry_out</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>168.606,161.6,991.045,-244.916</PageViewport></page 2>
<page 3>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 3>
<page 4>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 4>
<page 5>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 5>
<page 6>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 6>
<page 7>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 7>
<page 8>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 8>
<page 9>
<PageViewport>-3.20813e-005,384.093,1224,-220.907</PageViewport></page 9></circuit>