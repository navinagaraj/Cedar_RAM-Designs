<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-506.495,205.616,254.216,-170.389</PageViewport>
<gate>
<ID>778</ID>
<type>AA_AND2</type>
<position>-162,-1</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>779</ID>
<type>AA_AND2</type>
<position>-170.5,-12</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>780</ID>
<type>AA_AND2</type>
<position>-162.5,-17</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>-368,-23.5</position>
<gparam>LABEL_TEXT now we got every bytes cleared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>781</ID>
<type>AA_AND2</type>
<position>-170.5,-27</position>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>782</ID>
<type>AA_AND2</type>
<position>-162,-32</position>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>-369.5,-30</position>
<gparam>LABEL_TEXT we can write data to registers</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>783</ID>
<type>AA_AND2</type>
<position>-170.5,-42.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AA_AND2</type>
<position>-162,-47.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>521 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-276.5,24.5</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>786</ID>
<type>BE_DECODER_3x8</type>
<position>-243.5,20</position>
<input>
<ID>ENABLE</ID>625 </input>
<input>
<ID>IN_0</ID>629 </input>
<input>
<ID>IN_1</ID>628 </input>
<input>
<ID>IN_2</ID>626 </input>
<output>
<ID>OUT_0</ID>482 </output>
<output>
<ID>OUT_1</ID>481 </output>
<output>
<ID>OUT_2</ID>480 </output>
<output>
<ID>OUT_3</ID>479 </output>
<output>
<ID>OUT_4</ID>478 </output>
<output>
<ID>OUT_5</ID>477 </output>
<output>
<ID>OUT_6</ID>476 </output>
<output>
<ID>OUT_7</ID>475 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-360,-37</position>
<gparam>LABEL_TEXT always on to make decoder on</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>788</ID>
<type>AA_TOGGLE</type>
<position>-263.5,19</position>
<output>
<ID>OUT_0</ID>626 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-274,19</position>
<gparam>LABEL_TEXT i1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-274,14.5</position>
<gparam>LABEL_TEXT i2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>790</ID>
<type>AA_TOGGLE</type>
<position>-263.5,14.5</position>
<output>
<ID>OUT_0</ID>628 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>-274,10</position>
<gparam>LABEL_TEXT i3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>792</ID>
<type>AA_TOGGLE</type>
<position>-263.5,11.5</position>
<output>
<ID>OUT_0</ID>629 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-269.5,5.5</position>
<gparam>LABEL_TEXT input combitaions that is address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>794</ID>
<type>AA_TOGGLE</type>
<position>-272,23.5</position>
<output>
<ID>OUT_0</ID>625 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-285.5,-6</position>
<gparam>LABEL_TEXT fst comb 000</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>795</ID>
<type>BA_TRI_STATE</type>
<position>-143,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>483 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>796</ID>
<type>BA_TRI_STATE</type>
<position>-119.5,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>484 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-246.5,-35.5</position>
<gparam>LABEL_TEXT selected register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>797</ID>
<type>BA_TRI_STATE</type>
<position>-97,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>485 </input>
<output>
<ID>OUT_0</ID>531 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>798</ID>
<type>BA_TRI_STATE</type>
<position>-76.5,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>486 </input>
<output>
<ID>OUT_0</ID>533 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>-260.5,-6</position>
<gparam>LABEL_TEXT 00001111</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>799</ID>
<type>BA_TRI_STATE</type>
<position>-55,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>487 </input>
<output>
<ID>OUT_0</ID>535 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>800</ID>
<type>BA_TRI_STATE</type>
<position>-33.5,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>537 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>-289.5,0.5</position>
<gparam>LABEL_TEXT i/p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>801</ID>
<type>BA_TRI_STATE</type>
<position>-12,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>489 </input>
<output>
<ID>OUT_0</ID>539 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>802</ID>
<type>BA_TRI_STATE</type>
<position>8,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>490 </input>
<output>
<ID>OUT_0</ID>541 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>-261,-0.5</position>
<gparam>LABEL_TEXT DATA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>803</ID>
<type>BA_TRI_STATE</type>
<position>-123.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>492 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>804</ID>
<type>BA_TRI_STATE</type>
<position>-100,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>530 </input>
<output>
<ID>OUT_0</ID>493 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>-372,4.5</position>
<gparam>LABEL_TEXT WRITE using clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>805</ID>
<type>BA_TRI_STATE</type>
<position>-78.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>532 </input>
<output>
<ID>OUT_0</ID>494 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>-286,-12</position>
<gparam>LABEL_TEXT sec combo 011</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>806</ID>
<type>BA_TRI_STATE</type>
<position>-57.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>534 </input>
<output>
<ID>OUT_0</ID>495 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-260.5,-12.5</position>
<gparam>LABEL_TEXT 11110000</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>807</ID>
<type>BA_TRI_STATE</type>
<position>-36,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>536 </input>
<output>
<ID>OUT_0</ID>496 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>-286,-18.5</position>
<gparam>LABEL_TEXT third combo 111</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>808</ID>
<type>BA_TRI_STATE</type>
<position>-14.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>538 </input>
<output>
<ID>OUT_0</ID>497 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-261,-19</position>
<gparam>LABEL_TEXT 00111100</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>809</ID>
<type>BA_TRI_STATE</type>
<position>6,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>540 </input>
<output>
<ID>OUT_0</ID>498 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>810</ID>
<type>BA_TRI_STATE</type>
<position>30.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>542 </input>
<output>
<ID>OUT_0</ID>499 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>-275,47</position>
<gparam>LABEL_TEXT now we read wat data we gave</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>812</ID>
<type>DA_FROM</type>
<position>-143,-73</position>
<input>
<ID>IN_0</ID>483 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>-371,35.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>814</ID>
<type>DA_FROM</type>
<position>-119.5,-73</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>-361.5,35.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>-384.5,36.5</position>
<gparam>LABEL_TEXT without delay</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>823</ID>
<type>DA_FROM</type>
<position>-97,-72</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>824</ID>
<type>DA_FROM</type>
<position>-76.5,-73</position>
<input>
<ID>IN_0</ID>486 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>825</ID>
<type>DA_FROM</type>
<position>-55,-72.5</position>
<input>
<ID>IN_0</ID>487 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>826</ID>
<type>DA_FROM</type>
<position>-33.5,-73</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>827</ID>
<type>DA_FROM</type>
<position>-12,-72.5</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>828</ID>
<type>DA_FROM</type>
<position>8,-71.5</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>829</ID>
<type>DA_FROM</type>
<position>-160.5,-64</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>831</ID>
<type>DA_FROM</type>
<position>-145,93</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>-184,92.5</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>835</ID>
<type>DE_TO</type>
<position>-126,107.5</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>836</ID>
<type>DE_TO</type>
<position>-103,107.5</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>837</ID>
<type>DE_TO</type>
<position>-80,107.5</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>838</ID>
<type>DE_TO</type>
<position>-59.5,108</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>839</ID>
<type>DE_TO</type>
<position>-38,108</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>840</ID>
<type>DE_TO</type>
<position>-16.5,108.5</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>841</ID>
<type>DE_TO</type>
<position>5,108</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>842</ID>
<type>DE_TO</type>
<position>25,107.5</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>844</ID>
<type>DA_FROM</type>
<position>-187,-65.5</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>846</ID>
<type>AA_TOGGLE</type>
<position>-370,29</position>
<output>
<ID>OUT_0</ID>606 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>847</ID>
<type>AA_TOGGLE</type>
<position>-370,21.5</position>
<output>
<ID>OUT_0</ID>607 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>848</ID>
<type>AA_TOGGLE</type>
<position>-370,14.5</position>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>849</ID>
<type>AA_TOGGLE</type>
<position>-352,-3.5</position>
<output>
<ID>OUT_0</ID>609 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>850</ID>
<type>AA_TOGGLE</type>
<position>-344,-3.5</position>
<output>
<ID>OUT_0</ID>610 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>851</ID>
<type>AA_TOGGLE</type>
<position>-337,-3</position>
<output>
<ID>OUT_0</ID>611 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>852</ID>
<type>AA_TOGGLE</type>
<position>-331,-2.5</position>
<output>
<ID>OUT_0</ID>612 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>853</ID>
<type>AA_TOGGLE</type>
<position>-325,-3.5</position>
<output>
<ID>OUT_0</ID>613 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>854</ID>
<type>AA_TOGGLE</type>
<position>-319,-3.5</position>
<output>
<ID>OUT_0</ID>614 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>855</ID>
<type>AA_TOGGLE</type>
<position>-313,-3</position>
<output>
<ID>OUT_0</ID>615 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>856</ID>
<type>AA_TOGGLE</type>
<position>-306,-3</position>
<output>
<ID>OUT_0</ID>616 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>858</ID>
<type>GA_LED</type>
<position>-355,43</position>
<input>
<ID>N_in3</ID>617 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>861</ID>
<type>GA_LED</type>
<position>-346.5,43</position>
<input>
<ID>N_in3</ID>618 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>862</ID>
<type>GA_LED</type>
<position>-339,43</position>
<input>
<ID>N_in3</ID>619 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>863</ID>
<type>GA_LED</type>
<position>-333,43</position>
<input>
<ID>N_in3</ID>620 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>864</ID>
<type>GA_LED</type>
<position>-326.5,43</position>
<input>
<ID>N_in3</ID>621 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>865</ID>
<type>GA_LED</type>
<position>-320.5,43</position>
<input>
<ID>N_in3</ID>622 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>866</ID>
<type>GA_LED</type>
<position>-313.5,43</position>
<input>
<ID>N_in3</ID>623 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>867</ID>
<type>GA_LED</type>
<position>-308,43</position>
<input>
<ID>N_in3</ID>624 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>869</ID>
<type>DE_TO</type>
<position>-363,29</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>871</ID>
<type>DE_TO</type>
<position>-362,21.5</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>872</ID>
<type>DE_TO</type>
<position>-362,14.5</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>873</ID>
<type>DE_TO</type>
<position>-352,6</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>874</ID>
<type>DE_TO</type>
<position>-344,6</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>875</ID>
<type>DE_TO</type>
<position>-337,6</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>876</ID>
<type>DE_TO</type>
<position>-331,6</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>877</ID>
<type>DE_TO</type>
<position>-325,6.5</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>878</ID>
<type>DE_TO</type>
<position>-319,6</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>879</ID>
<type>DE_TO</type>
<position>-313,6</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>880</ID>
<type>DE_TO</type>
<position>-306,6</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>882</ID>
<type>DA_FROM</type>
<position>-355,54</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>883</ID>
<type>DA_FROM</type>
<position>-346.5,53.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>884</ID>
<type>DA_FROM</type>
<position>-339,53.5</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>885</ID>
<type>DA_FROM</type>
<position>-333,54</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>886</ID>
<type>DA_FROM</type>
<position>-326.5,54</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>887</ID>
<type>DA_FROM</type>
<position>-320.5,54</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>888</ID>
<type>DA_FROM</type>
<position>-313.5,54</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>889</ID>
<type>DA_FROM</type>
<position>-308,54</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>895</ID>
<type>AA_LABEL</type>
<position>-357,67</position>
<gparam>LABEL_TEXT OUTPUT READ HERE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>638</ID>
<type>AE_DFF_LOW</type>
<position>-136,69</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>578 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>639</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,69</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>573 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>640</ID>
<type>AE_DFF_LOW</type>
<position>-90,69</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>572 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_DFF_LOW</type>
<position>-71,69</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>563 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>642</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,69</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>562 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>643</ID>
<type>AE_DFF_LOW</type>
<position>-27,69</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>553 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>644</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,69</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>545 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_DFF_LOW</type>
<position>14.5,69</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>543 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>647</ID>
<type>BA_TRI_STATE</type>
<position>-129,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>578 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>648</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>573 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>649</ID>
<type>BA_TRI_STATE</type>
<position>-83,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>572 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>650</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>563 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>651</ID>
<type>BA_TRI_STATE</type>
<position>-41,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>562 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>652</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>553 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>653</ID>
<type>BA_TRI_STATE</type>
<position>2,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>545 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>654</ID>
<type>BA_TRI_STATE</type>
<position>22,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>543 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>655</ID>
<type>AE_DFF_LOW</type>
<position>-136,53.5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>579 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>656</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,53.5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>574 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>657</ID>
<type>AE_DFF_LOW</type>
<position>-90,53.5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>571 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>658</ID>
<type>AE_DFF_LOW</type>
<position>-71,53.5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>564 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>659</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,53.5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>561 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>660</ID>
<type>AE_DFF_LOW</type>
<position>-27,53.5</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>554 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>661</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,53.5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>546 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>662</ID>
<type>AE_DFF_LOW</type>
<position>14.5,53.5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>544 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>663</ID>
<type>BA_TRI_STATE</type>
<position>-129,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>579 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>664</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>574 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>665</ID>
<type>BA_TRI_STATE</type>
<position>-83,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>571 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>666</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>564 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>667</ID>
<type>BA_TRI_STATE</type>
<position>-41,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>668</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>554 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>669</ID>
<type>BA_TRI_STATE</type>
<position>2,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>546 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>670</ID>
<type>BA_TRI_STATE</type>
<position>22,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>544 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>671</ID>
<type>AE_DFF_LOW</type>
<position>-136,37</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>582 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>672</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,37</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>575 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>673</ID>
<type>AE_DFF_LOW</type>
<position>-90,37</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>570 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>674</ID>
<type>AE_DFF_LOW</type>
<position>-71,37</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>565 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>675</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,37</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>560 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>676</ID>
<type>AE_DFF_LOW</type>
<position>-27,37</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>555 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>677</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,37</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>550 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>678</ID>
<type>AE_DFF_LOW</type>
<position>14.5,37</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>549 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>679</ID>
<type>BA_TRI_STATE</type>
<position>-129,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>582 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>680</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>575 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>681</ID>
<type>BA_TRI_STATE</type>
<position>-83,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>570 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>682</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>565 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>683</ID>
<type>BA_TRI_STATE</type>
<position>-41,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>560 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>684</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>555 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>685</ID>
<type>BA_TRI_STATE</type>
<position>2,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>550 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>686</ID>
<type>BA_TRI_STATE</type>
<position>22,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>549 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_DFF_LOW</type>
<position>-136,21</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>581 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>688</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,21</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>576 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>689</ID>
<type>AE_DFF_LOW</type>
<position>-90,21</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>569 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_DFF_LOW</type>
<position>-71,21</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>566 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>691</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,21</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>559 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_DFF_LOW</type>
<position>-27,21</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>556 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>693</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,21</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>551 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>694</ID>
<type>AE_DFF_LOW</type>
<position>14.5,21</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>548 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>695</ID>
<type>BA_TRI_STATE</type>
<position>-129,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>581 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>696</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>576 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>697</ID>
<type>BA_TRI_STATE</type>
<position>-83,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>569 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>698</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>566 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>699</ID>
<type>BA_TRI_STATE</type>
<position>-41,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>559 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>700</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>556 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>701</ID>
<type>BA_TRI_STATE</type>
<position>2,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>551 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>702</ID>
<type>BA_TRI_STATE</type>
<position>22,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>548 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>703</ID>
<type>AE_DFF_LOW</type>
<position>-136,5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>580 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>704</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>577 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>705</ID>
<type>AE_DFF_LOW</type>
<position>-90,5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>568 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>706</ID>
<type>AE_DFF_LOW</type>
<position>-71,5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>567 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>707</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>558 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>708</ID>
<type>AE_DFF_LOW</type>
<position>-27,5</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>557 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>709</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>552 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>710</ID>
<type>AE_DFF_LOW</type>
<position>14.5,5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>547 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>711</ID>
<type>BA_TRI_STATE</type>
<position>-129,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>580 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>712</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>577 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>713</ID>
<type>BA_TRI_STATE</type>
<position>-83,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>568 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>714</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>567 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>715</ID>
<type>BA_TRI_STATE</type>
<position>-41,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>558 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>716</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>557 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>717</ID>
<type>BA_TRI_STATE</type>
<position>2,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>552 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>718</ID>
<type>BA_TRI_STATE</type>
<position>22,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>547 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>719</ID>
<type>AE_DFF_LOW</type>
<position>-136,-11</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>583 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>720</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,-11</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>586 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>721</ID>
<type>AE_DFF_LOW</type>
<position>-90,-11</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>587 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>722</ID>
<type>AE_DFF_LOW</type>
<position>-71,-11</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>591 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>723</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,-11</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>596 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>724</ID>
<type>AE_DFF_LOW</type>
<position>-27,-11</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>597 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>725</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,-11</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>601 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>726</ID>
<type>AE_DFF_LOW</type>
<position>14.5,-11</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>603 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>727</ID>
<type>BA_TRI_STATE</type>
<position>-129,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>583 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>728</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>586 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>729</ID>
<type>BA_TRI_STATE</type>
<position>-83,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>587 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>730</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>591 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>731</ID>
<type>BA_TRI_STATE</type>
<position>-41,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>596 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>732</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>597 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>733</ID>
<type>BA_TRI_STATE</type>
<position>2,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>601 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>734</ID>
<type>BA_TRI_STATE</type>
<position>22,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>735</ID>
<type>AE_DFF_LOW</type>
<position>-136,-26</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>523 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>736</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,-26</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>585 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>737</ID>
<type>AE_DFF_LOW</type>
<position>-90,-26</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>590 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>738</ID>
<type>AE_DFF_LOW</type>
<position>-71,-26</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>593 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>739</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,-26</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>594 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>740</ID>
<type>AE_DFF_LOW</type>
<position>-27,-26</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>598 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>741</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,-26</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>600 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>742</ID>
<type>AE_DFF_LOW</type>
<position>14.5,-26</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>604 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>743</ID>
<type>BA_TRI_STATE</type>
<position>-129,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>523 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>744</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>585 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>745</ID>
<type>BA_TRI_STATE</type>
<position>-83,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>590 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>746</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>593 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>747</ID>
<type>BA_TRI_STATE</type>
<position>-41,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>594 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>748</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>598 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>749</ID>
<type>BA_TRI_STATE</type>
<position>2,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>600 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>750</ID>
<type>BA_TRI_STATE</type>
<position>22,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>604 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_DFF_LOW</type>
<position>-136,-41.5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>524 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>752</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,-41.5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>584 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>753</ID>
<type>AE_DFF_LOW</type>
<position>-90,-41.5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>589 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>754</ID>
<type>AE_DFF_LOW</type>
<position>-71,-41.5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>592 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>755</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,-41.5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>595 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>756</ID>
<type>AE_DFF_LOW</type>
<position>-27,-41.5</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>599 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>757</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,-41.5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>602 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>758</ID>
<type>AE_DFF_LOW</type>
<position>14.5,-41.5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>605 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>759</ID>
<type>BA_TRI_STATE</type>
<position>-129,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>760</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>584 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>761</ID>
<type>BA_TRI_STATE</type>
<position>-83,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>589 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>762</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>592 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>763</ID>
<type>BA_TRI_STATE</type>
<position>-41,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>595 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>764</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>599 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>765</ID>
<type>BA_TRI_STATE</type>
<position>2,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>602 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>766</ID>
<type>BA_TRI_STATE</type>
<position>22,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>605 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>768</ID>
<type>AA_AND2</type>
<position>-170.5,68</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>503 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>770</ID>
<type>AA_AND2</type>
<position>-162,63</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>771</ID>
<type>AA_AND2</type>
<position>-170.5,52.5</position>
<input>
<ID>IN_0</ID>476 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>772</ID>
<type>AA_AND2</type>
<position>-162,47.5</position>
<input>
<ID>IN_0</ID>476 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>773</ID>
<type>AA_AND2</type>
<position>-170.5,36</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>774</ID>
<type>AA_AND2</type>
<position>-162,31</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>775</ID>
<type>AA_AND2</type>
<position>-170.5,20</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>776</ID>
<type>AA_AND2</type>
<position>-162,15</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_AND2</type>
<position>-170.5,4</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131.5,44.5,-131.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,55.5,-131.5,55.5</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>-131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-131.5,44.5,-129,44.5</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>-131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-133,-4,-133,7</points>
<connection>
<GID>703</GID>
<name>OUT_0</name></connection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-133,-4,-129,-4</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>-133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-369,35.5,-363.5,35.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,12,-132.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,23,-132.5,23</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,12,-129,12</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,28,-132.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,39,-132.5,39</points>
<connection>
<GID>671</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,28,-129,28</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,-20,-132,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-9,-132,-9</points>
<connection>
<GID>719</GID>
<name>OUT_0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132,-20,-129,-20</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-50.5,-109.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-39.5,-109.5,-39.5</points>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,-50.5,-105.5,-50.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-35,-110,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-24,-110,-24</points>
<connection>
<GID>736</GID>
<name>OUT_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-110,-35,-105.5,-35</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-20,-109.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-9,-109.5,-9</points>
<connection>
<GID>720</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,-20,-105.5,-20</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,-20,-86,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,-9,-86,-9</points>
<connection>
<GID>721</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-20,-83,-20</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,-50.5,-86,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,-39.5,-86,-39.5</points>
<connection>
<GID>753</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-50.5,-83,-50.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,-35,-87,-24</points>
<connection>
<GID>737</GID>
<name>OUT_0</name></connection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87,-35,-83,-35</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-20,-66.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-9,-66.5,-9</points>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,-20,-62.5,-20</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-50.5,-67,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-39.5,-67,-39.5</points>
<connection>
<GID>754</GID>
<name>OUT_0</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-67,-50.5,-62.5,-50.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-35,-66.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-24,-66.5,-24</points>
<connection>
<GID>738</GID>
<name>OUT_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,-35,-62.5,-35</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-35,-44.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-24,-44.5,-24</points>
<connection>
<GID>739</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-35,-41,-35</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-50.5,-44.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-39.5,-44.5,-39.5</points>
<connection>
<GID>755</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-50.5,-41,-50.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-20,-44.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-9,-44.5,-9</points>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-20,-41,-20</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-20,-23.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-9,-23.5,-9</points>
<connection>
<GID>724</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-20,-19.5,-20</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-35,-23,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-24,-23,-24</points>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-35,-19.5,-35</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-50.5,-23.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-39.5,-23.5,-39.5</points>
<connection>
<GID>756</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-50.5,-19.5,-50.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-35,-1,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-24,-1,-24</points>
<connection>
<GID>741</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-35,2,-35</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-20,-1.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-9,-1.5,-9</points>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-20,2,-20</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-50.5,-1,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-39.5,-1,-39.5</points>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-50.5,2,-50.5</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-20,18.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-9,18.5,-9</points>
<connection>
<GID>726</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-20,22,-20</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-35,18.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-24,18.5,-24</points>
<connection>
<GID>742</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-35,22,-35</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-50.5,18.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-39.5,18.5,-39.5</points>
<connection>
<GID>758</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-50.5,22,-50.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-368,29,-365,29</points>
<connection>
<GID>846</GID>
<name>OUT_0</name></connection>
<connection>
<GID>869</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-368,21.5,-364,21.5</points>
<connection>
<GID>847</GID>
<name>OUT_0</name></connection>
<connection>
<GID>871</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-368,14.5,-364,14.5</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<connection>
<GID>848</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-352,-1.5,-352,4</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<connection>
<GID>849</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-344,-1.5,-344,4</points>
<connection>
<GID>874</GID>
<name>IN_0</name></connection>
<connection>
<GID>850</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-337,-1,-337,4</points>
<connection>
<GID>851</GID>
<name>OUT_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-331,-0.5,-331,4</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<connection>
<GID>852</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-325,-1.5,-325,4.5</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<connection>
<GID>853</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-319,-1.5,-319,4</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<connection>
<GID>854</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-313,-1,-313,4</points>
<connection>
<GID>855</GID>
<name>OUT_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-306,-1,-306,4</points>
<connection>
<GID>856</GID>
<name>OUT_0</name></connection>
<connection>
<GID>880</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-355,44,-355,52</points>
<connection>
<GID>858</GID>
<name>N_in3</name></connection>
<connection>
<GID>882</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-346.5,44,-346.5,51.5</points>
<connection>
<GID>861</GID>
<name>N_in3</name></connection>
<connection>
<GID>883</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-339,44,-339,51.5</points>
<connection>
<GID>862</GID>
<name>N_in3</name></connection>
<connection>
<GID>884</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-333,44,-333,52</points>
<connection>
<GID>863</GID>
<name>N_in3</name></connection>
<connection>
<GID>885</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-326.5,44,-326.5,52</points>
<connection>
<GID>864</GID>
<name>N_in3</name></connection>
<connection>
<GID>886</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-320.5,44,-320.5,52</points>
<connection>
<GID>865</GID>
<name>N_in3</name></connection>
<connection>
<GID>887</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-313.5,44,-313.5,52</points>
<connection>
<GID>866</GID>
<name>N_in3</name></connection>
<connection>
<GID>888</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-308,44,-308,52</points>
<connection>
<GID>867</GID>
<name>N_in3</name></connection>
<connection>
<GID>889</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-270,23.5,-246.5,23.5</points>
<connection>
<GID>786</GID>
<name>ENABLE</name></connection>
<connection>
<GID>794</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-261.5,19,-246.5,19</points>
<connection>
<GID>788</GID>
<name>OUT_0</name></connection>
<intersection>-246.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-246.5,18.5,-246.5,19</points>
<connection>
<GID>786</GID>
<name>IN_2</name></connection>
<intersection>19 1</intersection></vsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254,14.5,-254,17.5</points>
<intersection>14.5 2</intersection>
<intersection>17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-254,17.5,-246.5,17.5</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>-254 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261.5,14.5,-254,14.5</points>
<connection>
<GID>790</GID>
<name>OUT_0</name></connection>
<intersection>-254 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-252.5,11.5,-252.5,16.5</points>
<intersection>11.5 2</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-252.5,16.5,-246.5,16.5</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>-252.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261.5,11.5,-252.5,11.5</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<intersection>-252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-229.5,23.5,-229.5,69</points>
<intersection>23.5 2</intersection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-229.5,69,-173.5,69</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>-229.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,23.5,-229.5,23.5</points>
<connection>
<GID>786</GID>
<name>OUT_7</name></connection>
<intersection>-229.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,64,-178,69</points>
<intersection>64 4</intersection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,64,-165,64</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227.5,22.5,-227.5,53.5</points>
<intersection>22.5 2</intersection>
<intersection>53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-227.5,53.5,-173.5,53.5</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<intersection>-227.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,22.5,-227.5,22.5</points>
<connection>
<GID>786</GID>
<name>OUT_6</name></connection>
<intersection>-227.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,48.5,-178,53.5</points>
<intersection>48.5 4</intersection>
<intersection>53.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,48.5,-165,48.5</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224.5,21.5,-224.5,37</points>
<intersection>21.5 2</intersection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-224.5,37,-173.5,37</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>-224.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,21.5,-224.5,21.5</points>
<connection>
<GID>786</GID>
<name>OUT_5</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,32,-178,37</points>
<intersection>32 4</intersection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,32,-165,32</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-240.5,21,-173.5,21</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>-240.5 6</intersection>
<intersection>-178 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,16,-178,21</points>
<intersection>16 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,16,-165,16</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-240.5,20.5,-240.5,21</points>
<connection>
<GID>786</GID>
<name>OUT_4</name></connection>
<intersection>21 1</intersection></vsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224,5,-224,19.5</points>
<intersection>5 1</intersection>
<intersection>19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-224,5,-173.5,5</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>-224 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,19.5,-224,19.5</points>
<connection>
<GID>786</GID>
<name>OUT_3</name></connection>
<intersection>-224 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,0,-178,5</points>
<intersection>0 4</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,0,-165,0</points>
<connection>
<GID>778</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227.5,-11,-227.5,18.5</points>
<intersection>-11 1</intersection>
<intersection>18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-227.5,-11,-173.5,-11</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-227.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,18.5,-227.5,18.5</points>
<connection>
<GID>786</GID>
<name>OUT_2</name></connection>
<intersection>-227.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,-16,-178,-11</points>
<intersection>-16 4</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,-16,-165.5,-16</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230,-26,-230,17.5</points>
<intersection>-26 1</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230,-26,-173.5,-26</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>-230 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,17.5,-230,17.5</points>
<connection>
<GID>786</GID>
<name>OUT_1</name></connection>
<intersection>-230 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,-31,-178,-26</points>
<intersection>-31 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,-31,-165,-31</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233.5,-41.5,-233.5,16.5</points>
<intersection>-41.5 1</intersection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233.5,-41.5,-173.5,-41.5</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>-233.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,16.5,-233.5,16.5</points>
<connection>
<GID>786</GID>
<name>OUT_0</name></connection>
<intersection>-233.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,-46.5,-178,-41.5</points>
<intersection>-46.5 4</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,-46.5,-165,-46.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143,-71,-143,-67</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<connection>
<GID>812</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-119.5,-71,-119.5,-67</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<connection>
<GID>814</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97,-70,-97,-67</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<connection>
<GID>823</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-71,-76.5,-67</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<connection>
<GID>824</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-70.5,-55,-67</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<connection>
<GID>825</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-71,-33.5,-67</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<connection>
<GID>826</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-70.5,-12,-67</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<connection>
<GID>827</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-69.5,8,-67</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<connection>
<GID>828</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-158.5,-64,6,-64</points>
<connection>
<GID>797</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>802</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>801</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>800</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>799</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>798</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>796</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>795</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>829</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-123.5,96,-123.5,105.5</points>
<connection>
<GID>803</GID>
<name>OUT_0</name></connection>
<intersection>105.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-126,105.5,-123.5,105.5</points>
<connection>
<GID>835</GID>
<name>IN_0</name></connection>
<intersection>-123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,96,-100,105.5</points>
<connection>
<GID>804</GID>
<name>OUT_0</name></connection>
<intersection>105.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103,105.5,-100,105.5</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>-100 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,96,-78.5,105.5</points>
<connection>
<GID>805</GID>
<name>OUT_0</name></connection>
<intersection>105.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-80,105.5,-78.5,105.5</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,96,-57.5,106</points>
<connection>
<GID>806</GID>
<name>OUT_0</name></connection>
<intersection>106 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-59.5,106,-57.5,106</points>
<connection>
<GID>838</GID>
<name>IN_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,96,-36,106</points>
<connection>
<GID>807</GID>
<name>OUT_0</name></connection>
<intersection>106 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-38,106,-36,106</points>
<connection>
<GID>839</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,96,-14.5,106.5</points>
<connection>
<GID>808</GID>
<name>OUT_0</name></connection>
<intersection>106.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-16.5,106.5,-14.5,106.5</points>
<connection>
<GID>840</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,96,6,106</points>
<connection>
<GID>809</GID>
<name>OUT_0</name></connection>
<intersection>106 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>5,106,6,106</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,96,30.5,105.5</points>
<connection>
<GID>810</GID>
<name>OUT_0</name></connection>
<intersection>105.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>25,105.5,30.5,105.5</points>
<connection>
<GID>842</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-143,93.5,28.5,93.5</points>
<connection>
<GID>809</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>807</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>803</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>804</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>805</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>806</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>808</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>810</GID>
<name>ENABLE_0</name></connection>
<intersection>-143 34</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>-143,93,-143,93.5</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>93.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-187,-63.5,-187,67</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>-43.5 8</intersection>
<intersection>-28 7</intersection>
<intersection>-13 6</intersection>
<intersection>3 5</intersection>
<intersection>19 4</intersection>
<intersection>35 3</intersection>
<intersection>51.5 2</intersection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-187,67,-173.5,67</points>
<connection>
<GID>768</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-187,51.5,-173.5,51.5</points>
<connection>
<GID>771</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-187,35,-173.5,35</points>
<connection>
<GID>773</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-187,19,-173.5,19</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-187,3,-173.5,3</points>
<connection>
<GID>777</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-187,-13,-173.5,-13</points>
<connection>
<GID>779</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-187,-28,-173.5,-28</points>
<connection>
<GID>781</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-187,-43.5,-173.5,-43.5</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-182,-48.5,-182,90.5</points>
<intersection>-48.5 1</intersection>
<intersection>-33 3</intersection>
<intersection>-18 5</intersection>
<intersection>-2 7</intersection>
<intersection>14 9</intersection>
<intersection>30 10</intersection>
<intersection>46.5 11</intersection>
<intersection>62 12</intersection>
<intersection>90.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-48.5,-165,-48.5</points>
<connection>
<GID>784</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-182,-33,-165,-33</points>
<connection>
<GID>782</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-182,-18,-165.5,-18</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-182,-2,-165,-2</points>
<connection>
<GID>778</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-184,90.5,-182,90.5</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-182,14,-165,14</points>
<connection>
<GID>776</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-182,30,-165,30</points>
<connection>
<GID>774</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-182,46.5,-165,46.5</points>
<connection>
<GID>772</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-182,62,-165,62</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,68,11.5,68</points>
<connection>
<GID>645</GID>
<name>clock</name></connection>
<connection>
<GID>644</GID>
<name>clock</name></connection>
<connection>
<GID>643</GID>
<name>clock</name></connection>
<connection>
<GID>642</GID>
<name>clock</name></connection>
<connection>
<GID>641</GID>
<name>clock</name></connection>
<connection>
<GID>640</GID>
<name>clock</name></connection>
<connection>
<GID>639</GID>
<name>clock</name></connection>
<connection>
<GID>638</GID>
<name>clock</name></connection>
<connection>
<GID>768</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,63,20,63</points>
<connection>
<GID>654</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>653</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>652</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>651</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>650</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>649</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>648</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>647</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>770</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,47.5,20,47.5</points>
<connection>
<GID>772</GID>
<name>OUT</name></connection>
<connection>
<GID>663</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>664</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>665</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>666</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>667</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>668</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>669</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>670</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,52.5,11.5,52.5</points>
<connection>
<GID>771</GID>
<name>OUT</name></connection>
<connection>
<GID>655</GID>
<name>clock</name></connection>
<connection>
<GID>656</GID>
<name>clock</name></connection>
<connection>
<GID>657</GID>
<name>clock</name></connection>
<connection>
<GID>658</GID>
<name>clock</name></connection>
<connection>
<GID>659</GID>
<name>clock</name></connection>
<connection>
<GID>660</GID>
<name>clock</name></connection>
<connection>
<GID>662</GID>
<name>clock</name></connection>
<connection>
<GID>661</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,36,11.5,36</points>
<connection>
<GID>678</GID>
<name>clock</name></connection>
<connection>
<GID>677</GID>
<name>clock</name></connection>
<connection>
<GID>676</GID>
<name>clock</name></connection>
<connection>
<GID>675</GID>
<name>clock</name></connection>
<connection>
<GID>674</GID>
<name>clock</name></connection>
<connection>
<GID>673</GID>
<name>clock</name></connection>
<connection>
<GID>672</GID>
<name>clock</name></connection>
<connection>
<GID>671</GID>
<name>clock</name></connection>
<connection>
<GID>773</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,31,20,31</points>
<connection>
<GID>686</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>685</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>684</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>683</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>682</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>681</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>679</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>774</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,20,11.5,20</points>
<connection>
<GID>775</GID>
<name>OUT</name></connection>
<connection>
<GID>687</GID>
<name>clock</name></connection>
<connection>
<GID>689</GID>
<name>clock</name></connection>
<connection>
<GID>690</GID>
<name>clock</name></connection>
<connection>
<GID>691</GID>
<name>clock</name></connection>
<connection>
<GID>692</GID>
<name>clock</name></connection>
<connection>
<GID>693</GID>
<name>clock</name></connection>
<connection>
<GID>694</GID>
<name>clock</name></connection>
<connection>
<GID>688</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,15,20,15</points>
<connection>
<GID>776</GID>
<name>OUT</name></connection>
<connection>
<GID>695</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>696</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>697</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>698</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>699</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>700</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>701</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>702</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,4,11.5,4</points>
<connection>
<GID>710</GID>
<name>clock</name></connection>
<connection>
<GID>709</GID>
<name>clock</name></connection>
<connection>
<GID>708</GID>
<name>clock</name></connection>
<connection>
<GID>707</GID>
<name>clock</name></connection>
<connection>
<GID>706</GID>
<name>clock</name></connection>
<connection>
<GID>705</GID>
<name>clock</name></connection>
<connection>
<GID>704</GID>
<name>clock</name></connection>
<connection>
<GID>777</GID>
<name>OUT</name></connection>
<connection>
<GID>703</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-159,-1,20,-1</points>
<connection>
<GID>718</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>717</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>716</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>715</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>714</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>713</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>712</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>778</GID>
<name>OUT</name></connection>
<connection>
<GID>711</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,-12,11.5,-12</points>
<connection>
<GID>779</GID>
<name>OUT</name></connection>
<connection>
<GID>719</GID>
<name>clock</name></connection>
<connection>
<GID>720</GID>
<name>clock</name></connection>
<connection>
<GID>721</GID>
<name>clock</name></connection>
<connection>
<GID>722</GID>
<name>clock</name></connection>
<connection>
<GID>723</GID>
<name>clock</name></connection>
<connection>
<GID>724</GID>
<name>clock</name></connection>
<connection>
<GID>725</GID>
<name>clock</name></connection>
<connection>
<GID>726</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159.5,-17,20,-17</points>
<connection>
<GID>780</GID>
<name>OUT</name></connection>
<connection>
<GID>727</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>728</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>729</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>730</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>731</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>732</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>733</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>734</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,-27,11.5,-27</points>
<connection>
<GID>735</GID>
<name>clock</name></connection>
<connection>
<GID>781</GID>
<name>OUT</name></connection>
<connection>
<GID>736</GID>
<name>clock</name></connection>
<connection>
<GID>737</GID>
<name>clock</name></connection>
<connection>
<GID>738</GID>
<name>clock</name></connection>
<connection>
<GID>739</GID>
<name>clock</name></connection>
<connection>
<GID>740</GID>
<name>clock</name></connection>
<connection>
<GID>742</GID>
<name>clock</name></connection>
<connection>
<GID>741</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,-42.5,11.5,-42.5</points>
<connection>
<GID>783</GID>
<name>OUT</name></connection>
<connection>
<GID>751</GID>
<name>clock</name></connection>
<connection>
<GID>752</GID>
<name>clock</name></connection>
<connection>
<GID>753</GID>
<name>clock</name></connection>
<connection>
<GID>754</GID>
<name>clock</name></connection>
<connection>
<GID>755</GID>
<name>clock</name></connection>
<connection>
<GID>756</GID>
<name>clock</name></connection>
<connection>
<GID>757</GID>
<name>clock</name></connection>
<connection>
<GID>758</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,-47.5,20,-47.5</points>
<connection>
<GID>784</GID>
<name>OUT</name></connection>
<connection>
<GID>759</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>760</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>761</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>762</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>763</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>764</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>765</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>766</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,-32,20,-32</points>
<connection>
<GID>750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>749</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>748</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>745</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>746</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>744</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>743</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>782</GID>
<name>OUT</name></connection>
<connection>
<GID>747</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,-35,-132.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-24,-132.5,-24</points>
<connection>
<GID>735</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,-35,-129,-35</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,-50.5,-132,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-39.5,-132,-39.5</points>
<connection>
<GID>751</GID>
<name>OUT_0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132,-50.5,-129,-50.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143,-61.5,-143,71</points>
<connection>
<GID>795</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-143,71,-139,71</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-143,55.5,-139,55.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-143,39,-139,39</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-143,23,-139,23</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-143,7,-139,7</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-143,-9,-139,-9</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-143,-24,-139,-24</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-143,-39.5,-139,-39.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-123.5,-45,-123.5,90.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 6</intersection>
<intersection>1.5 7</intersection>
<intersection>17.5 8</intersection>
<intersection>33.5 9</intersection>
<intersection>50 10</intersection>
<intersection>65.5 11</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-129,-45,-123.5,-45</points>
<connection>
<GID>759</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-129,-14.5,-123.5,-14.5</points>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-129,1.5,-123.5,1.5</points>
<connection>
<GID>711</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-129,17.5,-123.5,17.5</points>
<connection>
<GID>695</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-129,33.5,-123.5,33.5</points>
<connection>
<GID>679</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-129,50,-123.5,50</points>
<connection>
<GID>663</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-129,65.5,-123.5,65.5</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-129,-29.5,-123.5,-29.5</points>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-119.5,-61.5,-119.5,71</points>
<connection>
<GID>796</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 7</intersection>
<intersection>-24 8</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-119.5,71,-116.5,71</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,55.5,-116.5,55.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-119.5,39,-116.5,39</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-119.5,23,-116.5,23</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119.5,7,-116.5,7</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119.5,-9,-116.5,-9</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-119.5,-39.5,-116.5,-39.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-119.5,-24,-116.5,-24</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-45,-100,90.5</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 9</intersection>
<intersection>33.5 8</intersection>
<intersection>50 6</intersection>
<intersection>65.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-105.5,-45,-100,-45</points>
<connection>
<GID>760</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-105.5,50,-100,50</points>
<connection>
<GID>664</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-105.5,65.5,-100,65.5</points>
<connection>
<GID>648</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-105.5,33.5,-100,33.5</points>
<connection>
<GID>680</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-105.5,17.5,-100,17.5</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-105.5,1.5,-100,1.5</points>
<connection>
<GID>712</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-105.5,-14.5,-100,-14.5</points>
<connection>
<GID>728</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-105.5,-29.5,-100,-29.5</points>
<connection>
<GID>744</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97,-61.5,-97,71</points>
<connection>
<GID>797</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-97,71,-93,71</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,55.5,-93,55.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-97,39,-93,39</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-97,23,-93,23</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-97,7,-93,7</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-97,-9,-93,-9</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-97,-24,-93,-24</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-97,-39.5,-93,-39.5</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,-45,-78.5,90.5</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 7</intersection>
<intersection>1.5 11</intersection>
<intersection>17.5 10</intersection>
<intersection>33.5 8</intersection>
<intersection>50 9</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-83,-45,-78.5,-45</points>
<connection>
<GID>761</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-83,65.5,-78.5,65.5</points>
<connection>
<GID>649</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-83,-14.5,-78.5,-14.5</points>
<connection>
<GID>729</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-83,33.5,-78.5,33.5</points>
<connection>
<GID>681</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-83,50,-78.5,50</points>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-83,17.5,-78.5,17.5</points>
<connection>
<GID>697</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-83,1.5,-78.5,1.5</points>
<connection>
<GID>713</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-83,-29.5,-78.5,-29.5</points>
<connection>
<GID>745</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-61.5,-76.5,71</points>
<connection>
<GID>798</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 2</intersection>
<intersection>55.5 3</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,71,-74,71</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76.5,39,-74,39</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-76.5,55.5,-74,55.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-76.5,23,-74,23</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-76.5,7,-74,7</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-76.5,-9,-74,-9</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-76.5,-24,-74,-24</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-76.5,-39.5,-74,-39.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-45,-57.5,90.5</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 8</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 11</intersection>
<intersection>33.5 9</intersection>
<intersection>50 6</intersection>
<intersection>65.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-62.5,-45,-57.5,-45</points>
<connection>
<GID>762</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-62.5,50,-57.5,50</points>
<connection>
<GID>666</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-62.5,65.5,-57.5,65.5</points>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-62.5,-14.5,-57.5,-14.5</points>
<connection>
<GID>730</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-62.5,33.5,-57.5,33.5</points>
<connection>
<GID>682</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-62.5,1.5,-57.5,1.5</points>
<connection>
<GID>714</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-62.5,17.5,-57.5,17.5</points>
<connection>
<GID>698</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-62.5,-29.5,-57.5,-29.5</points>
<connection>
<GID>746</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-61.5,-55,71</points>
<connection>
<GID>799</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 3</intersection>
<intersection>7 4</intersection>
<intersection>23 5</intersection>
<intersection>39 6</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,71,-51.5,71</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,55.5,-51.5,55.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55,-9,-51.5,-9</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-55,7,-51.5,7</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-55,23,-51.5,23</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-55,39,-51.5,39</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-55,-24,-51.5,-24</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-55,-39.5,-51.5,-39.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-45,-36,90.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 9</intersection>
<intersection>33.5 8</intersection>
<intersection>50 7</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-41,-45,-36,-45</points>
<connection>
<GID>763</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-41,65.5,-36,65.5</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-41,50,-36,50</points>
<connection>
<GID>667</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-41,33.5,-36,33.5</points>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-41,17.5,-36,17.5</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-41,1.5,-36,1.5</points>
<connection>
<GID>715</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-41,-14.5,-36,-14.5</points>
<connection>
<GID>731</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-41,-29.5,-36,-29.5</points>
<connection>
<GID>747</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-61.5,-33.5,71</points>
<connection>
<GID>800</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 3</intersection>
<intersection>7 4</intersection>
<intersection>23 5</intersection>
<intersection>39 6</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,71,-30,71</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,55.5,-30,55.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-33.5,-9,-30,-9</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-33.5,7,-30,7</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-33.5,23,-30,23</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-33.5,39,-30,39</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-33.5,-24,-30,-24</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-33.5,-39.5,-30,-39.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-45,-14.5,90.5</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 10</intersection>
<intersection>-14.5 9</intersection>
<intersection>1.5 8</intersection>
<intersection>17.5 7</intersection>
<intersection>33.5 6</intersection>
<intersection>50 5</intersection>
<intersection>65.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-45,-14.5,-45</points>
<connection>
<GID>764</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-19.5,65.5,-14.5,65.5</points>
<connection>
<GID>652</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-19.5,50,-14.5,50</points>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-19.5,33.5,-14.5,33.5</points>
<connection>
<GID>684</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-19.5,17.5,-14.5,17.5</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-19.5,1.5,-14.5,1.5</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-19.5,-14.5,-14.5,-14.5</points>
<connection>
<GID>732</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-19.5,-29.5,-14.5,-29.5</points>
<connection>
<GID>748</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-61.5,-12,71</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,71,-8.5,71</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12,55.5,-8.5,55.5</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12,39,-8.5,39</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-12,23,-8.5,23</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12,7,-8.5,7</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-12,-9,-8.5,-9</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-12,-24,-8.5,-24</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-12,-39.5,-8.5,-39.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-45,6,90.5</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>-45 5</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 9</intersection>
<intersection>33.5 8</intersection>
<intersection>50 7</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>2,-45,6,-45</points>
<connection>
<GID>765</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>2,65.5,6,65.5</points>
<connection>
<GID>653</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>2,50,6,50</points>
<connection>
<GID>669</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>2,33.5,6,33.5</points>
<connection>
<GID>685</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>2,17.5,6,17.5</points>
<connection>
<GID>701</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>2,1.5,6,1.5</points>
<connection>
<GID>717</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>2,-14.5,6,-14.5</points>
<connection>
<GID>733</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>2,-29.5,6,-29.5</points>
<connection>
<GID>749</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-61.5,8,71</points>
<connection>
<GID>802</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 7</intersection>
<intersection>-24 5</intersection>
<intersection>-9 6</intersection>
<intersection>7 8</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,71,11.5,71</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,55.5,11.5,55.5</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,39,11.5,39</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8,23,11.5,23</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>8,-24,11.5,-24</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>8,-9,11.5,-9</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>8,-39.5,11.5,-39.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>8,7,11.5,7</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-45,30.5,90.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 8</intersection>
<intersection>33.5 9</intersection>
<intersection>50 7</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22,-45,30.5,-45</points>
<connection>
<GID>766</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>22,65.5,30.5,65.5</points>
<connection>
<GID>654</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22,50,30.5,50</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>22,17.5,30.5,17.5</points>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22,33.5,30.5,33.5</points>
<connection>
<GID>686</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>22,1.5,30.5,1.5</points>
<connection>
<GID>718</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>22,-14.5,30.5,-14.5</points>
<connection>
<GID>734</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>22,-29.5,30.5,-29.5</points>
<connection>
<GID>750</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,60,19,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,71,19,71</points>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,60,22,60</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,44.5,18.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,55.5,18.5,55.5</points>
<connection>
<GID>662</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,44.5,22,44.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,60,-2,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,71,-2,71</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,60,2,60</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,44.5,-2,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,55.5,-2,55.5</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,44.5,2,44.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-4,18,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,7,18,7</points>
<connection>
<GID>710</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-4,22,-4</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,12,18.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,23,18.5,23</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,12,22,12</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,28,18.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,39,18.5,39</points>
<connection>
<GID>678</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,28,22,28</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,28,-1.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,39,-1.5,39</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,28,2,28</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,12,-1.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,23,-1.5,23</points>
<connection>
<GID>693</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,12,2,12</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-4,-2,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,7,-2,7</points>
<connection>
<GID>709</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-4,2,-4</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,60,-23,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,71,-23,71</points>
<connection>
<GID>643</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,60,-19.5,60</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,44.5,-23,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,55.5,-23,55.5</points>
<connection>
<GID>660</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,44.5,-19.5,44.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,28,-22.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,39,-22.5,39</points>
<connection>
<GID>676</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,28,-19.5,28</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,12,-22,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,23,-22,23</points>
<connection>
<GID>692</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22,12,-19.5,12</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-4,-23,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,7,-23,7</points>
<connection>
<GID>708</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-4,-19.5,-4</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-4,-44,7</points>
<intersection>-4 2</intersection>
<intersection>7 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-44,-4,-41,-4</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-45.5,7,-44,7</points>
<connection>
<GID>707</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,12,-44.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,23,-44.5,23</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,12,-41,12</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,28,-44.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,39,-44.5,39</points>
<connection>
<GID>675</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,28,-41,28</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,44.5,-44.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,55.5,-44.5,55.5</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,44.5,-41,44.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,60,-44,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,71,-44,71</points>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44,60,-41,60</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,60,-65.5,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,71,-65.5,71</points>
<connection>
<GID>641</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,60,-62.5,60</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,44.5,-66,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,55.5,-66,55.5</points>
<connection>
<GID>658</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,44.5,-62.5,44.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,28,-66,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,39,-66,39</points>
<connection>
<GID>674</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,28,-62.5,28</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,12,-66,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,23,-66,23</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,12,-62.5,12</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,-4,-66,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,7,-66,7</points>
<connection>
<GID>706</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,-4,-62.5,-4</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,-4,-86.5,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,7,-86.5,7</points>
<connection>
<GID>705</GID>
<name>OUT_0</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-4,-83,-4</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>-86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,12,-87,23</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87,12,-83,12</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,28,-86,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,39,-86,39</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,28,-83,28</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,44.5,-86.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,55.5,-86.5,55.5</points>
<connection>
<GID>657</GID>
<name>OUT_0</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,44.5,-83,44.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>-86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,60,-86,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,71,-86,71</points>
<connection>
<GID>640</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,60,-83,60</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,60,-109.5,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,71,-109.5,71</points>
<connection>
<GID>639</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,60,-105.5,60</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,44.5,-109.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,55.5,-109.5,55.5</points>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,44.5,-105.5,44.5</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,28,-109,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,39,-109,39</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109,28,-105.5,28</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,12,-109.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,23,-109.5,23</points>
<connection>
<GID>688</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,12,-105.5,12</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-4,-109.5,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,7,-109.5,7</points>
<connection>
<GID>704</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,-4,-105.5,-4</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,60,-132,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,71,-132,71</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132,60,-129,60</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>565.807,125.608,1093.79,-135.365</PageViewport>
<gate>
<ID>1</ID>
<type>AI_XOR2</type>
<position>752.5,23.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>766.5,18</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>766.5,8.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AI_XOR2</type>
<position>711,18</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>776.5,5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>711,8.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_OR2</type>
<position>721,5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>718,18</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>678,27.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>678,22.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>773.5,18</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>692,4</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>727.5,2.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>720,16</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>HA_JUNC_2</type>
<position>679.5,5</position>
<input>
<ID>N_in0</ID>31 </input>
<input>
<ID>N_in1</ID>25 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>733,27.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AI_XOR2</type>
<position>977,23</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>733.5,22.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>AI_XOR2</type>
<position>991,17.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>747.5,4</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>991,8</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AI_XOR2</type>
<position>935.5,17.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>783,2.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AE_OR2</type>
<position>1001,4.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>935.5,8</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>775.5,16</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AE_OR2</type>
<position>945.5,4.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AI_XOR2</type>
<position>807.5,23.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>942.5,17.5</position>
<input>
<ID>N_in0</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AI_XOR2</type>
<position>821.5,18</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>821.5,8.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_OR2</type>
<position>831.5,5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>902.5,27</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>828.5,18</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>902.5,22</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>998,17.5</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>788.5,27.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>788.5,22.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>916.5,3.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND2</type>
<position>802.5,4</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>838,2.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>830.5,16</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>952,2</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>944.5,15.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>HA_JUNC_2</type>
<position>904,4.5</position>
<input>
<ID>N_in0</ID>62 </input>
<input>
<ID>N_in1</ID>56 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>958,27</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>958,22</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>972,3.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>1007.5,2</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>1000,15.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AI_XOR2</type>
<position>1032,23</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AI_XOR2</type>
<position>1046,17.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>1046,8</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR2</type>
<position>1056,4.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>HA_JUNC_2</type>
<position>790,5</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>10 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>1053,17.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AI_XOR2</type>
<position>642,23.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>1062,4.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AI_XOR2</type>
<position>656,18</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>1013,27</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>656,8.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>1013,22</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_OR2</type>
<position>666,5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>1027,3.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>663,18</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>1062.5,2</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>623,27.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>1055,15.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_TOGGLE</type>
<position>623,22.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>92</ID>
<type>HA_JUNC_2</type>
<position>1014.5,4.5</position>
<input>
<ID>N_in0</ID>47 </input>
<input>
<ID>N_in1</ID>40 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_AND2</type>
<position>637,4</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AI_XOR2</type>
<position>866.5,23</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>623,9.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AI_XOR2</type>
<position>880.5,17.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>672.5,2.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND2</type>
<position>880.5,8</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>665,16</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AE_OR2</type>
<position>890.5,4.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>887.5,17.5</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AI_XOR2</type>
<position>697,23.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>847.5,27</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>847.5,22</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>861.5,3.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>897,2</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>889.5,15.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AI_XOR2</type>
<position>921.5,23</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>HA_JUNC_2</type>
<position>734.5,5</position>
<input>
<ID>N_in0</ID>63 </input>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>HA_JUNC_2</type>
<position>843,5</position>
<input>
<ID>N_in0</ID>64 </input>
<input>
<ID>N_in1</ID>49 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>HA_JUNC_2</type>
<position>957.5,4.5</position>
<input>
<ID>N_in0</ID>65 </input>
<input>
<ID>N_in1</ID>33 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>771.5,6,771.5,8.5</points>
<intersection>6 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>771.5,6,773.5,6</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>771.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>769.5,8.5,771.5,8.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>771.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>762.5,17,763.5,17</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>762.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>762.5,9.5,762.5,17</points>
<intersection>9.5 4</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>735.5,9.5,763.5,9.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>735.5 10</intersection>
<intersection>762.5 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>735.5,5,735.5,9.5</points>
<connection>
<GID>109</GID>
<name>N_in1</name></connection>
<intersection>9.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>755.5,23.5,760,23.5</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>760 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>760,7.5,760,23.5</points>
<intersection>7.5 5</intersection>
<intersection>19 6</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>760,7.5,763.5,7.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>760 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>760,19,763.5,19</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>760 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>769.5,18,772.5,18</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>23</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>735,27.5,744.5,27.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>744.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>744.5,5,744.5,27.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>24.5 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>744.5,24.5,749.5,24.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>744.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>735.5,22.5,749.5,22.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>739 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>739,3,739,22.5</points>
<intersection>3 4</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>739,3,744.5,3</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>739 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>750.5,4,773.5,4</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>826.5,6,826.5,8.5</points>
<intersection>6 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>826.5,6,828.5,6</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>826.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>824.5,8.5,826.5,8.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>826.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>817.5,17,818.5,17</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>817.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>817.5,9.5,817.5,17</points>
<intersection>9.5 4</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>791,9.5,818.5,9.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>791 7</intersection>
<intersection>817.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>791,5,791,9.5</points>
<connection>
<GID>77</GID>
<name>N_in1</name></connection>
<intersection>9.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>810.5,23.5,815,23.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>815 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>815,7.5,815,23.5</points>
<intersection>7.5 5</intersection>
<intersection>19 6</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>815,7.5,818.5,7.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>815 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>815,19,818.5,19</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>815 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>824.5,18,827.5,18</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>56</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>790.5,27.5,799.5,27.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>799.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>799.5,5,799.5,27.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>24.5 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>799.5,24.5,804.5,24.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>799.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>790.5,22.5,804.5,22.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>794 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>794,3,794,22.5</points>
<intersection>3 4</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>794,3,799.5,3</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>794 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>805.5,4,828.5,4</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>779.5,5,789,5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>77</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>661,6,661,8.5</points>
<intersection>6 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>661,6,663,6</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>661 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,8.5,661,8.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>661 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>652,17,653,17</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>652 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>652,9.5,652,17</points>
<intersection>9.5 4</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>625,9.5,653,9.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>652 3</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>645,23.5,649.5,23.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>649.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>649.5,7.5,649.5,23.5</points>
<intersection>7.5 5</intersection>
<intersection>19 6</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>649.5,7.5,653,7.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>649.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>649.5,19,653,19</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>649.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>659,18,662,18</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>625,27.5,634,27.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>634 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>634,5,634,27.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>24.5 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>634,24.5,639,24.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>634 4</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>625,22.5,639,22.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>628 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>628,3,628,22.5</points>
<intersection>3 4</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>628,3,634,3</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>628 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,4,663,4</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>716,6,716,8.5</points>
<intersection>6 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>716,6,718,6</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>716 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>714,8.5,716,8.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>716 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>707,17,708,17</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>707 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>707,9.5,707,17</points>
<intersection>9.5 4</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>680.5,9.5,708,9.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>680.5 7</intersection>
<intersection>707 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>680.5,5,680.5,9.5</points>
<connection>
<GID>34</GID>
<name>N_in1</name></connection>
<intersection>9.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>700,23.5,704.5,23.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>704.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>704.5,7.5,704.5,23.5</points>
<intersection>7.5 5</intersection>
<intersection>19 6</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>704.5,7.5,708,7.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>704.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>704.5,19,708,19</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>704.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>714,18,717,18</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>680,27.5,689,27.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>689 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>689,5,689,27.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>24.5 6</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>689,24.5,694,24.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>689 4</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>680,22.5,694,22.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>684.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>684.5,3,684.5,22.5</points>
<intersection>3 4</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>684.5,3,689,3</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>684.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>695,4,718,4</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>669,5,678.5,5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<connection>
<GID>34</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>996,5.5,996,8</points>
<intersection>5.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>996,5.5,998,5.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>996 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>994,8,996,8</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>996 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>987,16.5,988,16.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>987 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>987,9,987,16.5</points>
<intersection>9 4</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>960,9,988,9</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>960 7</intersection>
<intersection>987 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>960,4.5,960,9</points>
<intersection>4.5 8</intersection>
<intersection>9 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>958.5,4.5,960,4.5</points>
<connection>
<GID>111</GID>
<name>N_in1</name></connection>
<intersection>960 7</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>980,23,984.5,23</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>984.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>984.5,7,984.5,23</points>
<intersection>7 5</intersection>
<intersection>18.5 6</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>984.5,7,988,7</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>984.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>984.5,18.5,988,18.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>984.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>994,17.5,997,17.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>960,27,969,27</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>969 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>969,4.5,969,27</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>24 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>969,24,974,24</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>969 4</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>960,22,974,22</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>963.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>963.5,2.5,963.5,22</points>
<intersection>2.5 4</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>963.5,2.5,969,2.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>963.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>975,3.5,998,3.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1051,5.5,1051,8</points>
<intersection>5.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1051,5.5,1053,5.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>1051 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1049,8,1051,8</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>1051 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1042,16.5,1043,16.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>1042 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1042,9,1042,16.5</points>
<intersection>9 4</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1015.5,9,1043,9</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>1015.5 7</intersection>
<intersection>1042 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1015.5,4.5,1015.5,9</points>
<connection>
<GID>92</GID>
<name>N_in1</name></connection>
<intersection>9 4</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1035,23,1039.5,23</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>1039.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1039.5,7,1039.5,23</points>
<intersection>7 5</intersection>
<intersection>18.5 6</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>1039.5,7,1043,7</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>1039.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>1039.5,18.5,1043,18.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>1039.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1049,17.5,1052,17.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<connection>
<GID>78</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1059,4.5,1061,4.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1015,27,1024,27</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>1024 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>1024,4.5,1024,27</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>24 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>1024,24,1029,24</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>1024 4</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>1015,22,1029,22</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>1018.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1018.5,2.5,1018.5,22</points>
<intersection>2.5 4</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1018.5,2.5,1024,2.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>1018.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1030,3.5,1053,3.5</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1004,4.5,1013.5,4.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>885.5,5.5,885.5,8</points>
<intersection>5.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>885.5,5.5,887.5,5.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>885.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>883.5,8,885.5,8</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>885.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>876.5,16.5,877.5,16.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>876.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>876.5,9,876.5,16.5</points>
<intersection>9 4</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>844,9,877.5,9</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>844 7</intersection>
<intersection>876.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>844,5,844,9</points>
<connection>
<GID>110</GID>
<name>N_in1</name></connection>
<intersection>9 4</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>869.5,23,874,23</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>874 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>874,7,874,23</points>
<intersection>7 5</intersection>
<intersection>18.5 6</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>874,7,877.5,7</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>874 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>874,18.5,877.5,18.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>874 3</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>883.5,17.5,886.5,17.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<connection>
<GID>101</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>849.5,27,858.5,27</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>858.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>858.5,4.5,858.5,27</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>24 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>858.5,24,863.5,24</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>858.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>849.5,22,863.5,22</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>852.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>852.5,2.5,852.5,22</points>
<intersection>2.5 4</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>852.5,2.5,858.5,2.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>852.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>864.5,3.5,887.5,3.5</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>940.5,5.5,940.5,8</points>
<intersection>5.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>940.5,5.5,942.5,5.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>940.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>938.5,8,940.5,8</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>940.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>931.5,16.5,932.5,16.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>931.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>931.5,9,931.5,16.5</points>
<intersection>9 4</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>905,9,932.5,9</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>905 7</intersection>
<intersection>931.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>905,4.5,905,9</points>
<connection>
<GID>67</GID>
<name>N_in1</name></connection>
<intersection>9 4</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>924.5,23,929,23</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>929 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>929,7,929,23</points>
<intersection>7 5</intersection>
<intersection>18.5 6</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>929,7,932.5,7</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>929 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>929,18.5,932.5,18.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>929 3</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>938.5,17.5,941.5,17.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>51</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>904.5,27,913.5,27</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>913.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>913.5,4.5,913.5,27</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>24 6</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>913.5,24,918.5,24</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>913.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>904.5,22,918.5,22</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>909 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>909,2.5,909,22</points>
<intersection>2.5 4</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>909,2.5,913.5,2.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>909 3</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>919.5,3.5,942.5,3.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>893.5,4.5,903,4.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724,5,733.5,5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>109</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>834.5,5,842,5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>948.5,4.5,956.5,4.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<connection>
<GID>111</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>85.312,165.484,308.056,55.3859</PageViewport>
<gate>
<ID>389</ID>
<type>AE_OR2</type>
<position>737,149.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>GA_LED</type>
<position>734,162.5</position>
<input>
<ID>N_in0</ID>224 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>393</ID>
<type>GA_LED</type>
<position>903.5,162</position>
<input>
<ID>N_in0</ID>247 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>AA_AND2</type>
<position>822,148</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_AND2</type>
<position>708,148.5</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>226 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_LABEL</type>
<position>743.5,147</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>399</ID>
<type>AA_LABEL</type>
<position>736,160.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>857.5,146.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>AA_LABEL</type>
<position>850,160</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>HA_JUNC_2</type>
<position>809.5,149</position>
<input>
<ID>N_in0</ID>274 </input>
<input>
<ID>N_in1</ID>268 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>877.5,148</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_LABEL</type>
<position>913,146.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>407</ID>
<type>AA_LABEL</type>
<position>905.5,160</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>408</ID>
<type>AI_XOR2</type>
<position>937.5,167.5</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>257 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AI_XOR2</type>
<position>951.5,162</position>
<input>
<ID>IN_0</ID>253 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>951.5,152.5</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AE_OR2</type>
<position>961.5,149</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>258 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>HA_JUNC_2</type>
<position>695.5,149.5</position>
<input>
<ID>N_in0</ID>228 </input>
<input>
<ID>N_in1</ID>222 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>413</ID>
<type>GA_LED</type>
<position>958.5,162</position>
<input>
<ID>N_in0</ID>254 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>414</ID>
<type>AI_XOR2</type>
<position>547.5,168</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>415</ID>
<type>GA_LED</type>
<position>967.5,149</position>
<input>
<ID>N_in0</ID>255 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>416</ID>
<type>AI_XOR2</type>
<position>561.5,162.5</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_AND2</type>
<position>561.5,153</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>AE_OR2</type>
<position>571.5,149.5</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>AA_AND2</type>
<position>932.5,148</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>257 </input>
<output>
<ID>OUT</ID>258 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>422</ID>
<type>GA_LED</type>
<position>568.5,162.5</position>
<input>
<ID>N_in0</ID>232 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>968,146.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>425</ID>
<type>AA_LABEL</type>
<position>960.5,160</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>HA_JUNC_2</type>
<position>920,149</position>
<input>
<ID>N_in0</ID>259 </input>
<input>
<ID>N_in1</ID>252 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>AA_AND2</type>
<position>542.5,148.5</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>AI_XOR2</type>
<position>772,167.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>AA_TOGGLE</type>
<position>528.5,154</position>
<output>
<ID>OUT_0</ID>230 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>431</ID>
<type>AI_XOR2</type>
<position>786,162</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>261 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>432</ID>
<type>AA_LABEL</type>
<position>578,147</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AA_AND2</type>
<position>786,152.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>262 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>570.5,160.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AE_OR2</type>
<position>796,149</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>266 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>GA_LED</type>
<position>793,162</position>
<input>
<ID>N_in0</ID>263 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AI_XOR2</type>
<position>602.5,168</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_AND2</type>
<position>767,148</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>441</ID>
<type>AA_LABEL</type>
<position>802.5,146.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>AA_LABEL</type>
<position>795,160</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>443</ID>
<type>AI_XOR2</type>
<position>827,167.5</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>444</ID>
<type>HA_JUNC_2</type>
<position>640,149.5</position>
<input>
<ID>N_in0</ID>275 </input>
<input>
<ID>N_in1</ID>215 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>445</ID>
<type>HA_JUNC_2</type>
<position>748.5,149.5</position>
<input>
<ID>N_in0</ID>276 </input>
<input>
<ID>N_in1</ID>261 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>446</ID>
<type>HA_JUNC_2</type>
<position>863,149</position>
<input>
<ID>N_in0</ID>277 </input>
<input>
<ID>N_in1</ID>245 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>513.5,191.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>569.5,191</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>626.5,191.5</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>679.5,191</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>740,191.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>794.5,190</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>453</ID>
<type>DA_FROM</type>
<position>849.5,190</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>904,190.5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>456</ID>
<type>BA_TRI_STATE</type>
<position>512.5,181</position>
<input>
<ID>ENABLE_0</ID>279 </input>
<input>
<ID>IN_0</ID>281 </input>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>457</ID>
<type>BA_TRI_STATE</type>
<position>522.5,181</position>
<input>
<ID>ENABLE_0</ID>284 </input>
<input>
<ID>IN_0</ID>281 </input>
<output>
<ID>OUT_0</ID>233 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>459</ID>
<type>AE_SMALL_INVERTER</type>
<position>518,181</position>
<input>
<ID>IN_0</ID>284 </input>
<output>
<ID>OUT_0</ID>279 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>468</ID>
<type>BA_TRI_STATE</type>
<position>568,181</position>
<input>
<ID>ENABLE_0</ID>285 </input>
<input>
<ID>IN_0</ID>286 </input>
<output>
<ID>OUT_0</ID>241 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>469</ID>
<type>BA_TRI_STATE</type>
<position>578,181</position>
<input>
<ID>ENABLE_0</ID>287 </input>
<input>
<ID>IN_0</ID>286 </input>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>470</ID>
<type>AE_SMALL_INVERTER</type>
<position>573.5,181</position>
<input>
<ID>IN_0</ID>287 </input>
<output>
<ID>OUT_0</ID>285 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>471</ID>
<type>BA_TRI_STATE</type>
<position>624.5,181</position>
<input>
<ID>ENABLE_0</ID>288 </input>
<input>
<ID>IN_0</ID>289 </input>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>472</ID>
<type>BA_TRI_STATE</type>
<position>634.5,181</position>
<input>
<ID>ENABLE_0</ID>290 </input>
<input>
<ID>IN_0</ID>289 </input>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>473</ID>
<type>AE_SMALL_INVERTER</type>
<position>630,181</position>
<input>
<ID>IN_0</ID>290 </input>
<output>
<ID>OUT_0</ID>288 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>474</ID>
<type>BA_TRI_STATE</type>
<position>678,180</position>
<input>
<ID>ENABLE_0</ID>291 </input>
<input>
<ID>IN_0</ID>292 </input>
<output>
<ID>OUT_0</ID>226 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>475</ID>
<type>BA_TRI_STATE</type>
<position>688,180</position>
<input>
<ID>ENABLE_0</ID>293 </input>
<input>
<ID>IN_0</ID>292 </input>
<output>
<ID>OUT_0</ID>225 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>476</ID>
<type>AE_SMALL_INVERTER</type>
<position>683.5,180</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>291 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>477</ID>
<type>BA_TRI_STATE</type>
<position>738,180</position>
<input>
<ID>ENABLE_0</ID>294 </input>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>265 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>478</ID>
<type>BA_TRI_STATE</type>
<position>748,180</position>
<input>
<ID>ENABLE_0</ID>296 </input>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>264 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>479</ID>
<type>AE_SMALL_INVERTER</type>
<position>743.5,180</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>294 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>480</ID>
<type>BA_TRI_STATE</type>
<position>793,179</position>
<input>
<ID>ENABLE_0</ID>297 </input>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>272 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>481</ID>
<type>BA_TRI_STATE</type>
<position>803,179</position>
<input>
<ID>ENABLE_0</ID>299 </input>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>271 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>482</ID>
<type>AE_SMALL_INVERTER</type>
<position>798.5,179</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>297 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>483</ID>
<type>BA_TRI_STATE</type>
<position>847.5,178.5</position>
<input>
<ID>ENABLE_0</ID>300 </input>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>484</ID>
<type>BA_TRI_STATE</type>
<position>857.5,178.5</position>
<input>
<ID>ENABLE_0</ID>302 </input>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>485</ID>
<type>AE_SMALL_INVERTER</type>
<position>853,178.5</position>
<input>
<ID>IN_0</ID>302 </input>
<output>
<ID>OUT_0</ID>300 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>486</ID>
<type>BA_TRI_STATE</type>
<position>902.5,178</position>
<input>
<ID>ENABLE_0</ID>303 </input>
<input>
<ID>IN_0</ID>304 </input>
<output>
<ID>OUT_0</ID>257 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>487</ID>
<type>BA_TRI_STATE</type>
<position>912.5,178</position>
<input>
<ID>ENABLE_0</ID>305 </input>
<input>
<ID>IN_0</ID>304 </input>
<output>
<ID>OUT_0</ID>256 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>488</ID>
<type>AE_SMALL_INVERTER</type>
<position>908,178</position>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>303 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>490</ID>
<type>DA_FROM</type>
<position>529,181</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>494</ID>
<type>DA_FROM</type>
<position>584,181</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>641,181</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>496</ID>
<type>DA_FROM</type>
<position>694.5,180</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>755,180</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>498</ID>
<type>DA_FROM</type>
<position>809.5,179</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>499</ID>
<type>DA_FROM</type>
<position>864.5,178.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>500</ID>
<type>DA_FROM</type>
<position>920.5,178</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>304,96.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>295.5,85.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>DE_TO</type>
<position>194,154</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOC</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_AND2</type>
<position>303.5,80.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>98,74</position>
<gparam>LABEL_TEXT now we got every bytes cleared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>AA_TOGGLE</type>
<position>180,154</position>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>295.5,70.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>304,65.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>96.5,67.5</position>
<gparam>LABEL_TEXT we can write data to registers</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>295.5,55</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>304,50</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>189.5,122</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>BE_DECODER_3x8</type>
<position>222.5,117.5</position>
<input>
<ID>ENABLE</ID>210 </input>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>212 </input>
<input>
<ID>IN_2</ID>211 </input>
<output>
<ID>OUT_0</ID>74 </output>
<output>
<ID>OUT_1</ID>73 </output>
<output>
<ID>OUT_2</ID>72 </output>
<output>
<ID>OUT_3</ID>71 </output>
<output>
<ID>OUT_4</ID>70 </output>
<output>
<ID>OUT_5</ID>69 </output>
<output>
<ID>OUT_6</ID>68 </output>
<output>
<ID>OUT_7</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>106,60.5</position>
<gparam>LABEL_TEXT always on to make decoder on</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>202.5,116.5</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>192,116.5</position>
<gparam>LABEL_TEXT i1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>192,112</position>
<gparam>LABEL_TEXT i2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_TOGGLE</type>
<position>202.5,112</position>
<output>
<ID>OUT_0</ID>212 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>192,107.5</position>
<gparam>LABEL_TEXT i3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_TOGGLE</type>
<position>202.5,109</position>
<output>
<ID>OUT_0</ID>213 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>196.5,103</position>
<gparam>LABEL_TEXT input combitaions that is address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>194,121</position>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>180.5,91.5</position>
<gparam>LABEL_TEXT fst comb 000</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>BA_TRI_STATE</type>
<position>323,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_TRI_STATE</type>
<position>346.5,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>219.5,62</position>
<gparam>LABEL_TEXT selected register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>BA_TRI_STATE</type>
<position>369,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>BA_TRI_STATE</type>
<position>389.5,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>205.5,91.5</position>
<gparam>LABEL_TEXT 00001111</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>BA_TRI_STATE</type>
<position>411,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>BA_TRI_STATE</type>
<position>432.5,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>123 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>176.5,98</position>
<gparam>LABEL_TEXT i/p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>BA_TRI_STATE</type>
<position>454,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>143</ID>
<type>BA_TRI_STATE</type>
<position>474,33.5</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>205,97</position>
<gparam>LABEL_TEXT DATA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>BA_TRI_STATE</type>
<position>342.5,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>146</ID>
<type>BA_TRI_STATE</type>
<position>366,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>116 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>94,102</position>
<gparam>LABEL_TEXT WRITE using clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>BA_TRI_STATE</type>
<position>387.5,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>118 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>180,85.5</position>
<gparam>LABEL_TEXT sec combo 011</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>BA_TRI_STATE</type>
<position>408.5,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>120 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>205.5,85</position>
<gparam>LABEL_TEXT 11110000</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>BA_TRI_STATE</type>
<position>430,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>122 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>180,79</position>
<gparam>LABEL_TEXT third combo 111</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>BA_TRI_STATE</type>
<position>451.5,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>205,78.5</position>
<gparam>LABEL_TEXT 00111100</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>BA_TRI_STATE</type>
<position>472,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>BA_TRI_STATE</type>
<position>496.5,191</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>128 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>191,144.5</position>
<gparam>LABEL_TEXT now we read wat data we gave</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>323,24.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_TOGGLE</type>
<position>95,133</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>346.5,24.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>104.5,133</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>81.5,134</position>
<gparam>LABEL_TEXT without delay</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>369,25.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>389.5,24.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>411,25</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>432.5,24.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>168</ID>
<type>DA_FROM</type>
<position>454,25</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>474,26</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>305.5,33.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>321,190.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>282,190</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>340,205</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>363,205</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>386,205</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>176</ID>
<type>DE_TO</type>
<position>406.5,205.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>177</ID>
<type>DE_TO</type>
<position>428,205.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>178</ID>
<type>DE_TO</type>
<position>449.5,206</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>471,205.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_TO</type>
<position>491,205</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>279,32</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_TOGGLE</type>
<position>96,126.5</position>
<output>
<ID>OUT_0</ID>191 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>96,119</position>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_TOGGLE</type>
<position>95.5,113.5</position>
<output>
<ID>OUT_0</ID>193 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_TOGGLE</type>
<position>114,94</position>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>186</ID>
<type>AA_TOGGLE</type>
<position>122,94</position>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_TOGGLE</type>
<position>129,94.5</position>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>135,95</position>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_TOGGLE</type>
<position>141,94</position>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>147.5,94</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>153,94.5</position>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>160,94.5</position>
<output>
<ID>OUT_0</ID>201 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>193</ID>
<type>GA_LED</type>
<position>111,140.5</position>
<input>
<ID>N_in3</ID>202 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>GA_LED</type>
<position>119.5,140.5</position>
<input>
<ID>N_in3</ID>203 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>GA_LED</type>
<position>127,140.5</position>
<input>
<ID>N_in3</ID>204 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>GA_LED</type>
<position>133,140.5</position>
<input>
<ID>N_in3</ID>205 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>GA_LED</type>
<position>139.5,140.5</position>
<input>
<ID>N_in3</ID>206 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>GA_LED</type>
<position>145.5,140.5</position>
<input>
<ID>N_in3</ID>207 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>GA_LED</type>
<position>152.5,140.5</position>
<input>
<ID>N_in3</ID>208 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>GA_LED</type>
<position>158,140.5</position>
<input>
<ID>N_in3</ID>209 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>DE_TO</type>
<position>103,126.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>202</ID>
<type>DE_TO</type>
<position>104,119</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>203</ID>
<type>DE_TO</type>
<position>104,112</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>204</ID>
<type>DE_TO</type>
<position>114,103.5</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>205</ID>
<type>DE_TO</type>
<position>122,103.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>206</ID>
<type>DE_TO</type>
<position>129,103.5</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>207</ID>
<type>DE_TO</type>
<position>135,103.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>208</ID>
<type>DE_TO</type>
<position>141,104</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>209</ID>
<type>DE_TO</type>
<position>147,103.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>153,103.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_TO</type>
<position>160,103.5</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>111,151.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>119.5,151</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>214</ID>
<type>DA_FROM</type>
<position>127,151</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>215</ID>
<type>DA_FROM</type>
<position>133,151.5</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>139.5,151.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>145.5,151.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>152.5,151.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>158,151.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>109,164.5</position>
<gparam>LABEL_TEXT OUTPUT READ HERE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AE_DFF_LOW</type>
<position>330,166.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>164 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>222</ID>
<type>AE_DFF_LOW</type>
<position>352.5,166.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>159 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_DFF_LOW</type>
<position>376,166.5</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>158 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>224</ID>
<type>AE_DFF_LOW</type>
<position>395,166.5</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>149 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_DFF_LOW</type>
<position>417.5,166.5</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>148 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>226</ID>
<type>AE_DFF_LOW</type>
<position>439,166.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>139 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>227</ID>
<type>AE_DFF_LOW</type>
<position>460.5,166.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>131 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_DFF_LOW</type>
<position>480.5,166.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>129 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>229</ID>
<type>BA_TRI_STATE</type>
<position>337,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>164 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>230</ID>
<type>BA_TRI_STATE</type>
<position>360.5,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>BA_TRI_STATE</type>
<position>383,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>232</ID>
<type>BA_TRI_STATE</type>
<position>403.5,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>149 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>233</ID>
<type>BA_TRI_STATE</type>
<position>425,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>234</ID>
<type>BA_TRI_STATE</type>
<position>446.5,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>139 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>235</ID>
<type>BA_TRI_STATE</type>
<position>468,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>236</ID>
<type>BA_TRI_STATE</type>
<position>488,160.5</position>
<input>
<ID>ENABLE_0</ID>96 </input>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>237</ID>
<type>AE_DFF_LOW</type>
<position>330,151</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>165 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_DFF_LOW</type>
<position>352.5,151</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>160 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>239</ID>
<type>AE_DFF_LOW</type>
<position>376,151</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>157 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_DFF_LOW</type>
<position>395,151</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>150 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_DFF_LOW</type>
<position>417.5,151</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>147 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_DFF_LOW</type>
<position>439,151</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>140 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>243</ID>
<type>AE_DFF_LOW</type>
<position>460.5,151</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>132 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_DFF_LOW</type>
<position>480.5,151</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>130 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>245</ID>
<type>BA_TRI_STATE</type>
<position>337,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>246</ID>
<type>BA_TRI_STATE</type>
<position>360.5,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>247</ID>
<type>BA_TRI_STATE</type>
<position>383,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>248</ID>
<type>BA_TRI_STATE</type>
<position>403.5,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>249</ID>
<type>BA_TRI_STATE</type>
<position>425,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>147 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>250</ID>
<type>BA_TRI_STATE</type>
<position>446.5,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>140 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>251</ID>
<type>BA_TRI_STATE</type>
<position>468,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>252</ID>
<type>BA_TRI_STATE</type>
<position>488,145</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>253</ID>
<type>AE_DFF_LOW</type>
<position>330,134.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>168 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_DFF_LOW</type>
<position>352.5,134.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>161 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_DFF_LOW</type>
<position>376,134.5</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>156 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>256</ID>
<type>AE_DFF_LOW</type>
<position>395,134.5</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>151 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>257</ID>
<type>AE_DFF_LOW</type>
<position>417.5,134.5</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>146 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>258</ID>
<type>AE_DFF_LOW</type>
<position>439,134.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>141 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>259</ID>
<type>AE_DFF_LOW</type>
<position>460.5,134.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>136 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_DFF_LOW</type>
<position>480.5,134.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>135 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>261</ID>
<type>BA_TRI_STATE</type>
<position>337,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>262</ID>
<type>BA_TRI_STATE</type>
<position>360.5,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>263</ID>
<type>BA_TRI_STATE</type>
<position>383,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>264</ID>
<type>BA_TRI_STATE</type>
<position>403.5,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>151 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>265</ID>
<type>BA_TRI_STATE</type>
<position>425,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>146 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>266</ID>
<type>BA_TRI_STATE</type>
<position>446.5,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>141 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>267</ID>
<type>BA_TRI_STATE</type>
<position>468,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>136 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>268</ID>
<type>BA_TRI_STATE</type>
<position>488,128.5</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_DFF_LOW</type>
<position>330,118.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>167 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_DFF_LOW</type>
<position>352.5,118.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>162 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>271</ID>
<type>AE_DFF_LOW</type>
<position>376,118.5</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>155 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>272</ID>
<type>AE_DFF_LOW</type>
<position>395,118.5</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>152 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>273</ID>
<type>AE_DFF_LOW</type>
<position>417.5,118.5</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>145 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>274</ID>
<type>AE_DFF_LOW</type>
<position>439,118.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>142 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>275</ID>
<type>AE_DFF_LOW</type>
<position>460.5,118.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>137 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>276</ID>
<type>AE_DFF_LOW</type>
<position>480.5,118.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clock</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>277</ID>
<type>BA_TRI_STATE</type>
<position>337,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>278</ID>
<type>BA_TRI_STATE</type>
<position>360.5,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>162 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>279</ID>
<type>BA_TRI_STATE</type>
<position>383,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>280</ID>
<type>BA_TRI_STATE</type>
<position>403.5,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>281</ID>
<type>BA_TRI_STATE</type>
<position>425,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>145 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>282</ID>
<type>BA_TRI_STATE</type>
<position>446.5,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>283</ID>
<type>BA_TRI_STATE</type>
<position>468,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>137 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>284</ID>
<type>BA_TRI_STATE</type>
<position>488,112.5</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>285</ID>
<type>AE_DFF_LOW</type>
<position>330,102.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>166 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_DFF_LOW</type>
<position>352.5,102.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>163 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>287</ID>
<type>AE_DFF_LOW</type>
<position>376,102.5</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>154 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_DFF_LOW</type>
<position>395,102.5</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>153 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_DFF_LOW</type>
<position>417.5,102.5</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>144 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_DFF_LOW</type>
<position>439,102.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>143 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_DFF_LOW</type>
<position>460.5,102.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>138 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_DFF_LOW</type>
<position>480.5,102.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>133 </output>
<input>
<ID>clock</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>293</ID>
<type>BA_TRI_STATE</type>
<position>337,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>166 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>294</ID>
<type>BA_TRI_STATE</type>
<position>360.5,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>295</ID>
<type>BA_TRI_STATE</type>
<position>383,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>296</ID>
<type>BA_TRI_STATE</type>
<position>403.5,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>297</ID>
<type>BA_TRI_STATE</type>
<position>425,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>298</ID>
<type>BA_TRI_STATE</type>
<position>446.5,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>143 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>299</ID>
<type>BA_TRI_STATE</type>
<position>468,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>138 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>300</ID>
<type>BA_TRI_STATE</type>
<position>488,96.5</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>301</ID>
<type>AE_DFF_LOW</type>
<position>330,86.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>169 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_DFF_LOW</type>
<position>352.5,86.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>172 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_DFF_LOW</type>
<position>376,86.5</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>173 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_DFF_LOW</type>
<position>395,86.5</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>176 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>305</ID>
<type>AE_DFF_LOW</type>
<position>417.5,86.5</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>181 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>439,86.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>182 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_DFF_LOW</type>
<position>460.5,86.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>186 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_DFF_LOW</type>
<position>480.5,86.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>188 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>309</ID>
<type>BA_TRI_STATE</type>
<position>337,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>310</ID>
<type>BA_TRI_STATE</type>
<position>360.5,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>311</ID>
<type>BA_TRI_STATE</type>
<position>383,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>173 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>312</ID>
<type>BA_TRI_STATE</type>
<position>403.5,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>176 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>313</ID>
<type>BA_TRI_STATE</type>
<position>425,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>181 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>314</ID>
<type>BA_TRI_STATE</type>
<position>446.5,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>315</ID>
<type>BA_TRI_STATE</type>
<position>468,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>186 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>316</ID>
<type>BA_TRI_STATE</type>
<position>488,80.5</position>
<input>
<ID>ENABLE_0</ID>106 </input>
<input>
<ID>IN_0</ID>188 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>317</ID>
<type>AE_DFF_LOW</type>
<position>330,71.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>111 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_DFF_LOW</type>
<position>352.5,71.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>171 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_DFF_LOW</type>
<position>376,71.5</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>175 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_DFF_LOW</type>
<position>395,71.5</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>178 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>321</ID>
<type>AE_DFF_LOW</type>
<position>417.5,71.5</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>179 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_DFF_LOW</type>
<position>439,71.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>183 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_DFF_LOW</type>
<position>460.5,71.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>185 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_DFF_LOW</type>
<position>480.5,71.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>189 </output>
<input>
<ID>clock</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>325</ID>
<type>BA_TRI_STATE</type>
<position>337,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>111 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>326</ID>
<type>BA_TRI_STATE</type>
<position>360.5,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>171 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>327</ID>
<type>BA_TRI_STATE</type>
<position>383,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>175 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>328</ID>
<type>BA_TRI_STATE</type>
<position>403.5,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>178 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>329</ID>
<type>BA_TRI_STATE</type>
<position>425,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>330</ID>
<type>BA_TRI_STATE</type>
<position>446.5,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>183 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>331</ID>
<type>BA_TRI_STATE</type>
<position>468,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>185 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>332</ID>
<type>BA_TRI_STATE</type>
<position>488,65.5</position>
<input>
<ID>ENABLE_0</ID>110 </input>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>333</ID>
<type>AE_DFF_LOW</type>
<position>330,56</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>112 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>334</ID>
<type>AE_DFF_LOW</type>
<position>352.5,56</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>170 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_DFF_LOW</type>
<position>376,56</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>174 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_DFF_LOW</type>
<position>395,56</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>177 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_DFF_LOW</type>
<position>417.5,56</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>180 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_DFF_LOW</type>
<position>439,56</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>184 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>339</ID>
<type>AE_DFF_LOW</type>
<position>460.5,56</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>187 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>340</ID>
<type>AE_DFF_LOW</type>
<position>480.5,56</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>190 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>341</ID>
<type>BA_TRI_STATE</type>
<position>337,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>342</ID>
<type>BA_TRI_STATE</type>
<position>360.5,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>343</ID>
<type>BA_TRI_STATE</type>
<position>383,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>174 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>BA_TRI_STATE</type>
<position>403.5,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>345</ID>
<type>BA_TRI_STATE</type>
<position>425,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>346</ID>
<type>BA_TRI_STATE</type>
<position>446.5,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>184 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>347</ID>
<type>BA_TRI_STATE</type>
<position>468,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>348</ID>
<type>BA_TRI_STATE</type>
<position>488,50</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_AND2</type>
<position>295.5,165.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_AND2</type>
<position>304,160.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_AND2</type>
<position>295.5,150</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND2</type>
<position>304,145</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_AND2</type>
<position>295.5,133.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>304,128.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>295.5,117.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_AND2</type>
<position>304,112.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_AND2</type>
<position>295.5,101.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AI_XOR2</type>
<position>658,168</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AI_XOR2</type>
<position>672,162.5</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_AND2</type>
<position>672,153</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AI_XOR2</type>
<position>616.5,162.5</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>237 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>AE_OR2</type>
<position>682,149.5</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>616.5,153</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_OR2</type>
<position>626.5,149.5</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>GA_LED</type>
<position>623.5,162.5</position>
<input>
<ID>N_in0</ID>239 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>GA_LED</type>
<position>679,162.5</position>
<input>
<ID>N_in0</ID>217 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>369</ID>
<type>AA_AND2</type>
<position>597.5,148.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_LABEL</type>
<position>633,147</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>AA_LABEL</type>
<position>625.5,160.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>HA_JUNC_2</type>
<position>585,149.5</position>
<input>
<ID>N_in0</ID>243 </input>
<input>
<ID>N_in1</ID>237 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>374</ID>
<type>AI_XOR2</type>
<position>882.5,167.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>246 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>AI_XOR2</type>
<position>896.5,162</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>245 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND2</type>
<position>653,148.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_AND2</type>
<position>896.5,152.5</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AI_XOR2</type>
<position>841,162</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_LABEL</type>
<position>688.5,147</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>381</ID>
<type>AE_OR2</type>
<position>906.5,149</position>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_AND2</type>
<position>841,152.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>269 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_LABEL</type>
<position>681,160.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>384</ID>
<type>AE_OR2</type>
<position>851,149</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>AI_XOR2</type>
<position>713,168</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>226 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>386</ID>
<type>GA_LED</type>
<position>848,162</position>
<input>
<ID>N_in0</ID>270 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>387</ID>
<type>AI_XOR2</type>
<position>727,162.5</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_AND2</type>
<position>727,153</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,133,102.5,133</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,121,236.5,166.5</points>
<intersection>121 2</intersection>
<intersection>166.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,166.5,292.5,166.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>236.5 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,121,236.5,121</points>
<connection>
<GID>122</GID>
<name>OUT_7</name></connection>
<intersection>236.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,161.5,288,166.5</points>
<intersection>161.5 4</intersection>
<intersection>166.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,161.5,301,161.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,120,238.5,151</points>
<intersection>120 2</intersection>
<intersection>151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,151,292.5,151</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,120,238.5,120</points>
<connection>
<GID>122</GID>
<name>OUT_6</name></connection>
<intersection>238.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,146,288,151</points>
<intersection>146 4</intersection>
<intersection>151 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,146,301,146</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,119,241.5,134.5</points>
<intersection>119 2</intersection>
<intersection>134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241.5,134.5,292.5,134.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,119,241.5,119</points>
<connection>
<GID>122</GID>
<name>OUT_5</name></connection>
<intersection>241.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,129.5,288,134.5</points>
<intersection>129.5 4</intersection>
<intersection>134.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,129.5,301,129.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225.5,118.5,292.5,118.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>225.5 6</intersection>
<intersection>288 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,113.5,288,118.5</points>
<intersection>113.5 4</intersection>
<intersection>118.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,113.5,301,113.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>225.5,118,225.5,118.5</points>
<connection>
<GID>122</GID>
<name>OUT_4</name></connection>
<intersection>118.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,102.5,242,117</points>
<intersection>102.5 1</intersection>
<intersection>117 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242,102.5,292.5,102.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>242 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,117,242,117</points>
<connection>
<GID>122</GID>
<name>OUT_3</name></connection>
<intersection>242 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,97.5,288,102.5</points>
<intersection>97.5 4</intersection>
<intersection>102.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,97.5,301,97.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,86.5,238.5,116</points>
<intersection>86.5 1</intersection>
<intersection>116 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,86.5,292.5,86.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>238.5 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,116,238.5,116</points>
<connection>
<GID>122</GID>
<name>OUT_2</name></connection>
<intersection>238.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,81.5,288,86.5</points>
<intersection>81.5 4</intersection>
<intersection>86.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,81.5,300.5,81.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,71.5,236,115</points>
<intersection>71.5 1</intersection>
<intersection>115 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,71.5,292.5,71.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>236 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,115,236,115</points>
<connection>
<GID>122</GID>
<name>OUT_1</name></connection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,66.5,288,71.5</points>
<intersection>66.5 4</intersection>
<intersection>71.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,66.5,301,66.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,56,232.5,114</points>
<intersection>56 1</intersection>
<intersection>114 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,56,292.5,56</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>232.5 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,114,232.5,114</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,51,288,56</points>
<intersection>51 4</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,51,301,51</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,26.5,323,30.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346.5,26.5,346.5,30.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,27.5,369,30.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389.5,26.5,389.5,30.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411,27,411,30.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,26.5,432.5,30.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,27,454,30.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>474,28,474,30.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307.5,33.5,472,33.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>143</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>142</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>140</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>139</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>137</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>136</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>134</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>133</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342.5,193.5,342.5,203</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>203 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>340,203,342.5,203</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>342.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366,193.5,366,203</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>203 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>363,203,366,203</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>366 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387.5,193.5,387.5,203</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>203 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>386,203,387.5,203</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>387.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,193.5,408.5,203.5</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>203.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>406.5,203.5,408.5,203.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,193.5,430,203.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>203.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>428,203.5,430,203.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>430 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451.5,193.5,451.5,204</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>204 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>449.5,204,451.5,204</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>451.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>472,193.5,472,203.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>203.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>471,203.5,472,203.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>472 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496.5,193.5,496.5,203</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>203 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>491,203,496.5,203</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>323,191,494.5,191</points>
<connection>
<GID>157</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>156</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>154</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>152</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>150</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>148</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>146</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>145</GID>
<name>ENABLE_0</name></connection>
<intersection>323 34</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>323,190.5,323,191</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>191 1</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,34,279,164.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>54 8</intersection>
<intersection>69.5 7</intersection>
<intersection>84.5 6</intersection>
<intersection>100.5 5</intersection>
<intersection>116.5 4</intersection>
<intersection>132.5 3</intersection>
<intersection>149 2</intersection>
<intersection>164.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,164.5,292.5,164.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>279,149,292.5,149</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>279,132.5,292.5,132.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279,116.5,292.5,116.5</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>279,100.5,292.5,100.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>279,84.5,292.5,84.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>279,69.5,292.5,69.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>279,54,292.5,54</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,49,284,188</points>
<intersection>49 1</intersection>
<intersection>64.5 3</intersection>
<intersection>79.5 5</intersection>
<intersection>95.5 7</intersection>
<intersection>111.5 9</intersection>
<intersection>127.5 10</intersection>
<intersection>144 11</intersection>
<intersection>159.5 12</intersection>
<intersection>188 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284,49,301,49</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>284,64.5,301,64.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>284,79.5,300.5,79.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>284,95.5,301,95.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>282,188,284,188</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>284,111.5,301,111.5</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>284,127.5,301,127.5</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>284,144,301,144</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>284,159.5,301,159.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,165.5,477.5,165.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<connection>
<GID>228</GID>
<name>clock</name></connection>
<connection>
<GID>227</GID>
<name>clock</name></connection>
<connection>
<GID>226</GID>
<name>clock</name></connection>
<connection>
<GID>225</GID>
<name>clock</name></connection>
<connection>
<GID>224</GID>
<name>clock</name></connection>
<connection>
<GID>223</GID>
<name>clock</name></connection>
<connection>
<GID>222</GID>
<name>clock</name></connection>
<connection>
<GID>221</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,160.5,486,160.5</points>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<connection>
<GID>236</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>235</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>234</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>233</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>232</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>231</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>230</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>229</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,145,486,145</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<connection>
<GID>252</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>251</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>250</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>249</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>248</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>247</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>246</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>245</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,150,477.5,150</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<connection>
<GID>244</GID>
<name>clock</name></connection>
<connection>
<GID>243</GID>
<name>clock</name></connection>
<connection>
<GID>242</GID>
<name>clock</name></connection>
<connection>
<GID>241</GID>
<name>clock</name></connection>
<connection>
<GID>240</GID>
<name>clock</name></connection>
<connection>
<GID>239</GID>
<name>clock</name></connection>
<connection>
<GID>238</GID>
<name>clock</name></connection>
<connection>
<GID>237</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,133.5,477.5,133.5</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<connection>
<GID>260</GID>
<name>clock</name></connection>
<connection>
<GID>259</GID>
<name>clock</name></connection>
<connection>
<GID>258</GID>
<name>clock</name></connection>
<connection>
<GID>257</GID>
<name>clock</name></connection>
<connection>
<GID>256</GID>
<name>clock</name></connection>
<connection>
<GID>255</GID>
<name>clock</name></connection>
<connection>
<GID>254</GID>
<name>clock</name></connection>
<connection>
<GID>253</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,128.5,486,128.5</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<connection>
<GID>268</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>267</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>266</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>265</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>264</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>263</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>262</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>261</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,117.5,477.5,117.5</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<connection>
<GID>276</GID>
<name>clock</name></connection>
<connection>
<GID>275</GID>
<name>clock</name></connection>
<connection>
<GID>274</GID>
<name>clock</name></connection>
<connection>
<GID>273</GID>
<name>clock</name></connection>
<connection>
<GID>272</GID>
<name>clock</name></connection>
<connection>
<GID>271</GID>
<name>clock</name></connection>
<connection>
<GID>270</GID>
<name>clock</name></connection>
<connection>
<GID>269</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,112.5,486,112.5</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<connection>
<GID>284</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>283</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>282</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>281</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>280</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>279</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>278</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>277</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,101.5,477.5,101.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<connection>
<GID>292</GID>
<name>clock</name></connection>
<connection>
<GID>291</GID>
<name>clock</name></connection>
<connection>
<GID>290</GID>
<name>clock</name></connection>
<connection>
<GID>289</GID>
<name>clock</name></connection>
<connection>
<GID>288</GID>
<name>clock</name></connection>
<connection>
<GID>287</GID>
<name>clock</name></connection>
<connection>
<GID>286</GID>
<name>clock</name></connection>
<connection>
<GID>285</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>307,96.5,486,96.5</points>
<connection>
<GID>300</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>299</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>298</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>297</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>296</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>295</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>294</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>293</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>112</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,85.5,477.5,85.5</points>
<connection>
<GID>308</GID>
<name>clock</name></connection>
<connection>
<GID>307</GID>
<name>clock</name></connection>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<connection>
<GID>305</GID>
<name>clock</name></connection>
<connection>
<GID>304</GID>
<name>clock</name></connection>
<connection>
<GID>303</GID>
<name>clock</name></connection>
<connection>
<GID>302</GID>
<name>clock</name></connection>
<connection>
<GID>301</GID>
<name>clock</name></connection>
<connection>
<GID>113</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>306.5,80.5,486,80.5</points>
<connection>
<GID>316</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>315</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>314</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>313</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>312</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>311</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>310</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>309</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>114</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,70.5,477.5,70.5</points>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<connection>
<GID>323</GID>
<name>clock</name></connection>
<connection>
<GID>322</GID>
<name>clock</name></connection>
<connection>
<GID>321</GID>
<name>clock</name></connection>
<connection>
<GID>320</GID>
<name>clock</name></connection>
<connection>
<GID>319</GID>
<name>clock</name></connection>
<connection>
<GID>318</GID>
<name>clock</name></connection>
<connection>
<GID>317</GID>
<name>clock</name></connection>
<connection>
<GID>116</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,55,477.5,55</points>
<connection>
<GID>340</GID>
<name>clock</name></connection>
<connection>
<GID>339</GID>
<name>clock</name></connection>
<connection>
<GID>338</GID>
<name>clock</name></connection>
<connection>
<GID>337</GID>
<name>clock</name></connection>
<connection>
<GID>336</GID>
<name>clock</name></connection>
<connection>
<GID>335</GID>
<name>clock</name></connection>
<connection>
<GID>334</GID>
<name>clock</name></connection>
<connection>
<GID>333</GID>
<name>clock</name></connection>
<connection>
<GID>119</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,50,486,50</points>
<connection>
<GID>348</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>347</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>346</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>345</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>344</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>343</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>342</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>341</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,65.5,486,65.5</points>
<connection>
<GID>332</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>331</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>330</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>329</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>328</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>327</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>326</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>325</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,62.5,333.5,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,73.5,333.5,73.5</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>333.5,62.5,337,62.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,47,334,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,58,334,58</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>334,47,337,47</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,36,323,168.5</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>58 8</intersection>
<intersection>73.5 7</intersection>
<intersection>88.5 6</intersection>
<intersection>104.5 5</intersection>
<intersection>120.5 4</intersection>
<intersection>136.5 3</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,168.5,327,168.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>323,153,327,153</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>323,136.5,327,136.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>323,120.5,327,120.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>323,104.5,327,104.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>323,88.5,327,88.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>323,73.5,327,73.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>323,58,327,58</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>323 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342.5,52.5,342.5,188</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 12</intersection>
<intersection>83 6</intersection>
<intersection>99 7</intersection>
<intersection>115 8</intersection>
<intersection>131 9</intersection>
<intersection>147.5 10</intersection>
<intersection>163 11</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>337,52.5,342.5,52.5</points>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>337,83,342.5,83</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>337,99,342.5,99</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>337,115,342.5,115</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>337,131,342.5,131</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>337,147.5,342.5,147.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>337,163,342.5,163</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>337,68,342.5,68</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346.5,36,346.5,168.5</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>58 7</intersection>
<intersection>73.5 8</intersection>
<intersection>88.5 6</intersection>
<intersection>104.5 5</intersection>
<intersection>120.5 4</intersection>
<intersection>136.5 3</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>346.5,168.5,349.5,168.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346.5,153,349.5,153</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>346.5,136.5,349.5,136.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>346.5,120.5,349.5,120.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>346.5,104.5,349.5,104.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>346.5,88.5,349.5,88.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>346.5,58,349.5,58</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>346.5,73.5,349.5,73.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>346.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366,52.5,366,188</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 12</intersection>
<intersection>83 11</intersection>
<intersection>99 10</intersection>
<intersection>115 9</intersection>
<intersection>131 8</intersection>
<intersection>147.5 6</intersection>
<intersection>163 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>360.5,52.5,366,52.5</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>360.5,147.5,366,147.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>360.5,163,366,163</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>360.5,131,366,131</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>360.5,115,366,115</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>360.5,99,366,99</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>360.5,83,366,83</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>360.5,68,366,68</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>366 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,36,369,168.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>58 8</intersection>
<intersection>73.5 7</intersection>
<intersection>88.5 6</intersection>
<intersection>104.5 5</intersection>
<intersection>120.5 4</intersection>
<intersection>136.5 3</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369,168.5,373,168.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>369,153,373,153</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>369,136.5,373,136.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>369,120.5,373,120.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>369,104.5,373,104.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>369,88.5,373,88.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>369,73.5,373,73.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>369,58,373,58</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387.5,52.5,387.5,188</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 12</intersection>
<intersection>83 7</intersection>
<intersection>99 11</intersection>
<intersection>115 10</intersection>
<intersection>131 8</intersection>
<intersection>147.5 9</intersection>
<intersection>163 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>383,52.5,387.5,52.5</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>383,163,387.5,163</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>383,83,387.5,83</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>383,131,387.5,131</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>383,147.5,387.5,147.5</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>383,115,387.5,115</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>383,99,387.5,99</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>383,68,387.5,68</points>
<connection>
<GID>327</GID>
<name>OUT_0</name></connection>
<intersection>387.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389.5,36,389.5,168.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>58 8</intersection>
<intersection>73.5 7</intersection>
<intersection>88.5 6</intersection>
<intersection>104.5 5</intersection>
<intersection>120.5 4</intersection>
<intersection>136.5 2</intersection>
<intersection>153 3</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>389.5,168.5,392,168.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>389.5,136.5,392,136.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>389.5,153,392,153</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>389.5,120.5,392,120.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>389.5,104.5,392,104.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>389.5,88.5,392,88.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>389.5,73.5,392,73.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>389.5,58,392,58</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>389.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,52.5,408.5,188</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 12</intersection>
<intersection>83 8</intersection>
<intersection>99 10</intersection>
<intersection>115 11</intersection>
<intersection>131 9</intersection>
<intersection>147.5 6</intersection>
<intersection>163 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>403.5,52.5,408.5,52.5</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>403.5,147.5,408.5,147.5</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>403.5,163,408.5,163</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>403.5,83,408.5,83</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>403.5,131,408.5,131</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>403.5,99,408.5,99</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>403.5,115,408.5,115</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>403.5,68,408.5,68</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411,36,411,168.5</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>58 8</intersection>
<intersection>73.5 7</intersection>
<intersection>88.5 3</intersection>
<intersection>104.5 4</intersection>
<intersection>120.5 5</intersection>
<intersection>136.5 6</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>411,168.5,414.5,168.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>411,153,414.5,153</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>411,88.5,414.5,88.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>411,104.5,414.5,104.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>411,120.5,414.5,120.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411,136.5,414.5,136.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>411,73.5,414.5,73.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>411,58,414.5,58</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,52.5,430,188</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 12</intersection>
<intersection>83 11</intersection>
<intersection>99 10</intersection>
<intersection>115 9</intersection>
<intersection>131 8</intersection>
<intersection>147.5 7</intersection>
<intersection>163 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>425,52.5,430,52.5</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>425,163,430,163</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>425,147.5,430,147.5</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>425,131,430,131</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>425,115,430,115</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>425,99,430,99</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>425,83,430,83</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>425,68,430,68</points>
<connection>
<GID>329</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,36,432.5,168.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>58 8</intersection>
<intersection>73.5 7</intersection>
<intersection>88.5 3</intersection>
<intersection>104.5 4</intersection>
<intersection>120.5 5</intersection>
<intersection>136.5 6</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,168.5,436,168.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432.5,153,436,153</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432.5,88.5,436,88.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>432.5,104.5,436,104.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>432.5,120.5,436,120.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>432.5,136.5,436,136.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>432.5,73.5,436,73.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>432.5,58,436,58</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451.5,52.5,451.5,188</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 10</intersection>
<intersection>83 9</intersection>
<intersection>99 8</intersection>
<intersection>115 7</intersection>
<intersection>131 6</intersection>
<intersection>147.5 5</intersection>
<intersection>163 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>446.5,52.5,451.5,52.5</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>446.5,163,451.5,163</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>446.5,147.5,451.5,147.5</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>446.5,131,451.5,131</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>446.5,115,451.5,115</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>446.5,99,451.5,99</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>446.5,83,451.5,83</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>446.5,68,451.5,68</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>451.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,36,454,168.5</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>58 8</intersection>
<intersection>73.5 7</intersection>
<intersection>88.5 6</intersection>
<intersection>104.5 5</intersection>
<intersection>120.5 4</intersection>
<intersection>136.5 3</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454,168.5,457.5,168.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>454,153,457.5,153</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>454,136.5,457.5,136.5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>454,120.5,457.5,120.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>454,104.5,457.5,104.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>454,88.5,457.5,88.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>454,73.5,457.5,73.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>454,58,457.5,58</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>472,52.5,472,188</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>52.5 5</intersection>
<intersection>68 12</intersection>
<intersection>83 11</intersection>
<intersection>99 10</intersection>
<intersection>115 9</intersection>
<intersection>131 8</intersection>
<intersection>147.5 7</intersection>
<intersection>163 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>468,52.5,472,52.5</points>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>468,163,472,163</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>468,147.5,472,147.5</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>468,131,472,131</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>468,115,472,115</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>468,99,472,99</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>468,83,472,83</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>468,68,472,68</points>
<connection>
<GID>331</GID>
<name>OUT_0</name></connection>
<intersection>472 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>474,36,474,168.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>58 7</intersection>
<intersection>73.5 5</intersection>
<intersection>88.5 6</intersection>
<intersection>104.5 8</intersection>
<intersection>120.5 4</intersection>
<intersection>136.5 3</intersection>
<intersection>153 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>474,168.5,477.5,168.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>474,153,477.5,153</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>474,136.5,477.5,136.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>474,120.5,477.5,120.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>474,73.5,477.5,73.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474,88.5,477.5,88.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>474,58,477.5,58</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>474,104.5,477.5,104.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>474 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496.5,52.5,496.5,188</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>68 12</intersection>
<intersection>83 11</intersection>
<intersection>99 10</intersection>
<intersection>115 8</intersection>
<intersection>131 9</intersection>
<intersection>147.5 7</intersection>
<intersection>163 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>488,52.5,496.5,52.5</points>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>488,163,496.5,163</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>488,147.5,496.5,147.5</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>488,115,496.5,115</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>488,131,496.5,131</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>488,99,496.5,99</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>488,83,496.5,83</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>488,68,496.5,68</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485,157.5,485,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,168.5,485,168.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>485 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>485,157.5,488,157.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>485 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,142,484.5,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,153,484.5,153</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>484.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,142,488,142</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464,157.5,464,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,168.5,464,168.5</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,157.5,468,157.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464,142,464,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,153,464,153</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,142,468,142</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484,93.5,484,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,104.5,484,104.5</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>484 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484,93.5,488,93.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>484 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,109.5,484.5,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,120.5,484.5,120.5</points>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection>
<intersection>484.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,109.5,488,109.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,125.5,484.5,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,136.5,484.5,136.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>484.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,125.5,488,125.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,125.5,464.5,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,136.5,464.5,136.5</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464.5,125.5,468,125.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,109.5,464.5,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,120.5,464.5,120.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464.5,109.5,468,109.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464,93.5,464,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,104.5,464,104.5</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,93.5,468,93.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,157.5,443,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,168.5,443,168.5</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443,157.5,446.5,157.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>443 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,142,443,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,153,443,153</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443,142,446.5,142</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>443 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443.5,125.5,443.5,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,136.5,443.5,136.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443.5,125.5,446.5,125.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>443.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,109.5,444,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,120.5,444,120.5</points>
<connection>
<GID>274</GID>
<name>OUT_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,109.5,446.5,109.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,93.5,443,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,104.5,443,104.5</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443,93.5,446.5,93.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>443 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422,93.5,422,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>422,93.5,425,93.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>422 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>420.5,104.5,422,104.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>422 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,109.5,421.5,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,120.5,421.5,120.5</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,109.5,425,109.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,125.5,421.5,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,136.5,421.5,136.5</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,125.5,425,125.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,142,421.5,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,153,421.5,153</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,142,425,142</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422,157.5,422,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,168.5,422,168.5</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>422 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422,157.5,425,157.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>422 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,157.5,400.5,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,168.5,400.5,168.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400.5,157.5,403.5,157.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,142,400,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,153,400,153</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400,142,403.5,142</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>400 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,125.5,400,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,136.5,400,136.5</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400,125.5,403.5,125.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>400 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,109.5,400,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,120.5,400,120.5</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400,109.5,403.5,109.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>400 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,93.5,400,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,104.5,400,104.5</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400,93.5,403.5,93.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>400 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,93.5,379.5,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,104.5,379.5,104.5</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>379.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>379.5,93.5,383,93.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,109.5,379,120.5</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>109.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>379,109.5,383,109.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,125.5,380,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,136.5,380,136.5</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>380,125.5,383,125.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,142,379.5,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,153,379.5,153</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>379.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>379.5,142,383,142</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,157.5,380,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,168.5,380,168.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>380,157.5,383,157.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,157.5,356.5,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,168.5,356.5,168.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,157.5,360.5,157.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,142,356.5,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,153,356.5,153</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,142,360.5,142</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,125.5,357,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,136.5,357,136.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,125.5,360.5,125.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,109.5,356.5,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,120.5,356.5,120.5</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,109.5,360.5,109.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,93.5,356.5,104.5</points>
<intersection>93.5 2</intersection>
<intersection>104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,104.5,356.5,104.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,93.5,360.5,93.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,157.5,334,168.5</points>
<intersection>157.5 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,168.5,334,168.5</points>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>334,157.5,337,157.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,142,334.5,153</points>
<intersection>142 2</intersection>
<intersection>153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,153,334.5,153</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>334.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>334.5,142,337,142</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>334.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,93.5,333,104.5</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>333,93.5,337,93.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>333 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,109.5,333.5,120.5</points>
<intersection>109.5 2</intersection>
<intersection>120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,120.5,333.5,120.5</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>333.5,109.5,337,109.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,125.5,333.5,136.5</points>
<intersection>125.5 2</intersection>
<intersection>136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,136.5,333.5,136.5</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>333.5,125.5,337,125.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,77.5,334,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333,88.5,334,88.5</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>334,77.5,337,77.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,47,356.5,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,58,356.5,58</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,47,360.5,47</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,62.5,356,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,73.5,356,73.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356,62.5,360.5,62.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,77.5,356.5,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,88.5,356.5,88.5</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,77.5,360.5,77.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,77.5,380,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,88.5,380,88.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>380,77.5,383,77.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,47,380,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,58,380,58</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>380,47,383,47</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,62.5,379,73.5</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>379,62.5,383,62.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,77.5,399.5,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,88.5,399.5,88.5</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399.5,77.5,403.5,77.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>399.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,47,399,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,58,399,58</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>399 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399,47,403.5,47</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>399 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,62.5,399.5,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,73.5,399.5,73.5</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399.5,62.5,403.5,62.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>399.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,62.5,421.5,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,73.5,421.5,73.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,62.5,425,62.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,47,421.5,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,58,421.5,58</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,47,425,47</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,77.5,421.5,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,88.5,421.5,88.5</points>
<connection>
<GID>305</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,77.5,425,77.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442.5,77.5,442.5,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,88.5,442.5,88.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>442.5,77.5,446.5,77.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,62.5,443,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,73.5,443,73.5</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443,62.5,446.5,62.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>443 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442.5,47,442.5,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,58,442.5,58</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>442.5,47,446.5,47</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,62.5,465,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,73.5,465,73.5</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>465,62.5,468,62.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>465 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,77.5,464.5,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,88.5,464.5,88.5</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464.5,77.5,468,77.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,47,465,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,58,465,58</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>465,47,468,47</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>465 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,77.5,484.5,88.5</points>
<intersection>77.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,88.5,484.5,88.5</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<intersection>484.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,77.5,488,77.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,62.5,484.5,73.5</points>
<intersection>62.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,73.5,484.5,73.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>484.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,62.5,488,62.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,47,484.5,58</points>
<intersection>47 2</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,58,484.5,58</points>
<connection>
<GID>340</GID>
<name>OUT_0</name></connection>
<intersection>484.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,47,488,47</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,126.5,101,126.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,119,102,119</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>102 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>102,119,102,119</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>119 1</intersection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,113.5,102,113.5</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>102 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>102,112,102,113.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>113.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,96,114,101.5</points>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection>
<connection>
<GID>204</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,96,122,101.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,96.5,129,101.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,97,135,101.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,96,141,102</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,96,147.5,101.5</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>101.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>147,101.5,147.5,101.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,96.5,153,101.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,96.5,160,101.5</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>101.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>160,101.5,160,101.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,141.5,111,149.5</points>
<connection>
<GID>193</GID>
<name>N_in3</name></connection>
<connection>
<GID>212</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,141.5,119.5,149</points>
<connection>
<GID>194</GID>
<name>N_in3</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,141.5,127,149</points>
<connection>
<GID>195</GID>
<name>N_in3</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,141.5,133,149.5</points>
<connection>
<GID>196</GID>
<name>N_in3</name></connection>
<connection>
<GID>215</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,141.5,139.5,149.5</points>
<connection>
<GID>197</GID>
<name>N_in3</name></connection>
<connection>
<GID>216</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,141.5,145.5,149.5</points>
<connection>
<GID>198</GID>
<name>N_in3</name></connection>
<connection>
<GID>217</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,141.5,152.5,149.5</points>
<connection>
<GID>199</GID>
<name>N_in3</name></connection>
<connection>
<GID>218</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,141.5,158,149.5</points>
<connection>
<GID>200</GID>
<name>N_in3</name></connection>
<connection>
<GID>219</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,121,219.5,121</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<connection>
<GID>122</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,116.5,219.5,116.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>219.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>219.5,116,219.5,116.5</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>116.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,112,212,115</points>
<intersection>112 2</intersection>
<intersection>115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212,115,219.5,115</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,112,212,112</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,109,213.5,114</points>
<intersection>109 2</intersection>
<intersection>114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,114,219.5,114</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,109,213.5,109</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>677,150.5,677,153</points>
<intersection>150.5 1</intersection>
<intersection>153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>677,150.5,679,150.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>677 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>675,153,677,153</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>677 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>668,161.5,669,161.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>668 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>668,154,668,161.5</points>
<intersection>154 4</intersection>
<intersection>161.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>641,154,669,154</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>641 10</intersection>
<intersection>668 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>641,149.5,641,154</points>
<connection>
<GID>444</GID>
<name>N_in1</name></connection>
<intersection>154 4</intersection></vsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,168,665.5,168</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>665.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>665.5,152,665.5,168</points>
<intersection>152 5</intersection>
<intersection>163.5 6</intersection>
<intersection>168 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>665.5,152,669,152</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>665.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>665.5,163.5,669,163.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>665.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>675,162.5,678,162.5</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<connection>
<GID>368</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>634.5,172,650,172</points>
<intersection>634.5 8</intersection>
<intersection>650 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>650,149.5,650,172</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>169 6</intersection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>650,169,655,169</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>650 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>634.5,172,634.5,178.5</points>
<connection>
<GID>472</GID>
<name>OUT_0</name></connection>
<intersection>172 1</intersection></vsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>624.5,167,655,167</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<intersection>624.5 7</intersection>
<intersection>645 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>645,147.5,645,167</points>
<intersection>147.5 4</intersection>
<intersection>167 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>645,147.5,650,147.5</points>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>645 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>624.5,167,624.5,178.5</points>
<connection>
<GID>471</GID>
<name>OUT_0</name></connection>
<intersection>167 2</intersection></vsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>656,148.5,679,148.5</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<connection>
<GID>362</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>732,150.5,732,153</points>
<intersection>150.5 1</intersection>
<intersection>153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>732,150.5,734,150.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>732 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>730,153,732,153</points>
<connection>
<GID>388</GID>
<name>OUT</name></connection>
<intersection>732 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>723,161.5,724,161.5</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>723 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>723,154,723,161.5</points>
<intersection>154 4</intersection>
<intersection>161.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>696.5,154,724,154</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>696.5 7</intersection>
<intersection>723 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>696.5,149.5,696.5,154</points>
<connection>
<GID>412</GID>
<name>N_in1</name></connection>
<intersection>154 4</intersection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,168,720.5,168</points>
<connection>
<GID>385</GID>
<name>OUT</name></connection>
<intersection>720.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>720.5,152,720.5,168</points>
<intersection>152 5</intersection>
<intersection>163.5 6</intersection>
<intersection>168 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>720.5,152,724,152</points>
<connection>
<GID>388</GID>
<name>IN_1</name></connection>
<intersection>720.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>720.5,163.5,724,163.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>720.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>730,162.5,733,162.5</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<connection>
<GID>391</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,172,705,172</points>
<intersection>688 8</intersection>
<intersection>705 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>705,149.5,705,172</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>169 6</intersection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>705,169,710,169</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>705 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>688,172,688,177.5</points>
<connection>
<GID>475</GID>
<name>OUT_0</name></connection>
<intersection>172 1</intersection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>678,167,710,167</points>
<connection>
<GID>385</GID>
<name>IN_1</name></connection>
<intersection>678 7</intersection>
<intersection>699.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>699.5,147.5,699.5,167</points>
<intersection>147.5 4</intersection>
<intersection>167 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>699.5,147.5,705,147.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>699.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>678,167,678,177.5</points>
<connection>
<GID>474</GID>
<name>OUT_0</name></connection>
<intersection>167 2</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>711,148.5,734,148.5</points>
<connection>
<GID>397</GID>
<name>OUT</name></connection>
<connection>
<GID>389</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>685,149.5,694.5,149.5</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<connection>
<GID>412</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>566.5,150.5,566.5,153</points>
<intersection>150.5 1</intersection>
<intersection>153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>566.5,150.5,568.5,150.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>566.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>564.5,153,566.5,153</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>566.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557.5,161.5,558.5,161.5</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>557.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>557.5,154,557.5,161.5</points>
<intersection>154 4</intersection>
<intersection>161.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>530.5,154,558.5,154</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<intersection>557.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>550.5,168,555,168</points>
<connection>
<GID>414</GID>
<name>OUT</name></connection>
<intersection>555 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>555,152,555,168</points>
<intersection>152 5</intersection>
<intersection>163.5 6</intersection>
<intersection>168 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>555,152,558.5,152</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<intersection>555 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>555,163.5,558.5,163.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>555 3</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>564.5,162.5,567.5,162.5</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<connection>
<GID>422</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522.5,172,539.5,172</points>
<intersection>522.5 8</intersection>
<intersection>539.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>539.5,149.5,539.5,172</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>169 6</intersection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>539.5,169,544.5,169</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>539.5 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>522.5,172,522.5,178.5</points>
<connection>
<GID>457</GID>
<name>OUT_0</name></connection>
<intersection>172 1</intersection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>512.5,167,544.5,167</points>
<connection>
<GID>414</GID>
<name>IN_1</name></connection>
<intersection>512.5 7</intersection>
<intersection>534 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>534,147.5,534,167</points>
<intersection>147.5 4</intersection>
<intersection>167 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>534,147.5,539.5,147.5</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>534 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>512.5,167,512.5,178.5</points>
<connection>
<GID>456</GID>
<name>OUT_0</name></connection>
<intersection>167 2</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>545.5,148.5,568.5,148.5</points>
<connection>
<GID>428</GID>
<name>OUT</name></connection>
<connection>
<GID>420</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621.5,150.5,621.5,153</points>
<intersection>150.5 1</intersection>
<intersection>153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>621.5,150.5,623.5,150.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>621.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>619.5,153,621.5,153</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>621.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612.5,161.5,613.5,161.5</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<intersection>612.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>612.5,154,612.5,161.5</points>
<intersection>154 4</intersection>
<intersection>161.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>586,154,613.5,154</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>586 7</intersection>
<intersection>612.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>586,149.5,586,154</points>
<connection>
<GID>372</GID>
<name>N_in1</name></connection>
<intersection>154 4</intersection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>605.5,168,610,168</points>
<connection>
<GID>437</GID>
<name>OUT</name></connection>
<intersection>610 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>610,152,610,168</points>
<intersection>152 5</intersection>
<intersection>163.5 6</intersection>
<intersection>168 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>610,152,613.5,152</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>610 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>610,163.5,613.5,163.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>610 3</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,162.5,622.5,162.5</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<connection>
<GID>365</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578,172,594.5,172</points>
<intersection>578 8</intersection>
<intersection>594.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>594.5,149.5,594.5,172</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>169 6</intersection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>594.5,169,599.5,169</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>594.5 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>578,172,578,178.5</points>
<connection>
<GID>469</GID>
<name>OUT_0</name></connection>
<intersection>172 1</intersection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>568,167,599.5,167</points>
<connection>
<GID>437</GID>
<name>IN_1</name></connection>
<intersection>568 7</intersection>
<intersection>590.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>590.5,147.5,590.5,167</points>
<intersection>147.5 4</intersection>
<intersection>167 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>590.5,147.5,594.5,147.5</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>590.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>568,167,568,178.5</points>
<connection>
<GID>468</GID>
<name>OUT_0</name></connection>
<intersection>167 2</intersection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,148.5,623.5,148.5</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<connection>
<GID>364</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,149.5,584,149.5</points>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<connection>
<GID>372</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>901.5,150,901.5,152.5</points>
<intersection>150 1</intersection>
<intersection>152.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>901.5,150,903.5,150</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>901.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>899.5,152.5,901.5,152.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>901.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>892.5,161,893.5,161</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<intersection>892.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>892.5,153.5,892.5,161</points>
<intersection>153.5 4</intersection>
<intersection>161 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>865.5,153.5,893.5,153.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>865.5 7</intersection>
<intersection>892.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>865.5,149,865.5,153.5</points>
<intersection>149 8</intersection>
<intersection>153.5 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>864,149,865.5,149</points>
<connection>
<GID>446</GID>
<name>N_in1</name></connection>
<intersection>865.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>885.5,167.5,890,167.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>890 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>890,151.5,890,167.5</points>
<intersection>151.5 5</intersection>
<intersection>163 6</intersection>
<intersection>167.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>890,151.5,893.5,151.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>890 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>890,163,893.5,163</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>890 3</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>899.5,162,902.5,162</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<connection>
<GID>393</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>857.5,171.5,874.5,171.5</points>
<intersection>857.5 8</intersection>
<intersection>874.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>874.5,149,874.5,171.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>168.5 6</intersection>
<intersection>171.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>874.5,168.5,879.5,168.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>874.5 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>857.5,171.5,857.5,176</points>
<connection>
<GID>484</GID>
<name>OUT_0</name></connection>
<intersection>171.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>847.5,166.5,879.5,166.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>847.5 7</intersection>
<intersection>869 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>869,147,869,166.5</points>
<intersection>147 4</intersection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>869,147,874.5,147</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>869 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>847.5,166.5,847.5,176</points>
<connection>
<GID>483</GID>
<name>OUT_0</name></connection>
<intersection>166.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>880.5,148,903.5,148</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<connection>
<GID>381</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>956.5,150,956.5,152.5</points>
<intersection>150 1</intersection>
<intersection>152.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>956.5,150,958.5,150</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>956.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>954.5,152.5,956.5,152.5</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>956.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>947.5,161,948.5,161</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>947.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>947.5,153.5,947.5,161</points>
<intersection>153.5 4</intersection>
<intersection>161 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>921,153.5,948.5,153.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>921 7</intersection>
<intersection>947.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>921,149,921,153.5</points>
<connection>
<GID>427</GID>
<name>N_in1</name></connection>
<intersection>153.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>940.5,167.5,945,167.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>945 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>945,151.5,945,167.5</points>
<intersection>151.5 5</intersection>
<intersection>163 6</intersection>
<intersection>167.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>945,151.5,948.5,151.5</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>945 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>945,163,948.5,163</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>945 3</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>954.5,162,957.5,162</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<connection>
<GID>413</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>964.5,149,966.5,149</points>
<connection>
<GID>411</GID>
<name>OUT</name></connection>
<connection>
<GID>415</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>912.5,171.5,929.5,171.5</points>
<intersection>912.5 8</intersection>
<intersection>929.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>929.5,149,929.5,171.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>168.5 6</intersection>
<intersection>171.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>929.5,168.5,934.5,168.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>929.5 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>912.5,171.5,912.5,175.5</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<intersection>171.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>902.5,166.5,934.5,166.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>902.5 7</intersection>
<intersection>924.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>924.5,147,924.5,166.5</points>
<intersection>147 4</intersection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>924.5,147,929.5,147</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>924.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>902.5,166.5,902.5,175.5</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>166.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>935.5,148,958.5,148</points>
<connection>
<GID>421</GID>
<name>OUT</name></connection>
<connection>
<GID>411</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>909.5,149,919,149</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<connection>
<GID>427</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>791,150,791,152.5</points>
<intersection>150 1</intersection>
<intersection>152.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>791,150,793,150</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>791 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>789,152.5,791,152.5</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<intersection>791 0</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>782,161,783,161</points>
<connection>
<GID>431</GID>
<name>IN_1</name></connection>
<intersection>782 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>782,153.5,782,161</points>
<intersection>153.5 4</intersection>
<intersection>161 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>749.5,153.5,783,153.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>749.5 7</intersection>
<intersection>782 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>749.5,149.5,749.5,153.5</points>
<connection>
<GID>445</GID>
<name>N_in1</name></connection>
<intersection>153.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>775,167.5,779.5,167.5</points>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<intersection>779.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>779.5,151.5,779.5,167.5</points>
<intersection>151.5 5</intersection>
<intersection>163 6</intersection>
<intersection>167.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>779.5,151.5,783,151.5</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>779.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>779.5,163,783,163</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>779.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>789,162,792,162</points>
<connection>
<GID>431</GID>
<name>OUT</name></connection>
<connection>
<GID>436</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>748,171.5,764,171.5</points>
<intersection>748 8</intersection>
<intersection>764 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>764,149,764,171.5</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>168.5 6</intersection>
<intersection>171.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>764,168.5,769,168.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>764 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>748,171.5,748,177.5</points>
<connection>
<GID>478</GID>
<name>OUT_0</name></connection>
<intersection>171.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>738,166.5,769,166.5</points>
<connection>
<GID>429</GID>
<name>IN_1</name></connection>
<intersection>738 7</intersection>
<intersection>758.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>758.5,147,758.5,166.5</points>
<intersection>147 4</intersection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>758.5,147,764,147</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<intersection>758.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>738,166.5,738,177.5</points>
<connection>
<GID>477</GID>
<name>OUT_0</name></connection>
<intersection>166.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>770,148,793,148</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<connection>
<GID>435</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>846,150,846,152.5</points>
<intersection>150 1</intersection>
<intersection>152.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>846,150,848,150</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>846 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>844,152.5,846,152.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>846 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>837,161,838,161</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<intersection>837 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>837,153.5,837,161</points>
<intersection>153.5 4</intersection>
<intersection>161 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>810.5,153.5,838,153.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>810.5 7</intersection>
<intersection>837 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>810.5,149,810.5,153.5</points>
<connection>
<GID>402</GID>
<name>N_in1</name></connection>
<intersection>153.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>830,167.5,834.5,167.5</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<intersection>834.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>834.5,151.5,834.5,167.5</points>
<intersection>151.5 5</intersection>
<intersection>163 6</intersection>
<intersection>167.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>834.5,151.5,838,151.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>834.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>834.5,163,838,163</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>834.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>844,162,847,162</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<connection>
<GID>386</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>803,171.5,819,171.5</points>
<intersection>803 8</intersection>
<intersection>819 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>819,149,819,171.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>168.5 6</intersection>
<intersection>171.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>819,168.5,824,168.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>819 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>803,171.5,803,176.5</points>
<connection>
<GID>481</GID>
<name>OUT_0</name></connection>
<intersection>171.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>793,166.5,824,166.5</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>793 7</intersection>
<intersection>814.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>814.5,147,814.5,166.5</points>
<intersection>147 4</intersection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>814.5,147,819,147</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>814.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>793,166.5,793,176.5</points>
<connection>
<GID>480</GID>
<name>OUT_0</name></connection>
<intersection>166.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>825,148,848,148</points>
<connection>
<GID>396</GID>
<name>OUT</name></connection>
<connection>
<GID>384</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>799,149,808.5,149</points>
<connection>
<GID>435</GID>
<name>OUT</name></connection>
<connection>
<GID>402</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>629.5,149.5,639,149.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<connection>
<GID>444</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>740,149.5,747.5,149.5</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<connection>
<GID>445</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>854,149,862,149</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<connection>
<GID>446</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>514.5,181,516,181</points>
<connection>
<GID>456</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>459</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,184,516,188</points>
<intersection>184 3</intersection>
<intersection>188 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>512.5,184,512.5,188</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>512.5,188,516,188</points>
<intersection>512.5 1</intersection>
<intersection>513.5 8</intersection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>516,184,522.5,184</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>513.5,188,513.5,189.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></vsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520,181,527,181</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<connection>
<GID>457</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>459</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>570,181,571.5,181</points>
<connection>
<GID>470</GID>
<name>OUT_0</name></connection>
<connection>
<GID>468</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,184,571.5,188</points>
<intersection>184 3</intersection>
<intersection>188 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>568,184,568,188</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>568,188,571.5,188</points>
<intersection>568 1</intersection>
<intersection>569.5 5</intersection>
<intersection>571.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>571.5,184,578,184</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>571.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>569.5,188,569.5,189</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></vsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>575.5,181,582,181</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<connection>
<GID>469</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>626.5,181,628,181</points>
<connection>
<GID>471</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>473</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>628,184,628,188</points>
<intersection>184 3</intersection>
<intersection>188 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>624.5,184,624.5,188</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>624.5,188,628,188</points>
<intersection>624.5 1</intersection>
<intersection>626.5 5</intersection>
<intersection>628 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>628,184,634.5,184</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>628 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>626.5,188,626.5,189.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></vsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>632,181,639,181</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<connection>
<GID>472</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>680,180,681.5,180</points>
<connection>
<GID>474</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>476</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>681.5,183,681.5,187</points>
<intersection>183 3</intersection>
<intersection>187 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>678,183,678,187</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>187 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>678,187,681.5,187</points>
<intersection>678 1</intersection>
<intersection>679.5 5</intersection>
<intersection>681.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>681.5,183,688,183</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>681.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>679.5,187,679.5,189</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>187 2</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>685.5,180,692.5,180</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<connection>
<GID>475</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>740,180,741.5,180</points>
<connection>
<GID>477</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>741.5,183,741.5,187</points>
<intersection>183 3</intersection>
<intersection>187 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>738,183,738,187</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>187 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>738,187,741.5,187</points>
<intersection>738 1</intersection>
<intersection>740 5</intersection>
<intersection>741.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>741.5,183,748,183</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>741.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>740,187,740,189.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>187 2</intersection></vsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,180,753,180</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<connection>
<GID>478</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>795,179,796.5,179</points>
<connection>
<GID>482</GID>
<name>OUT_0</name></connection>
<connection>
<GID>480</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>796.5,182,796.5,186</points>
<intersection>182 3</intersection>
<intersection>186 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>793,182,793,186</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>793,186,796.5,186</points>
<intersection>793 1</intersection>
<intersection>794.5 5</intersection>
<intersection>796.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>796.5,182,803,182</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>796.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>794.5,186,794.5,188</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>186 2</intersection></vsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>800.5,179,807.5,179</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<connection>
<GID>481</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>849.5,178.5,851,178.5</points>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection>
<connection>
<GID>483</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>851,181.5,851,185.5</points>
<intersection>181.5 3</intersection>
<intersection>185.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>847.5,181.5,847.5,185.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>185.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>847.5,185.5,851,185.5</points>
<intersection>847.5 1</intersection>
<intersection>849.5 5</intersection>
<intersection>851 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>851,181.5,857.5,181.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>851 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>849.5,185.5,849.5,188</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>185.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>855,178.5,862.5,178.5</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<connection>
<GID>484</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>904.5,178,906,178</points>
<connection>
<GID>486</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>906,181,906,185</points>
<intersection>181 3</intersection>
<intersection>185 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>902.5,181,902.5,185</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>185 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>902.5,185,906,185</points>
<intersection>902.5 1</intersection>
<intersection>904 4</intersection>
<intersection>906 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>906,181,912.5,181</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>906 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>904,185,904,188.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>185 2</intersection></vsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>910,178,918.5,178</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<connection>
<GID>487</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>488</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>182,154,192,154</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 3>
<page 4>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 4>
<page 5>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 5>
<page 6>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 6>
<page 7>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 7>
<page 8>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 8>
<page 9>
<PageViewport>-0.00025201,126.574,938.642,-337.379</PageViewport></page 9></circuit>