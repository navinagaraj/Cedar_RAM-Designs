<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW</type>
<position>68.5,-28</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>BA_TRI_STATE</type>
<position>88.5,-36</position>
<input>
<ID>ENABLE_0</ID>97 </input>
<input>
<ID>IN_0</ID>96 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_AND2</type>
<position>80.5,-36</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>33.5,-28</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>98 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-36</position>
<input>
<ID>ENABLE_0</ID>99 </input>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>45.5,-36</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_DFF_LOW</type>
<position>136.5,-28</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>100 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_TRI_STATE</type>
<position>156.5,-36.5</position>
<input>
<ID>ENABLE_0</ID>101 </input>
<input>
<ID>IN_0</ID>100 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>148.5,-36</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-28</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>102 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>11</ID>
<type>BA_TRI_STATE</type>
<position>121.5,-36</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>113.5,-36</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_DFF_LOW</type>
<position>206,-28</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>104 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_TRI_STATE</type>
<position>226,-36</position>
<input>
<ID>ENABLE_0</ID>105 </input>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>218,-36</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_DFF_LOW</type>
<position>171,-28</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>106 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>17</ID>
<type>BA_TRI_STATE</type>
<position>191,-36</position>
<input>
<ID>ENABLE_0</ID>107 </input>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>183,-36</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_DFF_LOW</type>
<position>274,-28</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>108 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>BA_TRI_STATE</type>
<position>294,-36</position>
<input>
<ID>ENABLE_0</ID>109 </input>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>286,-36</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_DFF_LOW</type>
<position>239,-28</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>110 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>BA_TRI_STATE</type>
<position>259,-36</position>
<input>
<ID>ENABLE_0</ID>111 </input>
<input>
<ID>IN_0</ID>110 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>251,-36</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>14.5,-29</position>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_TRI_STATE</type>
<position>17.5,-37</position>
<input>
<ID>ENABLE_0</ID>114 </input>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>69,-51.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>115 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>BA_TRI_STATE</type>
<position>89,-59.5</position>
<input>
<ID>ENABLE_0</ID>116 </input>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>81,-59.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_DFF_LOW</type>
<position>34,-51.5</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>117 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>31</ID>
<type>BA_TRI_STATE</type>
<position>54,-59.5</position>
<input>
<ID>ENABLE_0</ID>118 </input>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>46,-59.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>137,-51.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>119 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>BA_TRI_STATE</type>
<position>157,-59.5</position>
<input>
<ID>ENABLE_0</ID>120 </input>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>149,-59.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_DFF_LOW</type>
<position>102,-51.5</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>121 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>BA_TRI_STATE</type>
<position>122,-59.5</position>
<input>
<ID>ENABLE_0</ID>122 </input>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>114,-59.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>206.5,-51.5</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>123 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>BA_TRI_STATE</type>
<position>226.5,-59.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>218.5,-59.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_DFF_LOW</type>
<position>171.5,-51.5</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>125 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>43</ID>
<type>BA_TRI_STATE</type>
<position>191.5,-59.5</position>
<input>
<ID>ENABLE_0</ID>126 </input>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>183.5,-59.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>274.5,-51.5</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>127 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>BA_TRI_STATE</type>
<position>294.5,-59.5</position>
<input>
<ID>ENABLE_0</ID>128 </input>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>286.5,-59.5</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW</type>
<position>239.5,-51.5</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>129 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_TRI_STATE</type>
<position>259.5,-59.5</position>
<input>
<ID>ENABLE_0</ID>130 </input>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>251.5,-59.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>15,-52.5</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>BA_TRI_STATE</type>
<position>18,-60.5</position>
<input>
<ID>ENABLE_0</ID>133 </input>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_DFF_LOW</type>
<position>68.5,-74</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>BA_TRI_STATE</type>
<position>88.5,-82</position>
<input>
<ID>ENABLE_0</ID>135 </input>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>80.5,-82</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_DFF_LOW</type>
<position>33.5,-74</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>136 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>57</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-82</position>
<input>
<ID>ENABLE_0</ID>137 </input>
<input>
<ID>IN_0</ID>136 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>45.5,-82</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_DFF_LOW</type>
<position>136.5,-74</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>138 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_TRI_STATE</type>
<position>156.5,-82.5</position>
<input>
<ID>ENABLE_0</ID>139 </input>
<input>
<ID>IN_0</ID>138 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>148.5,-82</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-74</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>140 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>63</ID>
<type>BA_TRI_STATE</type>
<position>121.5,-82</position>
<input>
<ID>ENABLE_0</ID>141 </input>
<input>
<ID>IN_0</ID>140 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>113.5,-82</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_DFF_LOW</type>
<position>206,-74</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>142 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_TRI_STATE</type>
<position>226,-82</position>
<input>
<ID>ENABLE_0</ID>143 </input>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>218,-82</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_DFF_LOW</type>
<position>171,-74</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>144 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>BA_TRI_STATE</type>
<position>191,-82</position>
<input>
<ID>ENABLE_0</ID>145 </input>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>183,-82</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_DFF_LOW</type>
<position>274,-74</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>146 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>72</ID>
<type>BA_TRI_STATE</type>
<position>294,-82</position>
<input>
<ID>ENABLE_0</ID>147 </input>
<input>
<ID>IN_0</ID>146 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>286,-82</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_DFF_LOW</type>
<position>239,-74</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>148 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>BA_TRI_STATE</type>
<position>259,-82</position>
<input>
<ID>ENABLE_0</ID>149 </input>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>251,-82</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>14.5,-75</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>BA_TRI_STATE</type>
<position>17.5,-83</position>
<input>
<ID>ENABLE_0</ID>152 </input>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>79</ID>
<type>HA_JUNC_2</type>
<position>26,-101.5</position>
<input>
<ID>N_in1</ID>153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>80</ID>
<type>HA_JUNC_2</type>
<position>56.5,-96.5</position>
<input>
<ID>N_in1</ID>154 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>81</ID>
<type>HA_JUNC_2</type>
<position>61.5,-101.5</position>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>82</ID>
<type>HA_JUNC_2</type>
<position>91.5,-97</position>
<input>
<ID>N_in1</ID>156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>83</ID>
<type>HA_JUNC_2</type>
<position>95.5,-101.5</position>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>84</ID>
<type>HA_JUNC_2</type>
<position>126.5,-96.5</position>
<input>
<ID>N_in1</ID>158 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>85</ID>
<type>HA_JUNC_2</type>
<position>129.5,-101.5</position>
<input>
<ID>N_in1</ID>159 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>86</ID>
<type>HA_JUNC_2</type>
<position>161.5,-96.5</position>
<input>
<ID>N_in1</ID>160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>87</ID>
<type>HA_JUNC_2</type>
<position>164.5,-101.5</position>
<input>
<ID>N_in1</ID>161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>88</ID>
<type>HA_JUNC_2</type>
<position>195.5,-96</position>
<input>
<ID>N_in1</ID>162 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>89</ID>
<type>HA_JUNC_2</type>
<position>198.5,-101.5</position>
<input>
<ID>N_in1</ID>163 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>90</ID>
<type>HA_JUNC_2</type>
<position>230.5,-96.5</position>
<input>
<ID>N_in1</ID>164 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>91</ID>
<type>HA_JUNC_2</type>
<position>233.5,-101.5</position>
<input>
<ID>N_in1</ID>165 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>92</ID>
<type>HA_JUNC_2</type>
<position>262.5,-96</position>
<input>
<ID>N_in1</ID>166 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>93</ID>
<type>HA_JUNC_2</type>
<position>267.5,-101.5</position>
<input>
<ID>N_in1</ID>167 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>94</ID>
<type>HA_JUNC_2</type>
<position>299.5,-96</position>
<input>
<ID>N_in1</ID>168 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>95</ID>
<type>AE_DFF_LOW</type>
<position>102,44.5</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>96</ID>
<type>BE_DECODER_3x8</type>
<position>-75.5,7</position>
<output>
<ID>OUT_0</ID>152 </output>
<output>
<ID>OUT_1</ID>133 </output>
<output>
<ID>OUT_2</ID>114 </output>
<output>
<ID>OUT_3</ID>95 </output>
<output>
<ID>OUT_4</ID>76 </output>
<output>
<ID>OUT_5</ID>57 </output>
<output>
<ID>OUT_6</ID>38 </output>
<output>
<ID>OUT_7</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>67.5,84</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>1 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_TRI_STATE</type>
<position>87.5,76</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND2</type>
<position>79.5,76</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_DFF_LOW</type>
<position>32.5,84</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>BA_TRI_STATE</type>
<position>52.5,76</position>
<input>
<ID>ENABLE_0</ID>4 </input>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_AND2</type>
<position>44.5,76</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_DFF_LOW</type>
<position>135.5,84</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>104</ID>
<type>BA_TRI_STATE</type>
<position>155.5,76</position>
<input>
<ID>ENABLE_0</ID>6 </input>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>147.5,76</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_DFF_LOW</type>
<position>100.5,84</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_TRI_STATE</type>
<position>120.5,76</position>
<input>
<ID>ENABLE_0</ID>8 </input>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>112.5,76</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AE_DFF_LOW</type>
<position>205,84</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>110</ID>
<type>BA_TRI_STATE</type>
<position>225,76</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>217,76</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_DFF_LOW</type>
<position>170,84</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>11 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>113</ID>
<type>BA_TRI_STATE</type>
<position>190,76</position>
<input>
<ID>ENABLE_0</ID>12 </input>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_AND2</type>
<position>182,76</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_DFF_LOW</type>
<position>273,84</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>116</ID>
<type>BA_TRI_STATE</type>
<position>293,76</position>
<input>
<ID>ENABLE_0</ID>14 </input>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>285,76</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_DFF_LOW</type>
<position>238,84</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>119</ID>
<type>BA_TRI_STATE</type>
<position>258,76</position>
<input>
<ID>ENABLE_0</ID>16 </input>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>250,76</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>13.5,83</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>BA_TRI_STATE</type>
<position>16.5,75</position>
<input>
<ID>ENABLE_0</ID>19 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>123</ID>
<type>HA_JUNC_2</type>
<position>26,92</position>
<input>
<ID>N_in0</ID>153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>124</ID>
<type>HA_JUNC_2</type>
<position>56.5,97</position>
<input>
<ID>N_in0</ID>154 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>125</ID>
<type>HA_JUNC_2</type>
<position>61.5,92</position>
<input>
<ID>N_in0</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>126</ID>
<type>HA_JUNC_2</type>
<position>91.5,97</position>
<input>
<ID>N_in0</ID>156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>127</ID>
<type>HA_JUNC_2</type>
<position>95.5,92</position>
<input>
<ID>N_in0</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>128</ID>
<type>HA_JUNC_2</type>
<position>126.5,97</position>
<input>
<ID>N_in0</ID>158 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>129</ID>
<type>HA_JUNC_2</type>
<position>129.5,92</position>
<input>
<ID>N_in0</ID>159 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>130</ID>
<type>HA_JUNC_2</type>
<position>161.5,97</position>
<input>
<ID>N_in0</ID>160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>131</ID>
<type>HA_JUNC_2</type>
<position>164.5,92</position>
<input>
<ID>N_in0</ID>161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>132</ID>
<type>HA_JUNC_2</type>
<position>195.5,97</position>
<input>
<ID>N_in0</ID>162 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>133</ID>
<type>HA_JUNC_2</type>
<position>198.5,92</position>
<input>
<ID>N_in0</ID>163 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>134</ID>
<type>HA_JUNC_2</type>
<position>230.5,97</position>
<input>
<ID>N_in0</ID>164 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>135</ID>
<type>HA_JUNC_2</type>
<position>233.5,92</position>
<input>
<ID>N_in0</ID>165 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>136</ID>
<type>HA_JUNC_2</type>
<position>262.5,97</position>
<input>
<ID>N_in0</ID>166 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>137</ID>
<type>HA_JUNC_2</type>
<position>267.5,92</position>
<input>
<ID>N_in0</ID>167 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>138</ID>
<type>HA_JUNC_2</type>
<position>299.5,97</position>
<input>
<ID>N_in0</ID>168 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>139</ID>
<type>AE_DFF_LOW</type>
<position>68.5,65</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>140</ID>
<type>BA_TRI_STATE</type>
<position>88.5,57</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_AND2</type>
<position>80.5,57</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_DFF_LOW</type>
<position>33.5,65</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>143</ID>
<type>BA_TRI_STATE</type>
<position>53.5,57</position>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>45.5,57</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_DFF_LOW</type>
<position>136.5,65</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>146</ID>
<type>BA_TRI_STATE</type>
<position>156.5,57</position>
<input>
<ID>ENABLE_0</ID>25 </input>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND2</type>
<position>148.5,57</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_DFF_LOW</type>
<position>101.5,65</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>149</ID>
<type>BA_TRI_STATE</type>
<position>121.5,57</position>
<input>
<ID>ENABLE_0</ID>27 </input>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>113.5,57</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_DFF_LOW</type>
<position>206,65</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>152</ID>
<type>BA_TRI_STATE</type>
<position>226,57</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND2</type>
<position>218,57</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>AE_DFF_LOW</type>
<position>171,65</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>155</ID>
<type>BA_TRI_STATE</type>
<position>191,57</position>
<input>
<ID>ENABLE_0</ID>31 </input>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND2</type>
<position>183,57</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_DFF_LOW</type>
<position>274,65</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>158</ID>
<type>BA_TRI_STATE</type>
<position>294,57</position>
<input>
<ID>ENABLE_0</ID>33 </input>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>286,57</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_DFF_LOW</type>
<position>239,65</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clock</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>BA_TRI_STATE</type>
<position>259,57</position>
<input>
<ID>ENABLE_0</ID>35 </input>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_AND2</type>
<position>251,57</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_AND2</type>
<position>14.5,64</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>BA_TRI_STATE</type>
<position>17.5,56</position>
<input>
<ID>ENABLE_0</ID>38 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_DFF_LOW</type>
<position>69,44.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>BA_TRI_STATE</type>
<position>89,36.5</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_AND2</type>
<position>81,36.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_DFF_LOW</type>
<position>34,44.5</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>169</ID>
<type>BA_TRI_STATE</type>
<position>54,36.5</position>
<input>
<ID>ENABLE_0</ID>42 </input>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>46,36.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AE_DFF_LOW</type>
<position>137,44.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>172</ID>
<type>BA_TRI_STATE</type>
<position>157,36.5</position>
<input>
<ID>ENABLE_0</ID>44 </input>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>149,36.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>BA_TRI_STATE</type>
<position>122,36.5</position>
<input>
<ID>ENABLE_0</ID>46 </input>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>114,36.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_DFF_LOW</type>
<position>206.5,44.5</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>177</ID>
<type>BA_TRI_STATE</type>
<position>226.5,36.5</position>
<input>
<ID>ENABLE_0</ID>48 </input>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>218.5,36.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_DFF_LOW</type>
<position>171.5,44.5</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>180</ID>
<type>BA_TRI_STATE</type>
<position>191.5,36.5</position>
<input>
<ID>ENABLE_0</ID>50 </input>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_AND2</type>
<position>183.5,36.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AE_DFF_LOW</type>
<position>274.5,44.5</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>183</ID>
<type>BA_TRI_STATE</type>
<position>294.5,36.5</position>
<input>
<ID>ENABLE_0</ID>52 </input>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_AND2</type>
<position>286.5,36.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AE_DFF_LOW</type>
<position>239.5,44.5</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>186</ID>
<type>BA_TRI_STATE</type>
<position>259.5,36.5</position>
<input>
<ID>ENABLE_0</ID>54 </input>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND2</type>
<position>251.5,36.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>15,43.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>BA_TRI_STATE</type>
<position>18,35.5</position>
<input>
<ID>ENABLE_0</ID>57 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>190</ID>
<type>AE_DFF_LOW</type>
<position>68.5,21</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>191</ID>
<type>BA_TRI_STATE</type>
<position>88.5,13</position>
<input>
<ID>ENABLE_0</ID>59 </input>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND2</type>
<position>80.5,13</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>AE_DFF_LOW</type>
<position>33.5,21</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>194</ID>
<type>BA_TRI_STATE</type>
<position>53.5,13</position>
<input>
<ID>ENABLE_0</ID>61 </input>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_AND2</type>
<position>45.5,13</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_DFF_LOW</type>
<position>136.5,21</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>62 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_TRI_STATE</type>
<position>156.5,13</position>
<input>
<ID>ENABLE_0</ID>63 </input>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>148.5,13</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_DFF_LOW</type>
<position>101.5,21</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>200</ID>
<type>BA_TRI_STATE</type>
<position>121.5,13</position>
<input>
<ID>ENABLE_0</ID>65 </input>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>113.5,13</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_DFF_LOW</type>
<position>206,21</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>203</ID>
<type>BA_TRI_STATE</type>
<position>226,13</position>
<input>
<ID>ENABLE_0</ID>67 </input>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_AND2</type>
<position>218,13</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AE_DFF_LOW</type>
<position>171,21</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>206</ID>
<type>BA_TRI_STATE</type>
<position>191,13</position>
<input>
<ID>ENABLE_0</ID>69 </input>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_AND2</type>
<position>183,13</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_DFF_LOW</type>
<position>274,21</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>209</ID>
<type>BA_TRI_STATE</type>
<position>294,13</position>
<input>
<ID>ENABLE_0</ID>71 </input>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND2</type>
<position>286,13</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_DFF_LOW</type>
<position>239,21</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>72 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>212</ID>
<type>BA_TRI_STATE</type>
<position>259,13</position>
<input>
<ID>ENABLE_0</ID>73 </input>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>251,13</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>14.5,20</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>BA_TRI_STATE</type>
<position>17.5,12</position>
<input>
<ID>ENABLE_0</ID>76 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_DFF_LOW</type>
<position>68.5,-3.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>77 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>217</ID>
<type>BA_TRI_STATE</type>
<position>88.5,-11.5</position>
<input>
<ID>ENABLE_0</ID>78 </input>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>80.5,-11.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_DFF_LOW</type>
<position>33.5,-3.5</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>79 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>220</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-11.5</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>45.5,-11.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AE_DFF_LOW</type>
<position>136.5,-3.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>223</ID>
<type>BA_TRI_STATE</type>
<position>157,-11.5</position>
<input>
<ID>ENABLE_0</ID>82 </input>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_AND2</type>
<position>148.5,-11.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-3.5</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>83 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>226</ID>
<type>BA_TRI_STATE</type>
<position>121.5,-11.5</position>
<input>
<ID>ENABLE_0</ID>84 </input>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>113.5,-11.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_DFF_LOW</type>
<position>206,-3.5</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>85 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>229</ID>
<type>BA_TRI_STATE</type>
<position>226,-11.5</position>
<input>
<ID>ENABLE_0</ID>86 </input>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>218,-11.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>AE_DFF_LOW</type>
<position>171,-3.5</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>87 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>232</ID>
<type>BA_TRI_STATE</type>
<position>191,-11.5</position>
<input>
<ID>ENABLE_0</ID>88 </input>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>183,-11.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AE_DFF_LOW</type>
<position>274,-3.5</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>89 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>235</ID>
<type>BA_TRI_STATE</type>
<position>294,-11.5</position>
<input>
<ID>ENABLE_0</ID>90 </input>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>286,-11.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AE_DFF_LOW</type>
<position>239,-3.5</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>clock</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>238</ID>
<type>BA_TRI_STATE</type>
<position>259,-11.5</position>
<input>
<ID>ENABLE_0</ID>92 </input>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>251,-11.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>14.5,-4.5</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>BA_TRI_STATE</type>
<position>17.5,-12.5</position>
<input>
<ID>ENABLE_0</ID>95 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,73,72.5,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,77,76.5,77</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,86,72.5,86</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>72.5,73,87.5,73</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,76,85.5,76</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,73,37.5,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,77,41.5,77</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,86,37.5,86</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>37.5,73,52.5,73</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,76,50.5,76</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>101</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,73,140.5,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,77,144.5,77</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,86,140.5,86</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>140.5,73,155.5,73</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>140.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150.5,76,153.5,76</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<connection>
<GID>104</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,73,105.5,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,77,109.5,77</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,86,105.5,86</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>105.5,73,120.5,73</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115.5,76,118.5,76</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>107</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,73,210,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210,77,214,77</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>208,86,210,86</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>210,73,225,73</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,76,223,76</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,73,175,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,77,179,77</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>173,86,175,86</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>175,73,190,73</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,76,188,76</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<connection>
<GID>113</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,73,278,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,77,282,77</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,86,278,86</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>278,73,293,73</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,76,291,76</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,73,243,86</points>
<intersection>73 4</intersection>
<intersection>77 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,77,247,77</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241,86,243,86</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>243,73,258,73</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>253,76,256,76</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<connection>
<GID>119</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,75,282,75</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,83,270,83</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<connection>
<GID>115</GID>
<name>clock</name></connection>
<connection>
<GID>112</GID>
<name>clock</name></connection>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<connection>
<GID>106</GID>
<name>clock</name></connection>
<connection>
<GID>103</GID>
<name>clock</name></connection>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<connection>
<GID>97</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,10.5,-72.5,84</points>
<connection>
<GID>96</GID>
<name>OUT_7</name></connection>
<intersection>77 2</intersection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72.5,84,10.5,84</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-72.5,77,16.5,77</points>
<connection>
<GID>122</GID>
<name>ENABLE_0</name></connection>
<intersection>-72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,54,73.5,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,58,77.5,58</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,67,73.5,67</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,54,88.5,54</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,57,86.5,57</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<connection>
<GID>140</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,54,38.5,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,58,42.5,58</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,67,38.5,67</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38.5,54,53.5,54</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,57,51.5,57</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<connection>
<GID>143</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,54,141.5,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,58,145.5,58</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,67,141.5,67</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,54,156.5,54</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,57,154.5,57</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<connection>
<GID>146</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,54,106.5,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,58,110.5,58</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,67,106.5,67</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106.5,54,121.5,54</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,57,119.5,57</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<connection>
<GID>149</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,54,211,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211,58,215,58</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,67,211,67</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211,54,226,54</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,57,224,57</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<connection>
<GID>152</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,54,176,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,58,180,58</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,67,176,67</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,54,191,54</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186,57,189,57</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<connection>
<GID>155</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,54,279,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,58,283,58</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,67,279,67</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279,54,294,54</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,57,292,57</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<connection>
<GID>158</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,54,244,67</points>
<intersection>54 4</intersection>
<intersection>58 1</intersection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,58,248,58</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,67,244,67</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244,54,259,54</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254,57,257,57</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<connection>
<GID>161</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,56,283,56</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<connection>
<GID>141</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,64,271,64</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<connection>
<GID>157</GID>
<name>clock</name></connection>
<connection>
<GID>154</GID>
<name>clock</name></connection>
<connection>
<GID>151</GID>
<name>clock</name></connection>
<connection>
<GID>148</GID>
<name>clock</name></connection>
<connection>
<GID>145</GID>
<name>clock</name></connection>
<connection>
<GID>142</GID>
<name>clock</name></connection>
<connection>
<GID>139</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71.5,9.5,-71.5,65</points>
<intersection>9.5 4</intersection>
<intersection>58 2</intersection>
<intersection>65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,65,11.5,65</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,58,17.5,58</points>
<connection>
<GID>164</GID>
<name>ENABLE_0</name></connection>
<intersection>-71.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-72.5,9.5,-71.5,9.5</points>
<connection>
<GID>96</GID>
<name>OUT_6</name></connection>
<intersection>-71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,33.5,74,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,37.5,78,37.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,46.5,74,46.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>74,33.5,89,33.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,36.5,87,36.5</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<connection>
<GID>166</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,33.5,39,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,37.5,43,37.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,46.5,39,46.5</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,33.5,54,33.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,36.5,52,36.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,33.5,142,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,37.5,146,37.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,46.5,142,46.5</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142,33.5,157,33.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,36.5,155,36.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>172</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,33.5,107,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,37.5,111,37.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>107,33.5,122,33.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>105,46.5,107,46.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,36.5,120,36.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>174</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,33.5,211.5,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,37.5,215.5,37.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209.5,46.5,211.5,46.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211.5,33.5,226.5,33.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221.5,36.5,224.5,36.5</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<connection>
<GID>177</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,33.5,176.5,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176.5,37.5,180.5,37.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>176.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174.5,46.5,176.5,46.5</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>176.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176.5,33.5,191.5,33.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186.5,36.5,189.5,36.5</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<connection>
<GID>180</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,33.5,279.5,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,37.5,283.5,37.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277.5,46.5,279.5,46.5</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279.5,33.5,294.5,33.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,36.5,292.5,36.5</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<connection>
<GID>183</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,33.5,244.5,46.5</points>
<intersection>33.5 4</intersection>
<intersection>37.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,37.5,248.5,37.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242.5,46.5,244.5,46.5</points>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244.5,33.5,259.5,33.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254.5,36.5,257.5,36.5</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,35.5,283.5,35.5</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<connection>
<GID>167</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,43.5,271.5,43.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<connection>
<GID>185</GID>
<name>clock</name></connection>
<connection>
<GID>182</GID>
<name>clock</name></connection>
<connection>
<GID>179</GID>
<name>clock</name></connection>
<connection>
<GID>176</GID>
<name>clock</name></connection>
<connection>
<GID>171</GID>
<name>clock</name></connection>
<connection>
<GID>168</GID>
<name>clock</name></connection>
<connection>
<GID>165</GID>
<name>clock</name></connection>
<connection>
<GID>95</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,8.5,-70.5,44.5</points>
<intersection>8.5 4</intersection>
<intersection>37.5 2</intersection>
<intersection>44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70.5,44.5,12,44.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-70.5,37.5,18,37.5</points>
<connection>
<GID>189</GID>
<name>ENABLE_0</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-72.5,8.5,-70.5,8.5</points>
<connection>
<GID>96</GID>
<name>OUT_5</name></connection>
<intersection>-70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,10,73.5,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,14,77.5,14</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,23,73.5,23</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,10,88.5,10</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,13,86.5,13</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<connection>
<GID>191</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,10,38.5,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,14,42.5,14</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,23,38.5,23</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38.5,10,53.5,10</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,13,51.5,13</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<connection>
<GID>194</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,10,141.5,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,14,145.5,14</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,23,141.5,23</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,10,156.5,10</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,13,154.5,13</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<connection>
<GID>197</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,10,106.5,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,14,110.5,14</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,23,106.5,23</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106.5,10,121.5,10</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,13,119.5,13</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<connection>
<GID>200</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,10,211,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211,14,215,14</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,23,211,23</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211,10,226,10</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,13,224,13</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<connection>
<GID>203</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,10,176,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,14,180,14</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,23,176,23</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,10,191,10</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186,13,189,13</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<connection>
<GID>206</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,10,279,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,14,283,14</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,23,279,23</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279,10,294,10</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,13,292,13</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<connection>
<GID>209</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,10,244,23</points>
<intersection>10 4</intersection>
<intersection>14 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,14,248,14</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,23,244,23</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244,10,259,10</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254,13,257,13</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<connection>
<GID>212</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,12,283,12</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>192</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,20,271,20</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<connection>
<GID>211</GID>
<name>clock</name></connection>
<connection>
<GID>208</GID>
<name>clock</name></connection>
<connection>
<GID>205</GID>
<name>clock</name></connection>
<connection>
<GID>202</GID>
<name>clock</name></connection>
<connection>
<GID>199</GID>
<name>clock</name></connection>
<connection>
<GID>196</GID>
<name>clock</name></connection>
<connection>
<GID>193</GID>
<name>clock</name></connection>
<connection>
<GID>190</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,7.5,-69.5,21</points>
<intersection>7.5 4</intersection>
<intersection>14 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,21,11.5,21</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,14,17.5,14</points>
<connection>
<GID>215</GID>
<name>ENABLE_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-72.5,7.5,-69.5,7.5</points>
<connection>
<GID>96</GID>
<name>OUT_4</name></connection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-14.5,73.5,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-10.5,77.5,-10.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-1.5,73.5,-1.5</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-14.5,88.5,-14.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-11.5,86.5,-11.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>217</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-14.5,38.5,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-10.5,42.5,-10.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-1.5,38.5,-1.5</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38.5,-14.5,53.5,-14.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-11.5,51.5,-11.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>220</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-15,141.5,-1.5</points>
<intersection>-15 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-10.5,145.5,-10.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-1.5,141.5,-1.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,-15,157,-15</points>
<intersection>141.5 0</intersection>
<intersection>157 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>157,-15,157,-14.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-15 4</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-11.5,155,-11.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<connection>
<GID>223</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-14.5,106.5,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-10.5,110.5,-10.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-1.5,106.5,-1.5</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106.5,-14.5,121.5,-14.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-11.5,119.5,-11.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<connection>
<GID>226</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-14.5,211,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211,-10.5,215,-10.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,-1.5,211,-1.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211,-14.5,226,-14.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-11.5,224,-11.5</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>229</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-14.5,176,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-10.5,180,-10.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-1.5,176,-1.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,-14.5,191,-14.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186,-11.5,189,-11.5</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,-14.5,279,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,-10.5,283,-10.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-1.5,279,-1.5</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279,-14.5,294,-14.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-11.5,292,-11.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<connection>
<GID>235</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-14.5,244,-1.5</points>
<intersection>-14.5 4</intersection>
<intersection>-10.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-10.5,248,-10.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-1.5,244,-1.5</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244,-14.5,259,-14.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254,-11.5,257,-11.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<connection>
<GID>238</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-12.5,283,-12.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<connection>
<GID>218</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-4.5,271,-4.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<connection>
<GID>237</GID>
<name>clock</name></connection>
<connection>
<GID>234</GID>
<name>clock</name></connection>
<connection>
<GID>231</GID>
<name>clock</name></connection>
<connection>
<GID>228</GID>
<name>clock</name></connection>
<connection>
<GID>225</GID>
<name>clock</name></connection>
<connection>
<GID>222</GID>
<name>clock</name></connection>
<connection>
<GID>219</GID>
<name>clock</name></connection>
<connection>
<GID>216</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-10.5,-69.5,6.5</points>
<intersection>-10.5 2</intersection>
<intersection>-3.5 1</intersection>
<intersection>6.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-3.5,11.5,-3.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,-10.5,17.5,-10.5</points>
<connection>
<GID>241</GID>
<name>ENABLE_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-72.5,6.5,-69.5,6.5</points>
<connection>
<GID>96</GID>
<name>OUT_3</name></connection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-39,73.5,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-35,77.5,-35</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-26,73.5,-26</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-39,88.5,-39</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-36,86.5,-36</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-39,38.5,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-35,42.5,-35</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-26,38.5,-26</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38.5,-39,53.5,-39</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-36,51.5,-36</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>5</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-39,141.5,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-35,145.5,-35</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-26,141.5,-26</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,-39,156.5,-39</points>
<intersection>141.5 0</intersection>
<intersection>156.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>156.5,-39.5,156.5,-39</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-39 4</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-36.5,154.5,-36.5</points>
<connection>
<GID>8</GID>
<name>ENABLE_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-36.5,151.5,-36</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-39,106.5,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-35,110.5,-35</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-26,106.5,-26</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106.5,-39,121.5,-39</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-36,119.5,-36</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>11</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-39,211,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211,-35,215,-35</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,-26,211,-26</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211,-39,226,-39</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-36,224,-36</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-39,176,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-35,180,-35</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-26,176,-26</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,-39,191,-39</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186,-36,189,-36</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,-39,279,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,-35,283,-35</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-26,279,-26</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279,-39,294,-39</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-36,292,-36</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-39,244,-26</points>
<intersection>-39 4</intersection>
<intersection>-35 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-35,248,-35</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-26,244,-26</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244,-39,259,-39</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254,-36,257,-36</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>23</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-37,283,-37</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>3</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-29,271,-29</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<connection>
<GID>13</GID>
<name>clock</name></connection>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<connection>
<GID>1</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,-35,-70.5,5.5</points>
<intersection>-35 2</intersection>
<intersection>-28 1</intersection>
<intersection>5.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70.5,-28,11.5,-28</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-70.5,-35,17.5,-35</points>
<connection>
<GID>26</GID>
<name>ENABLE_0</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-72.5,5.5,-70.5,5.5</points>
<connection>
<GID>96</GID>
<name>OUT_2</name></connection>
<intersection>-70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-62.5,74,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-58.5,78,-58.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-49.5,74,-49.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>74,-62.5,89,-62.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-59.5,87,-59.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<connection>
<GID>28</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-62.5,39,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-58.5,43,-58.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-49.5,39,-49.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-62.5,54,-62.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-59.5,52,-59.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<connection>
<GID>31</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-62.5,142,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-58.5,146,-58.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,-49.5,142,-49.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142,-62.5,157,-62.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-59.5,155,-59.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<connection>
<GID>34</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-62.5,107,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-58.5,111,-58.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,-49.5,107,-49.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>107,-62.5,122,-62.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,-59.5,120,-59.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>37</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,-62.5,211.5,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-58.5,215.5,-58.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209.5,-49.5,211.5,-49.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211.5,-62.5,226.5,-62.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221.5,-59.5,224.5,-59.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-62.5,176.5,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176.5,-58.5,180.5,-58.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>176.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174.5,-49.5,176.5,-49.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>176.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176.5,-62.5,191.5,-62.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186.5,-59.5,189.5,-59.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-62.5,279.5,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,-58.5,283.5,-58.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277.5,-49.5,279.5,-49.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279.5,-62.5,294.5,-62.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,-59.5,292.5,-59.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-62.5,244.5,-49.5</points>
<intersection>-62.5 4</intersection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,-58.5,248.5,-58.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242.5,-49.5,244.5,-49.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244.5,-62.5,259.5,-62.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254.5,-59.5,257.5,-59.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<connection>
<GID>49</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-60.5,283.5,-60.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-52.5,271.5,-52.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<connection>
<GID>30</GID>
<name>clock</name></connection>
<connection>
<GID>27</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71.5,-58.5,-71.5,4.5</points>
<intersection>-58.5 2</intersection>
<intersection>-51.5 1</intersection>
<intersection>4.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-51.5,12,-51.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-58.5,18,-58.5</points>
<connection>
<GID>52</GID>
<name>ENABLE_0</name></connection>
<intersection>-71.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-72.5,4.5,-71.5,4.5</points>
<connection>
<GID>96</GID>
<name>OUT_1</name></connection>
<intersection>-71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-85,73.5,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-81,77.5,-81</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-72,73.5,-72</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-85,88.5,-85</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-82,86.5,-82</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-85,38.5,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-81,42.5,-81</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-72,38.5,-72</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38.5,-85,53.5,-85</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-82,51.5,-82</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>57</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-85,141.5,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-81,145.5,-81</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-72,141.5,-72</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,-85,156.5,-85</points>
<intersection>141.5 0</intersection>
<intersection>156.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>156.5,-85.5,156.5,-85</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-85 4</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-82.5,154.5,-82.5</points>
<connection>
<GID>60</GID>
<name>ENABLE_0</name></connection>
<intersection>151.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151.5,-82.5,151.5,-82</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-82.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-85,106.5,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-81,110.5,-81</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-72,106.5,-72</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106.5,-85,121.5,-85</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-82,119.5,-82</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>63</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-85,211,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211,-81,215,-81</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,-72,211,-72</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>211,-85,226,-85</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-82,224,-82</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<connection>
<GID>66</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-85,176,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-81,180,-81</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-72,176,-72</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,-85,191,-85</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186,-82,189,-82</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,-85,279,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,-81,283,-81</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-72,279,-72</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>279,-85,294,-85</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-82,292,-82</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>72</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-85,244,-72</points>
<intersection>-85 4</intersection>
<intersection>-81 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-81,248,-81</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242,-72,244,-72</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>244,-85,259,-85</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>254,-82,257,-82</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-83,283,-83</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<connection>
<GID>55</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-75,271,-75</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<connection>
<GID>65</GID>
<name>clock</name></connection>
<connection>
<GID>62</GID>
<name>clock</name></connection>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<connection>
<GID>53</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,-81,-72.5,3.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>-81 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72.5,-74,11.5,-74</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-72.5,-81,17.5,-81</points>
<connection>
<GID>78</GID>
<name>ENABLE_0</name></connection>
<intersection>-72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-100.5,26,91</points>
<connection>
<GID>79</GID>
<name>N_in1</name></connection>
<connection>
<GID>123</GID>
<name>N_in0</name></connection>
<intersection>-72 10</intersection>
<intersection>-49.5 9</intersection>
<intersection>-26 8</intersection>
<intersection>-1.5 7</intersection>
<intersection>23 6</intersection>
<intersection>46.5 5</intersection>
<intersection>67 4</intersection>
<intersection>86 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26,86,29.5,86</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26,67,30.5,67</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26,46.5,31,46.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>26,23,30.5,23</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>26,-1.5,30.5,-1.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>26,-26,30.5,-26</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>26,-49.5,31,-49.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>26,-72,30.5,-72</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-95.5,56.5,96</points>
<connection>
<GID>80</GID>
<name>N_in1</name></connection>
<connection>
<GID>124</GID>
<name>N_in0</name></connection>
<intersection>-79.5 6</intersection>
<intersection>-57 7</intersection>
<intersection>-33.5 8</intersection>
<intersection>-9 9</intersection>
<intersection>15.5 10</intersection>
<intersection>39 11</intersection>
<intersection>59.5 12</intersection>
<intersection>78.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>53.5,-79.5,56.5,-79.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54,-57,56.5,-57</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>53.5,-33.5,56.5,-33.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>53.5,-9,56.5,-9</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>53.5,15.5,56.5,15.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>54,39,56.5,39</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>53.5,59.5,56.5,59.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>52.5,78.5,56.5,78.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-100.5,61.5,91</points>
<connection>
<GID>81</GID>
<name>N_in1</name></connection>
<connection>
<GID>125</GID>
<name>N_in0</name></connection>
<intersection>-72 10</intersection>
<intersection>-49.5 9</intersection>
<intersection>-26 8</intersection>
<intersection>-1.5 7</intersection>
<intersection>23 6</intersection>
<intersection>46.5 5</intersection>
<intersection>67 4</intersection>
<intersection>86 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,86,64.5,86</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,67,65.5,67</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>61.5,46.5,66,46.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61.5,23,65.5,23</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>61.5,-1.5,65.5,-1.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>61.5,-26,65.5,-26</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>61.5,-49.5,66,-49.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61.5,-72,65.5,-72</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-96,91.5,96</points>
<connection>
<GID>82</GID>
<name>N_in1</name></connection>
<connection>
<GID>126</GID>
<name>N_in0</name></connection>
<intersection>-79.5 6</intersection>
<intersection>-57 7</intersection>
<intersection>-33.5 8</intersection>
<intersection>-9 9</intersection>
<intersection>15.5 10</intersection>
<intersection>39 11</intersection>
<intersection>59.5 12</intersection>
<intersection>78.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>88.5,-79.5,91.5,-79.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89,-57,91.5,-57</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>88.5,-33.5,91.5,-33.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>88.5,-9,91.5,-9</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>88.5,15.5,91.5,15.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>89,39,91.5,39</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>88.5,59.5,91.5,59.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>87.5,78.5,91.5,78.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-100.5,95.5,91</points>
<connection>
<GID>83</GID>
<name>N_in1</name></connection>
<connection>
<GID>127</GID>
<name>N_in0</name></connection>
<intersection>-72 3</intersection>
<intersection>-49.5 4</intersection>
<intersection>-26 5</intersection>
<intersection>-1.5 6</intersection>
<intersection>23 7</intersection>
<intersection>46.5 11</intersection>
<intersection>67 9</intersection>
<intersection>86 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95.5,-72,98.5,-72</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>95.5,-49.5,99,-49.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>95.5,-26,98.5,-26</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>95.5,-1.5,98.5,-1.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>95.5,23,98.5,23</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>95.5,67,98.5,67</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>95.5,86,97.5,86</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>95.5,46.5,99,46.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-95.5,126.5,96</points>
<connection>
<GID>84</GID>
<name>N_in1</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<intersection>-79.5 13</intersection>
<intersection>-57 12</intersection>
<intersection>-33.5 11</intersection>
<intersection>-9 10</intersection>
<intersection>15.5 9</intersection>
<intersection>39 8</intersection>
<intersection>59.5 7</intersection>
<intersection>78.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>120.5,78.5,126.5,78.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>121.5,59.5,126.5,59.5</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>122,39,126.5,39</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>121.5,15.5,126.5,15.5</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>121.5,-9,126.5,-9</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>121.5,-33.5,126.5,-33.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>122,-57,126.5,-57</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>121.5,-79.5,126.5,-79.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-100.5,129.5,91</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>-72 10</intersection>
<intersection>-49.5 9</intersection>
<intersection>-26 8</intersection>
<intersection>-1.5 7</intersection>
<intersection>23 6</intersection>
<intersection>46.5 5</intersection>
<intersection>67 4</intersection>
<intersection>86 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>129.5,86,132.5,86</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>129.5,67,133.5,67</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>129.5,46.5,134,46.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>129.5,23,133.5,23</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>129.5,-1.5,133.5,-1.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>129.5,-26,133.5,-26</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>129.5,-49.5,134,-49.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>129.5,-72,133.5,-72</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-95.5,161.5,96</points>
<connection>
<GID>86</GID>
<name>N_in1</name></connection>
<connection>
<GID>130</GID>
<name>N_in0</name></connection>
<intersection>-80 6</intersection>
<intersection>-57.5 7</intersection>
<intersection>-34 8</intersection>
<intersection>-9.5 9</intersection>
<intersection>15 10</intersection>
<intersection>39 11</intersection>
<intersection>60 12</intersection>
<intersection>78.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>156.5,-80,161.5,-80</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>157,-57.5,161.5,-57.5</points>
<intersection>157 19</intersection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>156.5,-34,161.5,-34</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,-9.5,161.5,-9.5</points>
<intersection>157 17</intersection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156.5,15,161.5,15</points>
<intersection>156.5 16</intersection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>157,39,161.5,39</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>156.5,60,161.5,60</points>
<intersection>156.5 15</intersection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>155.5,78.5,161.5,78.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>161.5 0</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>156.5,59.5,156.5,60</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>60 12</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>156.5,15,156.5,15.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>15 10</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>157,-9.5,157,-9</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 9</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>157,-57.5,157,-57</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-100.5,164.5,91</points>
<connection>
<GID>87</GID>
<name>N_in1</name></connection>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>-72 3</intersection>
<intersection>-49.5 4</intersection>
<intersection>-26 5</intersection>
<intersection>-1.5 6</intersection>
<intersection>23 7</intersection>
<intersection>46.5 8</intersection>
<intersection>67 9</intersection>
<intersection>86 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>164.5,-72,168,-72</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-49.5,168.5,-49.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>164.5,-26,168,-26</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>164.5,-1.5,168,-1.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>164.5,23,168,23</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>164.5,46.5,168.5,46.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>164.5,67,168,67</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>164.5,86,167,86</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-95,195.5,96</points>
<connection>
<GID>88</GID>
<name>N_in1</name></connection>
<connection>
<GID>132</GID>
<name>N_in0</name></connection>
<intersection>-79.5 13</intersection>
<intersection>-57 12</intersection>
<intersection>-33.5 11</intersection>
<intersection>-9 10</intersection>
<intersection>15.5 9</intersection>
<intersection>39 8</intersection>
<intersection>59.5 7</intersection>
<intersection>78.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>190,78.5,195.5,78.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>191,59.5,195.5,59.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>191.5,39,195.5,39</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>191,15.5,195.5,15.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>191,-9,195.5,-9</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>191,-33.5,195.5,-33.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>191.5,-57,195.5,-57</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>191,-79.5,195.5,-79.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-100.5,198.5,91</points>
<connection>
<GID>89</GID>
<name>N_in1</name></connection>
<connection>
<GID>133</GID>
<name>N_in0</name></connection>
<intersection>-72 10</intersection>
<intersection>-49.5 9</intersection>
<intersection>-26 8</intersection>
<intersection>-1.5 7</intersection>
<intersection>23 6</intersection>
<intersection>46.5 5</intersection>
<intersection>67 4</intersection>
<intersection>86 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198.5,86,202,86</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,67,203,67</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>198.5,46.5,203.5,46.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>198.5,23,203,23</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>198.5,-1.5,203,-1.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>198.5,-26,203,-26</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>198.5,-49.5,203.5,-49.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>198.5,-72,203,-72</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-95.5,230.5,96</points>
<connection>
<GID>90</GID>
<name>N_in1</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>-79.5 6</intersection>
<intersection>-57 7</intersection>
<intersection>-33.5 8</intersection>
<intersection>-9 9</intersection>
<intersection>15.5 10</intersection>
<intersection>39 11</intersection>
<intersection>59.5 12</intersection>
<intersection>78.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>226,-79.5,230.5,-79.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>226.5,-57,230.5,-57</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>226,-33.5,230.5,-33.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>226,-9,230.5,-9</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>226,15.5,230.5,15.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>226.5,39,230.5,39</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>226,59.5,230.5,59.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>225,78.5,230.5,78.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233.5,-100.5,233.5,91</points>
<connection>
<GID>91</GID>
<name>N_in1</name></connection>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<intersection>-72 3</intersection>
<intersection>-49.5 4</intersection>
<intersection>-26 5</intersection>
<intersection>-1.5 6</intersection>
<intersection>23 7</intersection>
<intersection>46.5 8</intersection>
<intersection>67 9</intersection>
<intersection>86 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>233.5,-72,236,-72</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>233.5,-49.5,236.5,-49.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>233.5,-26,236,-26</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>233.5,-1.5,236,-1.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>233.5,23,236,23</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>233.5,46.5,236.5,46.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>233.5,67,236,67</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>233.5,86,235,86</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>233.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-95,262.5,96</points>
<connection>
<GID>92</GID>
<name>N_in1</name></connection>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<intersection>-79.5 15</intersection>
<intersection>-57 14</intersection>
<intersection>-33.5 13</intersection>
<intersection>-9 12</intersection>
<intersection>15.5 11</intersection>
<intersection>39 10</intersection>
<intersection>59.5 9</intersection>
<intersection>78.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>258,78.5,262.5,78.5</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>259,59.5,262.5,59.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>259.5,39,262.5,39</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>259,15.5,262.5,15.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>259,-9,262.5,-9</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>259,-33.5,262.5,-33.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>259.5,-57,262.5,-57</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>259,-79.5,262.5,-79.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>262.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-100.5,267.5,91</points>
<connection>
<GID>93</GID>
<name>N_in1</name></connection>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<intersection>-72 10</intersection>
<intersection>-49.5 9</intersection>
<intersection>-26 8</intersection>
<intersection>-1.5 7</intersection>
<intersection>23 6</intersection>
<intersection>46.5 5</intersection>
<intersection>67 4</intersection>
<intersection>86 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>267.5,86,270,86</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>267.5,67,271,67</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>267.5,46.5,271.5,46.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>267.5,23,271,23</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>267.5,-1.5,271,-1.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>267.5,-26,271,-26</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>267.5,-49.5,271.5,-49.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>267.5,-72,271,-72</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299.5,-95,299.5,96</points>
<connection>
<GID>94</GID>
<name>N_in1</name></connection>
<connection>
<GID>138</GID>
<name>N_in0</name></connection>
<intersection>-79.5 6</intersection>
<intersection>-57 7</intersection>
<intersection>-33.5 8</intersection>
<intersection>-9 9</intersection>
<intersection>15.5 10</intersection>
<intersection>39 11</intersection>
<intersection>59.5 12</intersection>
<intersection>78.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>294,-79.5,299.5,-79.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>294.5,-57,299.5,-57</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>294,-33.5,299.5,-33.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>294,-9,299.5,-9</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>294,15.5,299.5,15.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>294.5,39,299.5,39</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>294,59.5,299.5,59.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>293,78.5,299.5,78.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>299.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>