<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 0>
<page 1>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 1>
<page 2>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 2>
<page 3>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 3>
<page 4>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 4>
<page 5>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 5>
<page 6>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 6>
<page 7>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 7>
<page 8>
<PageViewport>-72.0143,159.513,420.91,-84.1305</PageViewport>
<gate>
<ID>1</ID>
<type>AA_AND2</type>
<position>68,-24.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>BA_TRI_STATE</type>
<position>75,-24.5</position>
<input>
<ID>ENABLE_0</ID>1 </input>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_DFF_LOW</type>
<position>56,-17</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>2 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>HA_JUNC_2</type>
<position>52,-35.5</position>
<input>
<ID>N_in1</ID>205 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>6</ID>
<type>HA_JUNC_2</type>
<position>83,-36</position>
<input>
<ID>N_in1</ID>83 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>9</ID>
<type>HA_JUNC_2</type>
<position>115,-36</position>
<input>
<ID>N_in1</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>11</ID>
<type>HA_JUNC_2</type>
<position>146,-35</position>
<input>
<ID>N_in1</ID>85 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>13</ID>
<type>HA_JUNC_2</type>
<position>176,-34</position>
<input>
<ID>N_in1</ID>86 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>15</ID>
<type>HA_JUNC_2</type>
<position>207,-33.5</position>
<input>
<ID>N_in1</ID>87 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>17</ID>
<type>HA_JUNC_2</type>
<position>269,-34.5</position>
<input>
<ID>N_in1</ID>89 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>18</ID>
<type>HA_JUNC_2</type>
<position>238,-32.5</position>
<input>
<ID>N_in1</ID>88 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>19</ID>
<type>HA_JUNC_2</type>
<position>52,106</position>
<input>
<ID>N_in0</ID>205 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>20</ID>
<type>HA_JUNC_2</type>
<position>83,106</position>
<input>
<ID>N_in0</ID>83 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>21</ID>
<type>HA_JUNC_2</type>
<position>115,106</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>99.5,-24.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>BA_TRI_STATE</type>
<position>106.5,-24.5</position>
<input>
<ID>ENABLE_0</ID>15 </input>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>87,-17</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>130,-24.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_TRI_STATE</type>
<position>137,-24.5</position>
<input>
<ID>ENABLE_0</ID>17 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>118,-17</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>18 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>161.5,-24.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>BA_TRI_STATE</type>
<position>168.5,-24.5</position>
<input>
<ID>ENABLE_0</ID>19 </input>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_DFF_LOW</type>
<position>149,-17</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>191,-24.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>BA_TRI_STATE</type>
<position>198,-24.5</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>179,-17</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_AND2</type>
<position>222.5,-24.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>BA_TRI_STATE</type>
<position>229.5,-24.5</position>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_DFF_LOW</type>
<position>210,-17</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>253,-24.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BA_TRI_STATE</type>
<position>260,-24.5</position>
<input>
<ID>ENABLE_0</ID>25 </input>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>241,-17</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>284.5,-24.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>BA_TRI_STATE</type>
<position>291.5,-24.5</position>
<input>
<ID>ENABLE_0</ID>27 </input>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_DFF_LOW</type>
<position>272,-17</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clock</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>68.5,-7.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>BA_TRI_STATE</type>
<position>75.5,-7.5</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>56.5,0</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>100,-7.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>BA_TRI_STATE</type>
<position>107,-7.5</position>
<input>
<ID>ENABLE_0</ID>31 </input>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW</type>
<position>87.5,0</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>130.5,-7.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>BA_TRI_STATE</type>
<position>137.5,-7.5</position>
<input>
<ID>ENABLE_0</ID>33 </input>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_DFF_LOW</type>
<position>118.5,0</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>162,-7.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>BA_TRI_STATE</type>
<position>169,-7.5</position>
<input>
<ID>ENABLE_0</ID>35 </input>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_DFF_LOW</type>
<position>149.5,0</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>36 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>191.5,-7.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>BA_TRI_STATE</type>
<position>198.5,-7.5</position>
<input>
<ID>ENABLE_0</ID>37 </input>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_DFF_LOW</type>
<position>179.5,0</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>223,-7.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_TRI_STATE</type>
<position>230,-7.5</position>
<input>
<ID>ENABLE_0</ID>39 </input>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_DFF_LOW</type>
<position>210.5,0</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>253.5,-7.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_TRI_STATE</type>
<position>260.5,-7.5</position>
<input>
<ID>ENABLE_0</ID>41 </input>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_DFF_LOW</type>
<position>241.5,0</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>42 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>285,-7.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_TRI_STATE</type>
<position>292,-7.5</position>
<input>
<ID>ENABLE_0</ID>43 </input>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_DFF_LOW</type>
<position>272.5,0</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>69,8.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>BA_TRI_STATE</type>
<position>76,8.5</position>
<input>
<ID>ENABLE_0</ID>45 </input>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_DFF_LOW</type>
<position>57,16</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>100.5,8.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>BA_TRI_STATE</type>
<position>107.5,8.5</position>
<input>
<ID>ENABLE_0</ID>47 </input>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_DFF_LOW</type>
<position>88,16</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>131,8.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_TRI_STATE</type>
<position>138,8.5</position>
<input>
<ID>ENABLE_0</ID>49 </input>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_DFF_LOW</type>
<position>119,16</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>162.5,8.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>BA_TRI_STATE</type>
<position>169.5,8.5</position>
<input>
<ID>ENABLE_0</ID>51 </input>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>150,16</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>192,8.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>BA_TRI_STATE</type>
<position>199,8.5</position>
<input>
<ID>ENABLE_0</ID>53 </input>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_DFF_LOW</type>
<position>180,16</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>223.5,8.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>BA_TRI_STATE</type>
<position>230.5,8.5</position>
<input>
<ID>ENABLE_0</ID>55 </input>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_DFF_LOW</type>
<position>211,16</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>56 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND2</type>
<position>254,8.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>BA_TRI_STATE</type>
<position>261,8.5</position>
<input>
<ID>ENABLE_0</ID>57 </input>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_DFF_LOW</type>
<position>242,16</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND2</type>
<position>285.5,8.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>BA_TRI_STATE</type>
<position>292.5,8.5</position>
<input>
<ID>ENABLE_0</ID>59 </input>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_DFF_LOW</type>
<position>273,16</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>69.5,24</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>BA_TRI_STATE</type>
<position>76.5,24</position>
<input>
<ID>ENABLE_0</ID>61 </input>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_DFF_LOW</type>
<position>57.5,31.5</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>62 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND2</type>
<position>101,24</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>BA_TRI_STATE</type>
<position>108,24</position>
<input>
<ID>ENABLE_0</ID>63 </input>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_DFF_LOW</type>
<position>88.5,31.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>131.5,24</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_TRI_STATE</type>
<position>138.5,24</position>
<input>
<ID>ENABLE_0</ID>65 </input>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_DFF_LOW</type>
<position>119.5,31.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND2</type>
<position>163,24</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>BA_TRI_STATE</type>
<position>170,24</position>
<input>
<ID>ENABLE_0</ID>67 </input>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_DFF_LOW</type>
<position>150.5,31.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>192.5,24</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>BA_TRI_STATE</type>
<position>199.5,24</position>
<input>
<ID>ENABLE_0</ID>69 </input>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_DFF_LOW</type>
<position>180.5,31.5</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND2</type>
<position>224,24</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_TRI_STATE</type>
<position>231,24</position>
<input>
<ID>ENABLE_0</ID>71 </input>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_DFF_LOW</type>
<position>211.5,31.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>72 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>254.5,24</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>BA_TRI_STATE</type>
<position>261.5,24</position>
<input>
<ID>ENABLE_0</ID>73 </input>
<input>
<ID>IN_0</ID>74 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_DFF_LOW</type>
<position>242.5,31.5</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>286,24</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>BA_TRI_STATE</type>
<position>293,24</position>
<input>
<ID>ENABLE_0</ID>75 </input>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_DFF_LOW</type>
<position>273.5,31.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>115</ID>
<type>HA_JUNC_2</type>
<position>146,106</position>
<input>
<ID>N_in0</ID>85 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>116</ID>
<type>HA_JUNC_2</type>
<position>177,105.5</position>
<input>
<ID>N_in0</ID>86 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>117</ID>
<type>HA_JUNC_2</type>
<position>207,106</position>
<input>
<ID>N_in0</ID>87 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>118</ID>
<type>HA_JUNC_2</type>
<position>238,106</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>119</ID>
<type>HA_JUNC_2</type>
<position>269,105.5</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>120</ID>
<type>HA_JUNC_2</type>
<position>81,113</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>121</ID>
<type>HA_JUNC_2</type>
<position>81,-44</position>
<input>
<ID>N_in1</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>122</ID>
<type>HA_JUNC_2</type>
<position>112,-44.5</position>
<input>
<ID>N_in1</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>123</ID>
<type>HA_JUNC_2</type>
<position>144,-43</position>
<input>
<ID>N_in1</ID>92 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>124</ID>
<type>HA_JUNC_2</type>
<position>174.5,-42.5</position>
<input>
<ID>N_in1</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>125</ID>
<type>HA_JUNC_2</type>
<position>205,-42.5</position>
<input>
<ID>N_in1</ID>94 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>126</ID>
<type>HA_JUNC_2</type>
<position>236,-42.5</position>
<input>
<ID>N_in1</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>127</ID>
<type>HA_JUNC_2</type>
<position>267,-43</position>
<input>
<ID>N_in1</ID>96 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>128</ID>
<type>HA_JUNC_2</type>
<position>297.5,-42.5</position>
<input>
<ID>N_in1</ID>97 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>129</ID>
<type>HA_JUNC_2</type>
<position>297.5,114.5</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>130</ID>
<type>HA_JUNC_2</type>
<position>267,114</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>131</ID>
<type>HA_JUNC_2</type>
<position>236,113</position>
<input>
<ID>N_in0</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>132</ID>
<type>HA_JUNC_2</type>
<position>205,113</position>
<input>
<ID>N_in0</ID>94 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>133</ID>
<type>HA_JUNC_2</type>
<position>174.5,113</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>134</ID>
<type>HA_JUNC_2</type>
<position>144,113</position>
<input>
<ID>N_in0</ID>92 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>135</ID>
<type>HA_JUNC_2</type>
<position>112,113</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>136</ID>
<type>BE_DECODER_3x8</type>
<position>2,40.5</position>
<output>
<ID>OUT_0</ID>105 </output>
<output>
<ID>OUT_1</ID>104 </output>
<output>
<ID>OUT_2</ID>103 </output>
<output>
<ID>OUT_3</ID>102 </output>
<output>
<ID>OUT_4</ID>101 </output>
<output>
<ID>OUT_5</ID>100 </output>
<output>
<ID>OUT_6</ID>99 </output>
<output>
<ID>OUT_7</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>212</ID>
<type>BA_TRI_STATE</type>
<position>44,26</position>
<input>
<ID>ENABLE_0</ID>102 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>38,30.5</position>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>BA_TRI_STATE</type>
<position>44,10</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND2</type>
<position>38,15</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>BA_TRI_STATE</type>
<position>44,-6</position>
<input>
<ID>ENABLE_0</ID>104 </input>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>38,-1</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>BA_TRI_STATE</type>
<position>44,-23</position>
<input>
<ID>ENABLE_0</ID>105 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>38,-18</position>
<input>
<ID>IN_0</ID>105 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>69,40.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>BA_TRI_STATE</type>
<position>76,40.5</position>
<input>
<ID>ENABLE_0</ID>141 </input>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_DFF_LOW</type>
<position>57,48</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>142 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>224</ID>
<type>BA_TRI_STATE</type>
<position>45,91</position>
<input>
<ID>ENABLE_0</ID>98 </input>
<output>
<ID>OUT_0</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_AND2</type>
<position>38.5,95.5</position>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>BA_TRI_STATE</type>
<position>45,75</position>
<input>
<ID>ENABLE_0</ID>99 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>100.5,40.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_AND2</type>
<position>38,80</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>BA_TRI_STATE</type>
<position>107.5,40.5</position>
<input>
<ID>ENABLE_0</ID>143 </input>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>230</ID>
<type>BA_TRI_STATE</type>
<position>45,59</position>
<input>
<ID>ENABLE_0</ID>100 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AE_DFF_LOW</type>
<position>88,48</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>144 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_AND2</type>
<position>38,64</position>
<input>
<ID>IN_0</ID>100 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>131,40.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>BA_TRI_STATE</type>
<position>45,42</position>
<input>
<ID>ENABLE_0</ID>101 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>235</ID>
<type>BA_TRI_STATE</type>
<position>138,40.5</position>
<input>
<ID>ENABLE_0</ID>145 </input>
<input>
<ID>IN_0</ID>146 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>38,47</position>
<input>
<ID>IN_0</ID>101 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AE_DFF_LOW</type>
<position>119,48</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>146 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_AND2</type>
<position>162.5,40.5</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>BA_TRI_STATE</type>
<position>169.5,40.5</position>
<input>
<ID>ENABLE_0</ID>147 </input>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_DFF_LOW</type>
<position>150,48</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>148 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_AND2</type>
<position>192,40.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>BA_TRI_STATE</type>
<position>199,40.5</position>
<input>
<ID>ENABLE_0</ID>149 </input>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>243</ID>
<type>AE_DFF_LOW</type>
<position>180,48</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>150 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_AND2</type>
<position>223.5,40.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>BA_TRI_STATE</type>
<position>230.5,40.5</position>
<input>
<ID>ENABLE_0</ID>151 </input>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>246</ID>
<type>AE_DFF_LOW</type>
<position>211,48</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>152 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_AND2</type>
<position>254,40.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>BA_TRI_STATE</type>
<position>261,40.5</position>
<input>
<ID>ENABLE_0</ID>153 </input>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>249</ID>
<type>AE_DFF_LOW</type>
<position>242,48</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>154 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>285.5,40.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>BA_TRI_STATE</type>
<position>292.5,40.5</position>
<input>
<ID>ENABLE_0</ID>155 </input>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AE_DFF_LOW</type>
<position>273,48</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>156 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>69.5,57.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>BA_TRI_STATE</type>
<position>76.5,57.5</position>
<input>
<ID>ENABLE_0</ID>157 </input>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_DFF_LOW</type>
<position>57.5,65</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>158 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>101,57.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>BA_TRI_STATE</type>
<position>108,57.5</position>
<input>
<ID>ENABLE_0</ID>159 </input>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>258</ID>
<type>AE_DFF_LOW</type>
<position>88.5,65</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>160 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_AND2</type>
<position>131.5,57.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>BA_TRI_STATE</type>
<position>138.5,57.5</position>
<input>
<ID>ENABLE_0</ID>161 </input>
<input>
<ID>IN_0</ID>162 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>261</ID>
<type>AE_DFF_LOW</type>
<position>119.5,65</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>162 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>163,57.5</position>
<input>
<ID>IN_0</ID>164 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>BA_TRI_STATE</type>
<position>170,57.5</position>
<input>
<ID>ENABLE_0</ID>163 </input>
<input>
<ID>IN_0</ID>164 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_DFF_LOW</type>
<position>150.5,65</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>164 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>192.5,57.5</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>BA_TRI_STATE</type>
<position>199.5,57.5</position>
<input>
<ID>ENABLE_0</ID>165 </input>
<input>
<ID>IN_0</ID>166 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>267</ID>
<type>AE_DFF_LOW</type>
<position>180.5,65</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>166 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>224,57.5</position>
<input>
<ID>IN_0</ID>168 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>BA_TRI_STATE</type>
<position>231,57.5</position>
<input>
<ID>ENABLE_0</ID>167 </input>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_DFF_LOW</type>
<position>211.5,65</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>168 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND2</type>
<position>254.5,57.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>BA_TRI_STATE</type>
<position>261.5,57.5</position>
<input>
<ID>ENABLE_0</ID>169 </input>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>273</ID>
<type>AE_DFF_LOW</type>
<position>242.5,65</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>170 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_AND2</type>
<position>286,57.5</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>BA_TRI_STATE</type>
<position>293,57.5</position>
<input>
<ID>ENABLE_0</ID>171 </input>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>276</ID>
<type>AE_DFF_LOW</type>
<position>273.5,65</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>172 </output>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_AND2</type>
<position>70,73.5</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>BA_TRI_STATE</type>
<position>77,73.5</position>
<input>
<ID>ENABLE_0</ID>173 </input>
<input>
<ID>IN_0</ID>174 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>279</ID>
<type>AE_DFF_LOW</type>
<position>58,81</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>174 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_AND2</type>
<position>101.5,73.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>BA_TRI_STATE</type>
<position>108.5,73.5</position>
<input>
<ID>ENABLE_0</ID>175 </input>
<input>
<ID>IN_0</ID>176 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>282</ID>
<type>AE_DFF_LOW</type>
<position>89,81</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>176 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_AND2</type>
<position>132,73.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>284</ID>
<type>BA_TRI_STATE</type>
<position>139,73.5</position>
<input>
<ID>ENABLE_0</ID>177 </input>
<input>
<ID>IN_0</ID>178 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>285</ID>
<type>AE_DFF_LOW</type>
<position>120,81</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>178 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_AND2</type>
<position>163.5,73.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>BA_TRI_STATE</type>
<position>170.5,73.5</position>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_DFF_LOW</type>
<position>151,81</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>180 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>289</ID>
<type>AA_AND2</type>
<position>193,73.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>290</ID>
<type>BA_TRI_STATE</type>
<position>200,73.5</position>
<input>
<ID>ENABLE_0</ID>181 </input>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_DFF_LOW</type>
<position>181,81</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>182 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_AND2</type>
<position>224.5,73.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>293</ID>
<type>BA_TRI_STATE</type>
<position>231.5,73.5</position>
<input>
<ID>ENABLE_0</ID>183 </input>
<input>
<ID>IN_0</ID>184 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_DFF_LOW</type>
<position>212,81</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>184 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_AND2</type>
<position>255,73.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>296</ID>
<type>BA_TRI_STATE</type>
<position>262,73.5</position>
<input>
<ID>ENABLE_0</ID>185 </input>
<input>
<ID>IN_0</ID>186 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>297</ID>
<type>AE_DFF_LOW</type>
<position>243,81</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>186 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND2</type>
<position>286.5,73.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>BA_TRI_STATE</type>
<position>293.5,73.5</position>
<input>
<ID>ENABLE_0</ID>187 </input>
<input>
<ID>IN_0</ID>188 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_DFF_LOW</type>
<position>274,81</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>188 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_AND2</type>
<position>70.5,89</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>BA_TRI_STATE</type>
<position>77.5,89</position>
<input>
<ID>ENABLE_0</ID>189 </input>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_DFF_LOW</type>
<position>58.5,96.5</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>190 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>102,89</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>BA_TRI_STATE</type>
<position>109,89</position>
<input>
<ID>ENABLE_0</ID>191 </input>
<input>
<ID>IN_0</ID>192 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>89.5,96.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>192 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_AND2</type>
<position>132.5,89</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>BA_TRI_STATE</type>
<position>139.5,89</position>
<input>
<ID>ENABLE_0</ID>193 </input>
<input>
<ID>IN_0</ID>194 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_DFF_LOW</type>
<position>120.5,96.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>194 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_AND2</type>
<position>164,89</position>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>BA_TRI_STATE</type>
<position>171,89</position>
<input>
<ID>ENABLE_0</ID>195 </input>
<input>
<ID>IN_0</ID>196 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>312</ID>
<type>AE_DFF_LOW</type>
<position>151.5,96.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>196 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>193.5,89</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>BA_TRI_STATE</type>
<position>200.5,89</position>
<input>
<ID>ENABLE_0</ID>197 </input>
<input>
<ID>IN_0</ID>198 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>315</ID>
<type>AE_DFF_LOW</type>
<position>181.5,96.5</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>198 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>225,89</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>BA_TRI_STATE</type>
<position>232,89</position>
<input>
<ID>ENABLE_0</ID>199 </input>
<input>
<ID>IN_0</ID>200 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_DFF_LOW</type>
<position>212.5,96.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>200 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>255.5,89</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>BA_TRI_STATE</type>
<position>262.5,89</position>
<input>
<ID>ENABLE_0</ID>201 </input>
<input>
<ID>IN_0</ID>202 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>321</ID>
<type>AE_DFF_LOW</type>
<position>243.5,96.5</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>202 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>322</ID>
<type>AA_AND2</type>
<position>287,89</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>BA_TRI_STATE</type>
<position>294,89</position>
<input>
<ID>ENABLE_0</ID>203 </input>
<input>
<ID>IN_0</ID>204 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_DFF_LOW</type>
<position>274.5,96.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>204 </output>
<input>
<ID>clock</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>135.5,89,137.5,89</points>
<connection>
<GID>308</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>307</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,85.5,139.5,86</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,85.5,139.5,85.5</points>
<intersection>125.5 2</intersection>
<intersection>139.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>125.5,85.5,125.5,98.5</points>
<intersection>85.5 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>125.5,90,129.5,90</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>125.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>123.5,98.5,125.5,98.5</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>125.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>71,-24.5,73,-24.5</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>167,89,169,89</points>
<connection>
<GID>311</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>310</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-28,75,-27.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-28,75,-28</points>
<intersection>61 2</intersection>
<intersection>75 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>61,-28,61,-15</points>
<intersection>-28 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>61,-23.5,65,-23.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>61 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59,-15,61,-15</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>61 2</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,72.5,283.5,72.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<connection>
<GID>289</GID>
<name>IN_1</name></connection>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,72.5,47.5,75</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,86,171,86</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>157 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>157,86,157,98.5</points>
<intersection>86 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>157,90,161,90</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>157 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>154.5,98.5,157,98.5</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>157 2</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,80,271,80</points>
<connection>
<GID>300</GID>
<name>clock</name></connection>
<connection>
<GID>297</GID>
<name>clock</name></connection>
<connection>
<GID>294</GID>
<name>clock</name></connection>
<connection>
<GID>291</GID>
<name>clock</name></connection>
<connection>
<GID>288</GID>
<name>clock</name></connection>
<connection>
<GID>285</GID>
<name>clock</name></connection>
<connection>
<GID>282</GID>
<name>clock</name></connection>
<connection>
<GID>279</GID>
<name>clock</name></connection>
<connection>
<GID>228</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>196.5,89,198.5,89</points>
<connection>
<GID>314</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>313</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,85.5,200.5,86</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,85.5,200.5,85.5</points>
<intersection>186.5 2</intersection>
<intersection>200.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>186.5,85.5,186.5,98.5</points>
<intersection>85.5 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>186.5,90,190.5,90</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>186.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>184.5,98.5,186.5,98.5</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>186.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,56.5,283,56.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,56.5,47.5,59</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>228,89,230,89</points>
<connection>
<GID>317</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>316</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,64,270.5,64</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<connection>
<GID>255</GID>
<name>clock</name></connection>
<connection>
<GID>258</GID>
<name>clock</name></connection>
<connection>
<GID>261</GID>
<name>clock</name></connection>
<connection>
<GID>264</GID>
<name>clock</name></connection>
<connection>
<GID>267</GID>
<name>clock</name></connection>
<connection>
<GID>273</GID>
<name>clock</name></connection>
<connection>
<GID>276</GID>
<name>clock</name></connection>
<connection>
<GID>270</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218,86,232,86</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,86,218,98.5</points>
<intersection>86 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>218,90,222,90</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>218 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>215.5,98.5,218,98.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,47,270,47</points>
<connection>
<GID>252</GID>
<name>clock</name></connection>
<connection>
<GID>249</GID>
<name>clock</name></connection>
<connection>
<GID>246</GID>
<name>clock</name></connection>
<connection>
<GID>243</GID>
<name>clock</name></connection>
<connection>
<GID>240</GID>
<name>clock</name></connection>
<connection>
<GID>237</GID>
<name>clock</name></connection>
<connection>
<GID>231</GID>
<name>clock</name></connection>
<connection>
<GID>223</GID>
<name>clock</name></connection>
<connection>
<GID>236</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>258.5,89,260.5,89</points>
<connection>
<GID>320</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>319</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,39.5,282.5,39.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,39.5,47.5,42</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,85.5,262.5,86</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248.5,85.5,262.5,85.5</points>
<intersection>248.5 2</intersection>
<intersection>262.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>248.5,85.5,248.5,98.5</points>
<intersection>85.5 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>248.5,90,252.5,90</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>248.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>246.5,98.5,248.5,98.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>248.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>290,89,292,89</points>
<connection>
<GID>323</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>322</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,30.5,270.5,30.5</points>
<connection>
<GID>114</GID>
<name>clock</name></connection>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<connection>
<GID>108</GID>
<name>clock</name></connection>
<connection>
<GID>105</GID>
<name>clock</name></connection>
<connection>
<GID>102</GID>
<name>clock</name></connection>
<connection>
<GID>99</GID>
<name>clock</name></connection>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<connection>
<GID>93</GID>
<name>clock</name></connection>
<connection>
<GID>214</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>280,86,294,86</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>280 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>280,86,280,98.5</points>
<intersection>86 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>280,90,284,90</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>280 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>277.5,98.5,280,98.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>280 2</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,23,283,23</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>46.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46.5,23,46.5,26</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>23 1</intersection></vsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-34.5,52,105</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>N_in1</name></connection>
<intersection>-15 14</intersection>
<intersection>2 12</intersection>
<intersection>18 10</intersection>
<intersection>33.5 8</intersection>
<intersection>50 6</intersection>
<intersection>67 4</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,98.5,55.5,98.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,83,55,83</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52,67,54.5,67</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>52,50,54,50</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>52,33.5,54.5,33.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>52,18,54,18</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>52,2,53.5,2</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>52,-15,53,-15</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,15,270,15</points>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<connection>
<GID>87</GID>
<name>clock</name></connection>
<connection>
<GID>84</GID>
<name>clock</name></connection>
<connection>
<GID>81</GID>
<name>clock</name></connection>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<connection>
<GID>75</GID>
<name>clock</name></connection>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<connection>
<GID>216</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,88,284,88</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,88,47.5,91</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>88 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,7.5,282.5,7.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>46.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46.5,7.5,46.5,10</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<intersection>7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,95.5,271.5,95.5</points>
<connection>
<GID>303</GID>
<name>clock</name></connection>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<connection>
<GID>315</GID>
<name>clock</name></connection>
<connection>
<GID>318</GID>
<name>clock</name></connection>
<connection>
<GID>321</GID>
<name>clock</name></connection>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<connection>
<GID>225</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>102.5,-24.5,104.5,-24.5</points>
<connection>
<GID>23</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92.5,-27.5,106.5,-27.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>92.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>92.5,-27.5,92.5,-15</points>
<intersection>-27.5 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>92.5,-23.5,96.5,-23.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>92.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>90,-15,92.5,-15</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>92.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>133,-24.5,135,-24.5</points>
<connection>
<GID>26</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>25</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-28,137,-27.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-28,137,-28</points>
<intersection>123 2</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-28,123,-15</points>
<intersection>-28 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>123,-23.5,127,-23.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>121,-15,123,-15</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>164.5,-24.5,166.5,-24.5</points>
<connection>
<GID>29</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154.5,-27.5,168.5,-27.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>154.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>154.5,-27.5,154.5,-15</points>
<intersection>-27.5 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>154.5,-23.5,158.5,-23.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>154.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>152,-15,154.5,-15</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>154.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>194,-24.5,196,-24.5</points>
<connection>
<GID>32</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-28,198,-27.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-28,198,-28</points>
<intersection>184 2</intersection>
<intersection>198 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>184,-28,184,-15</points>
<intersection>-28 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>184,-23.5,188,-23.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>184 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>182,-15,184,-15</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>184 2</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>225.5,-24.5,227.5,-24.5</points>
<connection>
<GID>35</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215.5,-27.5,229.5,-27.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>215.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>215.5,-27.5,215.5,-15</points>
<intersection>-27.5 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>215.5,-23.5,219.5,-23.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>215.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>213,-15,215.5,-15</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>215.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>256,-24.5,258,-24.5</points>
<connection>
<GID>38</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>37</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-28,260,-27.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246,-28,260,-28</points>
<intersection>246 2</intersection>
<intersection>260 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>246,-28,246,-15</points>
<intersection>-28 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>246,-23.5,250,-23.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>246 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>244,-15,246,-15</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>246 2</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>287.5,-24.5,289.5,-24.5</points>
<connection>
<GID>41</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-27.5,291.5,-27.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>277.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>277.5,-27.5,277.5,-15</points>
<intersection>-27.5 1</intersection>
<intersection>-23.5 4</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>277.5,-23.5,281.5,-23.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>277.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>275,-15,277.5,-15</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>277.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>71.5,-7.5,73.5,-7.5</points>
<connection>
<GID>44</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>43</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-11,75.5,-10.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-11,75.5,-11</points>
<intersection>61.5 2</intersection>
<intersection>75.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>61.5,-11,61.5,2</points>
<intersection>-11 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-6.5,65.5,-6.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>61.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59.5,2,61.5,2</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>61.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>103,-7.5,105,-7.5</points>
<connection>
<GID>47</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93,-10.5,107,-10.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>93 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>93,-10.5,93,2</points>
<intersection>-10.5 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>93,-6.5,97,-6.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>93 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>90.5,2,93,2</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>93 2</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>133.5,-7.5,135.5,-7.5</points>
<connection>
<GID>50</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-11,137.5,-10.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-11,137.5,-11</points>
<intersection>123.5 2</intersection>
<intersection>137.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123.5,-11,123.5,2</points>
<intersection>-11 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>123.5,-6.5,127.5,-6.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>123.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>121.5,2,123.5,2</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>123.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>165,-7.5,167,-7.5</points>
<connection>
<GID>53</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>52</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155,-10.5,169,-10.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>155 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>155,-10.5,155,2</points>
<intersection>-10.5 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>155,-6.5,159,-6.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>155 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>152.5,2,155,2</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>155 2</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>194.5,-7.5,196.5,-7.5</points>
<connection>
<GID>56</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>55</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-11,198.5,-10.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-11,198.5,-11</points>
<intersection>184.5 2</intersection>
<intersection>198.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>184.5,-11,184.5,2</points>
<intersection>-11 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>184.5,-6.5,188.5,-6.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>184.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>182.5,2,184.5,2</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>184.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>226,-7.5,228,-7.5</points>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>58</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-10.5,230,-10.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>216 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>216,-10.5,216,2</points>
<intersection>-10.5 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>216,-6.5,220,-6.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>216 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>213.5,2,216,2</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>216 2</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>256.5,-7.5,258.5,-7.5</points>
<connection>
<GID>62</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>61</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-11,260.5,-10.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246.5,-11,260.5,-11</points>
<intersection>246.5 2</intersection>
<intersection>260.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>246.5,-11,246.5,2</points>
<intersection>-11 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>246.5,-6.5,250.5,-6.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>246.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>244.5,2,246.5,2</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>246.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>288,-7.5,290,-7.5</points>
<connection>
<GID>65</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>64</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>278,-10.5,292,-10.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>278 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>278,-10.5,278,2</points>
<intersection>-10.5 1</intersection>
<intersection>-6.5 4</intersection>
<intersection>2 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>278,-6.5,282,-6.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>278 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>275.5,2,278,2</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>278 2</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>72,8.5,74,8.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<connection>
<GID>68</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,5,76,5.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,5,76,5</points>
<intersection>62 2</intersection>
<intersection>76 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,5,62,18</points>
<intersection>5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,9.5,66,9.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60,18,62,18</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>103.5,8.5,105.5,8.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>71</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,5.5,107.5,5.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>93.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>93.5,5.5,93.5,18</points>
<intersection>5.5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>93.5,9.5,97.5,9.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>93.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>91,18,93.5,18</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>93.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>134,8.5,136,8.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,5,138,5.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,5,138,5</points>
<intersection>124 2</intersection>
<intersection>138 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,5,124,18</points>
<intersection>5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124,9.5,128,9.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>122,18,124,18</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>165.5,8.5,167.5,8.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>77</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155.5,5.5,169.5,5.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>155.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>155.5,5.5,155.5,18</points>
<intersection>5.5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>155.5,9.5,159.5,9.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>155.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>153,18,155.5,18</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>155.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>195,8.5,197,8.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,5,199,5.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,5,199,5</points>
<intersection>185 2</intersection>
<intersection>199 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>185,5,185,18</points>
<intersection>5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>185,9.5,189,9.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>185 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>183,18,185,18</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>185 2</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>226.5,8.5,228.5,8.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<connection>
<GID>83</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216.5,5.5,230.5,5.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>216.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>216.5,5.5,216.5,18</points>
<intersection>5.5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>216.5,9.5,220.5,9.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>216.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>214,18,216.5,18</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>216.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>257,8.5,259,8.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,5,261,5.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,5,261,5</points>
<intersection>247 2</intersection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>247,5,247,18</points>
<intersection>5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>247,9.5,251,9.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>247 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>245,18,247,18</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>247 2</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>288.5,8.5,290.5,8.5</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>278.5,5.5,292.5,5.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>278.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>278.5,5.5,278.5,18</points>
<intersection>5.5 1</intersection>
<intersection>9.5 4</intersection>
<intersection>18 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>278.5,9.5,282.5,9.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>278.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>276,18,278.5,18</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>278.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>72.5,24,74.5,24</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,20.5,76.5,21</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,20.5,76.5,20.5</points>
<intersection>62.5 2</intersection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,20.5,62.5,33.5</points>
<intersection>20.5 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62.5,25,66.5,25</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60.5,33.5,62.5,33.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>104,24,106,24</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<connection>
<GID>95</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,21,108,21</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>94 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>94,21,94,33.5</points>
<intersection>21 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94,25,98,25</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>94 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>91.5,33.5,94,33.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>94 2</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>134.5,24,136.5,24</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,20.5,138.5,21</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,20.5,138.5,20.5</points>
<intersection>124.5 2</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124.5,20.5,124.5,33.5</points>
<intersection>20.5 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124.5,25,128.5,25</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>124.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>122.5,33.5,124.5,33.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>124.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166,24,168,24</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<connection>
<GID>101</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,21,170,21</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,21,156,33.5</points>
<intersection>21 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>156,25,160,25</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>153.5,33.5,156,33.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>195.5,24,197.5,24</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>104</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,20.5,199.5,21</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,20.5,199.5,20.5</points>
<intersection>185.5 2</intersection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>185.5,20.5,185.5,33.5</points>
<intersection>20.5 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>185.5,25,189.5,25</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>185.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>183.5,33.5,185.5,33.5</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>185.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>227,24,229,24</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<connection>
<GID>107</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,21,231,21</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,21,217,33.5</points>
<intersection>21 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>217,25,221,25</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>214.5,33.5,217,33.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>257.5,24,259.5,24</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,20.5,261.5,21</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247.5,20.5,261.5,20.5</points>
<intersection>247.5 2</intersection>
<intersection>261.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>247.5,20.5,247.5,33.5</points>
<intersection>20.5 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>247.5,25,251.5,25</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>247.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>245.5,33.5,247.5,33.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>247.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>289,24,291,24</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<connection>
<GID>113</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>279,21,293,21</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>279 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>279,21,279,33.5</points>
<intersection>21 1</intersection>
<intersection>25 4</intersection>
<intersection>33.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>279,25,283,25</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>279 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>276.5,33.5,279,33.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>279 2</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-1,269.5,-1</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<connection>
<GID>60</GID>
<name>clock</name></connection>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<connection>
<GID>54</GID>
<name>clock</name></connection>
<connection>
<GID>57</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-8.5,282,-8.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>46.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46.5,-8.5,46.5,-6</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-18,269,-18</points>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<connection>
<GID>30</GID>
<name>clock</name></connection>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<connection>
<GID>220</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-25.5,47.5,-23</points>
<intersection>-25.5 2</intersection>
<intersection>-23 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-25.5,281.5,-25.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46.5,-23,47.5,-23</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-35,83,105</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<connection>
<GID>6</GID>
<name>N_in1</name></connection>
<intersection>-15 1</intersection>
<intersection>2 3</intersection>
<intersection>18 4</intersection>
<intersection>33.5 5</intersection>
<intersection>50 6</intersection>
<intersection>67 7</intersection>
<intersection>83 8</intersection>
<intersection>98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-15,84,-15</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,98.5,86.5,98.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83,2,84.5,2</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>83,18,85,18</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>83,33.5,85.5,33.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>83,50,85,50</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>83,67,85.5,67</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>83,83,86,83</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-35,115,105</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>N_in1</name></connection>
<intersection>2 9</intersection>
<intersection>18 10</intersection>
<intersection>33.5 7</intersection>
<intersection>50 11</intersection>
<intersection>67 5</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,98.5,117.5,98.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,83,117,83</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>115,67,116.5,67</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>115,33.5,116.5,33.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>115,2,115.5,2</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>115,18,116,18</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>115,50,116,50</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-34,146,105</points>
<connection>
<GID>11</GID>
<name>N_in1</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>2 38</intersection>
<intersection>18 21</intersection>
<intersection>33.5 7</intersection>
<intersection>50 20</intersection>
<intersection>67 5</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146,98.5,148.5,98.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146,83,148,83</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>146,67,147.5,67</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>146,33.5,147.5,33.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>146,50,147,50</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>146,18,147,18</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>146,2,146.5,2</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,2,177,104.5</points>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>2 9</intersection>
<intersection>33.5 7</intersection>
<intersection>67 5</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,98.5,178.5,98.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,83,178,83</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>177,67,177.5,67</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>177,33.5,177.5,33.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>176,2,177,2</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>176 10</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>176,-33,176,2</points>
<connection>
<GID>13</GID>
<name>N_in1</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>2 9</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-32.5,207,105</points>
<connection>
<GID>117</GID>
<name>N_in0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>N_in1</name></connection>
<intersection>2 13</intersection>
<intersection>18 11</intersection>
<intersection>33.5 9</intersection>
<intersection>50 7</intersection>
<intersection>67 5</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,98.5,209.5,98.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,83,209,83</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>207,67,208.5,67</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>207,50,208,50</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>207,33.5,208.5,33.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>207,18,208,18</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>207,2,207.5,2</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-31.5,238,105</points>
<connection>
<GID>118</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>N_in1</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>2 13</intersection>
<intersection>18 11</intersection>
<intersection>33.5 9</intersection>
<intersection>50 7</intersection>
<intersection>67 5</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,98.5,240.5,98.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238,83,240,83</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>238,67,239.5,67</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>238,50,239,50</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>238,33.5,239.5,33.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>238,18,239,18</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>238,2,238.5,2</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-33.5,269,104.5</points>
<connection>
<GID>119</GID>
<name>N_in0</name></connection>
<connection>
<GID>17</GID>
<name>N_in1</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>2 13</intersection>
<intersection>18 10</intersection>
<intersection>33.5 8</intersection>
<intersection>50 6</intersection>
<intersection>67 4</intersection>
<intersection>83 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269,98.5,271.5,98.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269,83,271,83</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>269,67,270.5,67</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>269,50,270,50</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>269,33.5,270.5,33.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>269,18,270,18</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>269,2,269.5,2</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-43,81,112</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<connection>
<GID>121</GID>
<name>N_in1</name></connection>
<intersection>-22 13</intersection>
<intersection>-5 12</intersection>
<intersection>11 11</intersection>
<intersection>26.5 10</intersection>
<intersection>43 9</intersection>
<intersection>60 8</intersection>
<intersection>76 7</intersection>
<intersection>91.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77.5,91.5,81,91.5</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>77,76,81,76</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>76.5,60,81,60</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>76,43,81,43</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>76.5,26.5,81,26.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>76,11,81,11</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>75.5,-5,81,-5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>75,-22,81,-22</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-43.5,112,112</points>
<connection>
<GID>122</GID>
<name>N_in1</name></connection>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<intersection>-22 13</intersection>
<intersection>-5 12</intersection>
<intersection>11 11</intersection>
<intersection>26.5 10</intersection>
<intersection>43 9</intersection>
<intersection>60 8</intersection>
<intersection>76 7</intersection>
<intersection>91.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>109,91.5,112,91.5</points>
<connection>
<GID>305</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>108.5,76,112,76</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>108,60,112,60</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>107.5,43,112,43</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>108,26.5,112,26.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>107.5,11,112,11</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>107,-5,112,-5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>106.5,-22,112,-22</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-42,144,112</points>
<connection>
<GID>123</GID>
<name>N_in1</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>-22 13</intersection>
<intersection>-5 12</intersection>
<intersection>11 11</intersection>
<intersection>26.5 10</intersection>
<intersection>43 9</intersection>
<intersection>60 8</intersection>
<intersection>76 7</intersection>
<intersection>91.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139.5,91.5,144,91.5</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,76,144,76</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>138.5,60,144,60</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>138,43,144,43</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>138.5,26.5,144,26.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>138,11,144,11</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>137.5,-5,144,-5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>137,-22,144,-22</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-41.5,174.5,112</points>
<connection>
<GID>124</GID>
<name>N_in1</name></connection>
<connection>
<GID>133</GID>
<name>N_in0</name></connection>
<intersection>-22 18</intersection>
<intersection>-5 17</intersection>
<intersection>11 16</intersection>
<intersection>26.5 15</intersection>
<intersection>43 14</intersection>
<intersection>60 13</intersection>
<intersection>76 12</intersection>
<intersection>91.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>171,91.5,174.5,91.5</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>170.5,76,174.5,76</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>170,60,174.5,60</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>169.5,43,174.5,43</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>170,26.5,174.5,26.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>169.5,11,174.5,11</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>169,-5,174.5,-5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>168.5,-22,174.5,-22</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-41.5,205,112</points>
<connection>
<GID>125</GID>
<name>N_in1</name></connection>
<connection>
<GID>132</GID>
<name>N_in0</name></connection>
<intersection>-22 9</intersection>
<intersection>-5 10</intersection>
<intersection>11 11</intersection>
<intersection>26.5 12</intersection>
<intersection>43 13</intersection>
<intersection>60 14</intersection>
<intersection>76 15</intersection>
<intersection>91.5 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>198,-22,205,-22</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>198.5,-5,205,-5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>199,11,205,11</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>199.5,26.5,205,26.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>199,43,205,43</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>199.5,60,205,60</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>200,76,205,76</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>200.5,91.5,205,91.5</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-41.5,236,112</points>
<connection>
<GID>126</GID>
<name>N_in1</name></connection>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>-22 6</intersection>
<intersection>-5 7</intersection>
<intersection>11 8</intersection>
<intersection>26.5 9</intersection>
<intersection>43 10</intersection>
<intersection>60 11</intersection>
<intersection>76 12</intersection>
<intersection>91.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>229.5,-22,236,-22</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>230,-5,236,-5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>230.5,11,236,11</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>231,26.5,236,26.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>230.5,43,236,43</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>231,60,236,60</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>231.5,76,236,76</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>232,91.5,236,91.5</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<intersection>236 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267,-42,267,113</points>
<connection>
<GID>127</GID>
<name>N_in1</name></connection>
<connection>
<GID>130</GID>
<name>N_in0</name></connection>
<intersection>-22 6</intersection>
<intersection>-5 7</intersection>
<intersection>11 8</intersection>
<intersection>26.5 9</intersection>
<intersection>43 10</intersection>
<intersection>60 11</intersection>
<intersection>76 12</intersection>
<intersection>91.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>260,-22,267,-22</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>260.5,-5,267,-5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>261,11,267,11</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>261.5,26.5,267,26.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>261,43,267,43</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>261.5,60,267,60</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>262,76,267,76</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>262.5,91.5,267,91.5</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>267 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-41.5,297.5,113.5</points>
<connection>
<GID>128</GID>
<name>N_in1</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>-22 3</intersection>
<intersection>-5 4</intersection>
<intersection>11 5</intersection>
<intersection>26.5 6</intersection>
<intersection>43 7</intersection>
<intersection>60 8</intersection>
<intersection>76 9</intersection>
<intersection>91.5 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-22,297.5,-22</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>292,-5,297.5,-5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>292.5,11,297.5,11</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>293,26.5,297.5,26.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>292.5,43,297.5,43</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>293,60,297.5,60</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>293.5,76,297.5,76</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>294,91.5,297.5,91.5</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,44,6,93</points>
<intersection>44 2</intersection>
<intersection>93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,93,45,93</points>
<connection>
<GID>224</GID>
<name>ENABLE_0</name></connection>
<intersection>6 0</intersection>
<intersection>31 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,44,6,44</points>
<connection>
<GID>136</GID>
<name>OUT_7</name></connection>
<intersection>6 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31,93,31,96.5</points>
<intersection>93 1</intersection>
<intersection>96.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,96.5,35.5,96.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,43,8,77.5</points>
<intersection>43 2</intersection>
<intersection>77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,77.5,45,77.5</points>
<intersection>8 0</intersection>
<intersection>31 4</intersection>
<intersection>45 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,43,8,43</points>
<connection>
<GID>136</GID>
<name>OUT_6</name></connection>
<intersection>8 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45,77,45,77.5</points>
<connection>
<GID>226</GID>
<name>ENABLE_0</name></connection>
<intersection>77.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>31,77.5,31,81</points>
<intersection>77.5 1</intersection>
<intersection>81 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,81,35,81</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,42,10,65</points>
<intersection>42 2</intersection>
<intersection>65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,65,35,65</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection>
<intersection>31 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,42,10,42</points>
<connection>
<GID>136</GID>
<name>OUT_5</name></connection>
<intersection>10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,61,31,65</points>
<intersection>61 4</intersection>
<intersection>65 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31,61,45,61</points>
<connection>
<GID>230</GID>
<name>ENABLE_0</name></connection>
<intersection>31 3</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,41,12,48</points>
<intersection>41 2</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,48,35,48</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection>
<intersection>31 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,41,12,41</points>
<connection>
<GID>136</GID>
<name>OUT_4</name></connection>
<intersection>12 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,44,31,48</points>
<intersection>44 4</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31,44,45,44</points>
<connection>
<GID>234</GID>
<name>ENABLE_0</name></connection>
<intersection>31 3</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,28,12,40</points>
<intersection>28 1</intersection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,28,44,28</points>
<connection>
<GID>212</GID>
<name>ENABLE_0</name></connection>
<intersection>12 0</intersection>
<intersection>31 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,40,12,40</points>
<connection>
<GID>136</GID>
<name>OUT_3</name></connection>
<intersection>12 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31,28,31,31.5</points>
<intersection>28 1</intersection>
<intersection>31.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,31.5,35,31.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,12,10,39</points>
<intersection>12 1</intersection>
<intersection>39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,12,44,12</points>
<connection>
<GID>215</GID>
<name>ENABLE_0</name></connection>
<intersection>10 0</intersection>
<intersection>31 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,39,10,39</points>
<connection>
<GID>136</GID>
<name>OUT_2</name></connection>
<intersection>10 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31,12,31,16</points>
<intersection>12 1</intersection>
<intersection>16 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,16,35,16</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-3.5,8,38</points>
<intersection>-3.5 1</intersection>
<intersection>38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-3.5,44,-3.5</points>
<intersection>8 0</intersection>
<intersection>31 4</intersection>
<intersection>44 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,38,8,38</points>
<connection>
<GID>136</GID>
<name>OUT_1</name></connection>
<intersection>8 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-4,44,-3.5</points>
<connection>
<GID>217</GID>
<name>ENABLE_0</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>31,-3.5,31,0</points>
<intersection>-3.5 1</intersection>
<intersection>0 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,0,35,0</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-21,6,37</points>
<intersection>-21 1</intersection>
<intersection>37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-21,44,-21</points>
<connection>
<GID>219</GID>
<name>ENABLE_0</name></connection>
<intersection>6 0</intersection>
<intersection>31 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,37,6,37</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31,-21,31,-17</points>
<intersection>-21 1</intersection>
<intersection>-17 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,-17,35,-17</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>72,40.5,74,40.5</points>
<connection>
<GID>222</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,37,76,37.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,37,76,37</points>
<intersection>62 2</intersection>
<intersection>76 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,37,62,50</points>
<intersection>37 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,41.5,66,41.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60,50,62,50</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>103.5,40.5,105.5,40.5</points>
<connection>
<GID>229</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>227</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,37.5,107.5,37.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>93.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>93.5,37.5,93.5,50</points>
<intersection>37.5 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>93.5,41.5,97.5,41.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>93.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>91,50,93.5,50</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>93.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>134,40.5,136,40.5</points>
<connection>
<GID>235</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>233</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,37,138,37.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,37,138,37</points>
<intersection>124 2</intersection>
<intersection>138 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,37,124,50</points>
<intersection>37 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124,41.5,128,41.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>124 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>122,50,124,50</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>165.5,40.5,167.5,40.5</points>
<connection>
<GID>239</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>238</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155.5,37.5,169.5,37.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>155.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>155.5,37.5,155.5,50</points>
<intersection>37.5 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>155.5,41.5,159.5,41.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>155.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>153,50,155.5,50</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>155.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>195,40.5,197,40.5</points>
<connection>
<GID>242</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>241</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,37,199,37.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,37,199,37</points>
<intersection>185 2</intersection>
<intersection>199 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>185,37,185,50</points>
<intersection>37 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>185,41.5,189,41.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>185 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>183,50,185,50</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>185 2</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>226.5,40.5,228.5,40.5</points>
<connection>
<GID>245</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>244</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216.5,37.5,230.5,37.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>216.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>216.5,37.5,216.5,50</points>
<intersection>37.5 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>216.5,41.5,220.5,41.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>216.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>214,50,216.5,50</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>216.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>257,40.5,259,40.5</points>
<connection>
<GID>248</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>247</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,37,261,37.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,37,261,37</points>
<intersection>247 2</intersection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>247,37,247,50</points>
<intersection>37 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>247,41.5,251,41.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>247 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>245,50,247,50</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>247 2</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>288.5,40.5,290.5,40.5</points>
<connection>
<GID>251</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>250</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>278.5,37.5,292.5,37.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>278.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>278.5,37.5,278.5,50</points>
<intersection>37.5 1</intersection>
<intersection>41.5 4</intersection>
<intersection>50 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>278.5,41.5,282.5,41.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>278.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>276,50,278.5,50</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>278.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>72.5,57.5,74.5,57.5</points>
<connection>
<GID>254</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>253</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,54,76.5,54.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,54,76.5,54</points>
<intersection>62.5 2</intersection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62.5,54,62.5,67</points>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62.5,58.5,66.5,58.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60.5,67,62.5,67</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>104,57.5,106,57.5</points>
<connection>
<GID>257</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>256</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,54.5,108,54.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>94 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>94,54.5,94,67</points>
<intersection>54.5 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94,58.5,98,58.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>94 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>91.5,67,94,67</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>94 2</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>134.5,57.5,136.5,57.5</points>
<connection>
<GID>260</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>259</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,54,138.5,54.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,54,138.5,54</points>
<intersection>124.5 2</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124.5,54,124.5,67</points>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124.5,58.5,128.5,58.5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>124.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>122.5,67,124.5,67</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>124.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166,57.5,168,57.5</points>
<connection>
<GID>263</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>262</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,54.5,170,54.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,54.5,156,67</points>
<intersection>54.5 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>156,58.5,160,58.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>156 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>153.5,67,156,67</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>195.5,57.5,197.5,57.5</points>
<connection>
<GID>266</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>265</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,54,199.5,54.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,54,199.5,54</points>
<intersection>185.5 2</intersection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>185.5,54,185.5,67</points>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>185.5,58.5,189.5,58.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>185.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>183.5,67,185.5,67</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>185.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>227,57.5,229,57.5</points>
<connection>
<GID>269</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>268</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,54.5,231,54.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,54.5,217,67</points>
<intersection>54.5 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>217,58.5,221,58.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>217 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>214.5,67,217,67</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>257.5,57.5,259.5,57.5</points>
<connection>
<GID>272</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>271</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,54,261.5,54.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247.5,54,261.5,54</points>
<intersection>247.5 2</intersection>
<intersection>261.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>247.5,54,247.5,67</points>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>247.5,58.5,251.5,58.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>247.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>245.5,67,247.5,67</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>247.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>289,57.5,291,57.5</points>
<connection>
<GID>275</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>274</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>279,54.5,293,54.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>279 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>279,54.5,279,67</points>
<intersection>54.5 1</intersection>
<intersection>58.5 4</intersection>
<intersection>67 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>279,58.5,283,58.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>279 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>276.5,67,279,67</points>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection>
<intersection>279 2</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>73,73.5,75,73.5</points>
<connection>
<GID>278</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>277</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,70,77,70.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,70,77,70</points>
<intersection>63 2</intersection>
<intersection>77 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>63,70,63,83</points>
<intersection>70 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63,74.5,67,74.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>63 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61,83,63,83</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>63 2</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>104.5,73.5,106.5,73.5</points>
<connection>
<GID>281</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>280</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,70.5,108.5,70.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>94.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>94.5,70.5,94.5,83</points>
<intersection>70.5 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94.5,74.5,98.5,74.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>94.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>92,83,94.5,83</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>94.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>135,73.5,137,73.5</points>
<connection>
<GID>284</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>283</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,70,139,70.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,70,139,70</points>
<intersection>125 2</intersection>
<intersection>139 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>125,70,125,83</points>
<intersection>70 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>125,74.5,129,74.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>125 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>123,83,125,83</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>125 2</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>166.5,73.5,168.5,73.5</points>
<connection>
<GID>287</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>286</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,70.5,170.5,70.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,70.5,156.5,83</points>
<intersection>70.5 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>156.5,74.5,160.5,74.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>156.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>154,83,156.5,83</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>156.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>196,73.5,198,73.5</points>
<connection>
<GID>290</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>289</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200,70,200,70.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186,70,200,70</points>
<intersection>186 2</intersection>
<intersection>200 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>186,70,186,83</points>
<intersection>70 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>186,74.5,190,74.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>186 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>184,83,186,83</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<intersection>186 2</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>227.5,73.5,229.5,73.5</points>
<connection>
<GID>293</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>292</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217.5,70.5,231.5,70.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>217.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217.5,70.5,217.5,83</points>
<intersection>70.5 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>217.5,74.5,221.5,74.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>217.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>215,83,217.5,83</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>217.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>258,73.5,260,73.5</points>
<connection>
<GID>296</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>295</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,70,262,70.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,70,262,70</points>
<intersection>248 2</intersection>
<intersection>262 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>248,70,248,83</points>
<intersection>70 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>248,74.5,252,74.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>248 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>246,83,248,83</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>248 2</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>289.5,73.5,291.5,73.5</points>
<connection>
<GID>299</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>298</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>279.5,70.5,293.5,70.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>279.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>279.5,70.5,279.5,83</points>
<intersection>70.5 1</intersection>
<intersection>74.5 4</intersection>
<intersection>83 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>279.5,74.5,283.5,74.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>279.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>277,83,279.5,83</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>279.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>73.5,89,75.5,89</points>
<connection>
<GID>302</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>301</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,85.5,77.5,86</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,85.5,77.5,85.5</points>
<intersection>63.5 2</intersection>
<intersection>77.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>63.5,85.5,63.5,98.5</points>
<intersection>85.5 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,90,67.5,90</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>63.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>61.5,98.5,63.5,98.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<intersection>63.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>105,89,107,89</points>
<connection>
<GID>305</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>304</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,86,109,86</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>95,86,95,98.5</points>
<intersection>86 1</intersection>
<intersection>90 4</intersection>
<intersection>98.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95,90,99,90</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>95 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>92.5,98.5,95,98.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>95 2</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>0,46.8715,492.369,-196.497</PageViewport></page 9></circuit>