<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0.624102,593.912,207.407,491.703</PageViewport></page 0>
<page 1>
<PageViewport>-550.8,271.8,673.2,-333.2</PageViewport></page 1>
<page 2>
<PageViewport>-601.579,-2886.97,622.421,-3491.97</PageViewport></page 2>
<page 3>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,5.6566e-007,122.4,-60.5</PageViewport></page 9></circuit>