<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-429.803,89.9354,-185.719,-30.7108</PageViewport>
<gate>
<ID>770</ID>
<type>AA_AND2</type>
<position>-162,63</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>771</ID>
<type>AA_AND2</type>
<position>-170.5,52.5</position>
<input>
<ID>IN_0</ID>476 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>772</ID>
<type>AA_AND2</type>
<position>-162,47.5</position>
<input>
<ID>IN_0</ID>476 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>773</ID>
<type>AA_AND2</type>
<position>-170.5,36</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>774</ID>
<type>AA_AND2</type>
<position>-162,31</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>775</ID>
<type>AA_AND2</type>
<position>-170.5,20</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-276.5,24.5</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>776</ID>
<type>AA_AND2</type>
<position>-162,15</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_AND2</type>
<position>-170.5,4</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>778</ID>
<type>AA_AND2</type>
<position>-162,-1</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-274,19</position>
<gparam>LABEL_TEXT i1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>779</ID>
<type>AA_AND2</type>
<position>-170.5,-12</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-274,14.5</position>
<gparam>LABEL_TEXT i2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>780</ID>
<type>AA_AND2</type>
<position>-162.5,-17</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>-274,10</position>
<gparam>LABEL_TEXT i3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>781</ID>
<type>AA_AND2</type>
<position>-170.5,-27</position>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>782</ID>
<type>AA_AND2</type>
<position>-162,-32</position>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-269.5,5.5</position>
<gparam>LABEL_TEXT input combitaions that is address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>783</ID>
<type>AA_AND2</type>
<position>-170.5,-42.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AA_AND2</type>
<position>-162,-47.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>521 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>786</ID>
<type>BE_DECODER_3x8</type>
<position>-243.5,20</position>
<input>
<ID>ENABLE</ID>625 </input>
<input>
<ID>IN_0</ID>629 </input>
<input>
<ID>IN_1</ID>628 </input>
<input>
<ID>IN_2</ID>626 </input>
<output>
<ID>OUT_0</ID>482 </output>
<output>
<ID>OUT_1</ID>481 </output>
<output>
<ID>OUT_2</ID>480 </output>
<output>
<ID>OUT_3</ID>479 </output>
<output>
<ID>OUT_4</ID>478 </output>
<output>
<ID>OUT_5</ID>477 </output>
<output>
<ID>OUT_6</ID>476 </output>
<output>
<ID>OUT_7</ID>475 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-246.5,-35.5</position>
<gparam>LABEL_TEXT selected register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>788</ID>
<type>AA_TOGGLE</type>
<position>-263.5,19</position>
<output>
<ID>OUT_0</ID>626 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>790</ID>
<type>AA_TOGGLE</type>
<position>-263.5,14.5</position>
<output>
<ID>OUT_0</ID>628 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>792</ID>
<type>AA_TOGGLE</type>
<position>-263.5,11.5</position>
<output>
<ID>OUT_0</ID>629 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>794</ID>
<type>AA_TOGGLE</type>
<position>-272,23.5</position>
<output>
<ID>OUT_0</ID>625 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>-372,4.5</position>
<gparam>LABEL_TEXT WRITE using clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>795</ID>
<type>BA_TRI_STATE</type>
<position>-143,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>483 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>796</ID>
<type>BA_TRI_STATE</type>
<position>-119.5,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>484 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>797</ID>
<type>BA_TRI_STATE</type>
<position>-97,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>485 </input>
<output>
<ID>OUT_0</ID>531 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>798</ID>
<type>BA_TRI_STATE</type>
<position>-76.5,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>486 </input>
<output>
<ID>OUT_0</ID>533 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>799</ID>
<type>BA_TRI_STATE</type>
<position>-55,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>487 </input>
<output>
<ID>OUT_0</ID>535 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>800</ID>
<type>BA_TRI_STATE</type>
<position>-33.5,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>537 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>801</ID>
<type>BA_TRI_STATE</type>
<position>-12,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>489 </input>
<output>
<ID>OUT_0</ID>539 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>802</ID>
<type>BA_TRI_STATE</type>
<position>8,-64</position>
<input>
<ID>ENABLE_0</ID>491 </input>
<input>
<ID>IN_0</ID>490 </input>
<output>
<ID>OUT_0</ID>541 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>803</ID>
<type>BA_TRI_STATE</type>
<position>-123.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>492 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>-371,35.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>804</ID>
<type>BA_TRI_STATE</type>
<position>-100,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>530 </input>
<output>
<ID>OUT_0</ID>493 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>-361.5,35.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>805</ID>
<type>BA_TRI_STATE</type>
<position>-78.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>532 </input>
<output>
<ID>OUT_0</ID>494 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>806</ID>
<type>BA_TRI_STATE</type>
<position>-57.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>534 </input>
<output>
<ID>OUT_0</ID>495 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>-384.5,36.5</position>
<gparam>LABEL_TEXT without delay</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>807</ID>
<type>BA_TRI_STATE</type>
<position>-36,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>536 </input>
<output>
<ID>OUT_0</ID>496 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>808</ID>
<type>BA_TRI_STATE</type>
<position>-14.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>538 </input>
<output>
<ID>OUT_0</ID>497 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>809</ID>
<type>BA_TRI_STATE</type>
<position>6,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>540 </input>
<output>
<ID>OUT_0</ID>498 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>810</ID>
<type>BA_TRI_STATE</type>
<position>30.5,93.5</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>542 </input>
<output>
<ID>OUT_0</ID>499 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>812</ID>
<type>DA_FROM</type>
<position>-143,-73</position>
<input>
<ID>IN_0</ID>483 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>814</ID>
<type>DA_FROM</type>
<position>-119.5,-73</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>823</ID>
<type>DA_FROM</type>
<position>-97,-72</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>824</ID>
<type>DA_FROM</type>
<position>-76.5,-73</position>
<input>
<ID>IN_0</ID>486 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>825</ID>
<type>DA_FROM</type>
<position>-55,-72.5</position>
<input>
<ID>IN_0</ID>487 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>826</ID>
<type>DA_FROM</type>
<position>-33.5,-73</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>827</ID>
<type>DA_FROM</type>
<position>-12,-72.5</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>828</ID>
<type>DA_FROM</type>
<position>8,-71.5</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>829</ID>
<type>DA_FROM</type>
<position>-160.5,-64</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>831</ID>
<type>DA_FROM</type>
<position>-145,93</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>-184,92.5</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>835</ID>
<type>DE_TO</type>
<position>-126,107.5</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>836</ID>
<type>DE_TO</type>
<position>-103,107.5</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>837</ID>
<type>DE_TO</type>
<position>-80,107.5</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>838</ID>
<type>DE_TO</type>
<position>-59.5,108</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>839</ID>
<type>DE_TO</type>
<position>-38,108</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>840</ID>
<type>DE_TO</type>
<position>-16.5,108.5</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>841</ID>
<type>DE_TO</type>
<position>5,108</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>842</ID>
<type>DE_TO</type>
<position>25,107.5</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>844</ID>
<type>DA_FROM</type>
<position>-187,-65.5</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>846</ID>
<type>AA_TOGGLE</type>
<position>-370,29</position>
<output>
<ID>OUT_0</ID>606 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>847</ID>
<type>AA_TOGGLE</type>
<position>-370,21.5</position>
<output>
<ID>OUT_0</ID>607 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>848</ID>
<type>AA_TOGGLE</type>
<position>-370,14.5</position>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>849</ID>
<type>AA_TOGGLE</type>
<position>-352,-3.5</position>
<output>
<ID>OUT_0</ID>609 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>850</ID>
<type>AA_TOGGLE</type>
<position>-344,-3.5</position>
<output>
<ID>OUT_0</ID>610 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>851</ID>
<type>AA_TOGGLE</type>
<position>-337,-3</position>
<output>
<ID>OUT_0</ID>611 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>852</ID>
<type>AA_TOGGLE</type>
<position>-331,-2.5</position>
<output>
<ID>OUT_0</ID>612 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>853</ID>
<type>AA_TOGGLE</type>
<position>-325,-3.5</position>
<output>
<ID>OUT_0</ID>613 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>854</ID>
<type>AA_TOGGLE</type>
<position>-319,-3.5</position>
<output>
<ID>OUT_0</ID>614 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>855</ID>
<type>AA_TOGGLE</type>
<position>-313,-3</position>
<output>
<ID>OUT_0</ID>615 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>856</ID>
<type>AA_TOGGLE</type>
<position>-306,-3</position>
<output>
<ID>OUT_0</ID>616 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>858</ID>
<type>GA_LED</type>
<position>-355,43</position>
<input>
<ID>N_in3</ID>617 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>861</ID>
<type>GA_LED</type>
<position>-346.5,43</position>
<input>
<ID>N_in3</ID>618 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>862</ID>
<type>GA_LED</type>
<position>-339,43</position>
<input>
<ID>N_in3</ID>619 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>863</ID>
<type>GA_LED</type>
<position>-333,43</position>
<input>
<ID>N_in3</ID>620 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>864</ID>
<type>GA_LED</type>
<position>-326.5,43</position>
<input>
<ID>N_in3</ID>621 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>865</ID>
<type>GA_LED</type>
<position>-320.5,43</position>
<input>
<ID>N_in3</ID>622 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>866</ID>
<type>GA_LED</type>
<position>-313.5,43</position>
<input>
<ID>N_in3</ID>623 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>867</ID>
<type>GA_LED</type>
<position>-308,43</position>
<input>
<ID>N_in3</ID>624 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>869</ID>
<type>DE_TO</type>
<position>-363,29</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>871</ID>
<type>DE_TO</type>
<position>-362,21.5</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>872</ID>
<type>DE_TO</type>
<position>-362,14.5</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>873</ID>
<type>DE_TO</type>
<position>-352,6</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>874</ID>
<type>DE_TO</type>
<position>-344,6</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>875</ID>
<type>DE_TO</type>
<position>-337,6</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>876</ID>
<type>DE_TO</type>
<position>-331,6</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>877</ID>
<type>DE_TO</type>
<position>-325,6.5</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>878</ID>
<type>DE_TO</type>
<position>-319,6</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>879</ID>
<type>DE_TO</type>
<position>-313,6</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>880</ID>
<type>DE_TO</type>
<position>-306,6</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>882</ID>
<type>DA_FROM</type>
<position>-355,54</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>883</ID>
<type>DA_FROM</type>
<position>-346.5,53.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>884</ID>
<type>DA_FROM</type>
<position>-339,53.5</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>885</ID>
<type>DA_FROM</type>
<position>-333,54</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>886</ID>
<type>DA_FROM</type>
<position>-326.5,54</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>887</ID>
<type>DA_FROM</type>
<position>-320.5,54</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>888</ID>
<type>DA_FROM</type>
<position>-313.5,54</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>889</ID>
<type>DA_FROM</type>
<position>-308,54</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>895</ID>
<type>AA_LABEL</type>
<position>-357,67</position>
<gparam>LABEL_TEXT OUTPUT READ HERE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-258.5,52.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>88 </input>
<input>
<ID>IN_3</ID>87 </input>
<input>
<ID>IN_4</ID>86 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>84 </input>
<input>
<ID>IN_7</ID>83 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>-278.5,61</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L1</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>-278.5,58.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L2</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>-278.5,56</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L3</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>-278.5,53.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L4</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-278.5,51</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L5</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>-278.5,48</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L6</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>-278.5,45</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L7</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>-278.5,42.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L8</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_TOGGLE</type>
<position>-300,33</position>
<output>
<ID>OUT_0</ID>315 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_DFF_LOW</type>
<position>86.5,3</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>159 </output>
<input>
<ID>clock</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>231</ID>
<type>AE_DFF_LOW</type>
<position>75,3.5</position>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUT_0</ID>160 </output>
<input>
<ID>clock</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>232</ID>
<type>AE_DFF_LOW</type>
<position>121,-8</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>164 </output>
<input>
<ID>clock</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>233</ID>
<type>AE_SMALL_INVERTER</type>
<position>84,21</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>234</ID>
<type>DE_TO</type>
<position>130.5,-6</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L1</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>76,29</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>51,2.5</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>51,0</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>100.5,23.5</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>51,-5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>240</ID>
<type>AI_XOR2</type>
<position>94.5,-1</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AI_XOR2</type>
<position>110.5,-6</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_AND2</type>
<position>110.5,-15</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>94.5,-22</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_OR2</type>
<position>123,-19</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_TOGGLE</type>
<position>70,-10.5</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_AND2</type>
<position>83,12.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_AND2</type>
<position>71.5,11.5</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>165 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AE_DFF_LOW</type>
<position>175,3</position>
<input>
<ID>IN_0</ID>173 </input>
<output>
<ID>OUT_0</ID>175 </output>
<input>
<ID>clock</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>249</ID>
<type>AE_DFF_LOW</type>
<position>163.5,3.5</position>
<input>
<ID>IN_0</ID>174 </input>
<output>
<ID>OUT_0</ID>176 </output>
<input>
<ID>clock</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>250</ID>
<type>AE_DFF_LOW</type>
<position>209.5,-8</position>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>180 </output>
<input>
<ID>clock</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>251</ID>
<type>AE_SMALL_INVERTER</type>
<position>172.5,21</position>
<input>
<ID>IN_0</ID>181 </input>
<output>
<ID>OUT_0</ID>178 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>252</ID>
<type>DE_TO</type>
<position>219,-6</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L2</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>164.5,29</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>139.5,2.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>139.5,0</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>189,23.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>139.5,-5</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>258</ID>
<type>AI_XOR2</type>
<position>183,-1</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>259</ID>
<type>AI_XOR2</type>
<position>199,-6</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_AND2</type>
<position>199,-15</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>169 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_AND2</type>
<position>183,-22</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_OR2</type>
<position>211.5,-19</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_AND2</type>
<position>171.5,12.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>179 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>160,11.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_DFF_LOW</type>
<position>265.5,3</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>191 </output>
<input>
<ID>clock</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>267</ID>
<type>AE_DFF_LOW</type>
<position>254,3.5</position>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUT_0</ID>192 </output>
<input>
<ID>clock</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>268</ID>
<type>AE_DFF_LOW</type>
<position>300,-8</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>196 </output>
<input>
<ID>clock</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_SMALL_INVERTER</type>
<position>263,21</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>DE_TO</type>
<position>309.5,-6</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L3</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>255,29</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>230,2.5</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>273</ID>
<type>DA_FROM</type>
<position>230,0</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>274</ID>
<type>DA_FROM</type>
<position>279.5,23.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>275</ID>
<type>DA_FROM</type>
<position>230,-5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>276</ID>
<type>AI_XOR2</type>
<position>273.5,-1</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AI_XOR2</type>
<position>289.5,-6</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>289.5,-15</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_AND2</type>
<position>273.5,-22</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AE_OR2</type>
<position>302,-19</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND2</type>
<position>262,12.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_AND2</type>
<position>250.5,11.5</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>AE_DFF_LOW</type>
<position>353,3</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>207 </output>
<input>
<ID>clock</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>284</ID>
<type>AE_DFF_LOW</type>
<position>341.5,3.5</position>
<input>
<ID>IN_0</ID>206 </input>
<output>
<ID>OUT_0</ID>208 </output>
<input>
<ID>clock</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>285</ID>
<type>AE_DFF_LOW</type>
<position>387.5,-8</position>
<input>
<ID>IN_0</ID>209 </input>
<output>
<ID>OUT_0</ID>212 </output>
<input>
<ID>clock</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_SMALL_INVERTER</type>
<position>350.5,21</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>287</ID>
<type>DE_TO</type>
<position>397,-6</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L4</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>342.5,29</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>317.5,2.5</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>317.5,0</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>367,23.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>292</ID>
<type>DA_FROM</type>
<position>317.5,-5</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>293</ID>
<type>AI_XOR2</type>
<position>361,-1</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>AI_XOR2</type>
<position>377,-6</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_AND2</type>
<position>377,-15</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND2</type>
<position>361,-22</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>AE_OR2</type>
<position>389.5,-19</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND2</type>
<position>349.5,12.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>338,11.5</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_DFF_LOW</type>
<position>440,3</position>
<input>
<ID>IN_0</ID>221 </input>
<output>
<ID>OUT_0</ID>223 </output>
<input>
<ID>clock</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>301</ID>
<type>AE_DFF_LOW</type>
<position>428.5,3.5</position>
<input>
<ID>IN_0</ID>222 </input>
<output>
<ID>OUT_0</ID>224 </output>
<input>
<ID>clock</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_DFF_LOW</type>
<position>474.5,-8</position>
<input>
<ID>IN_0</ID>225 </input>
<output>
<ID>OUT_0</ID>228 </output>
<input>
<ID>clock</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_SMALL_INVERTER</type>
<position>437.5,21</position>
<input>
<ID>IN_0</ID>229 </input>
<output>
<ID>OUT_0</ID>226 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>304</ID>
<type>DE_TO</type>
<position>484,-6</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L5</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>429.5,29</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q5</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>404.5,2.5</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>404.5,0</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>454,23.5</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>404.5,-5</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>310</ID>
<type>AI_XOR2</type>
<position>448,-1</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>AI_XOR2</type>
<position>464,-6</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_AND2</type>
<position>464,-15</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>448,-22</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>AE_OR2</type>
<position>476.5,-19</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_AND2</type>
<position>436.5,12.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>425,11.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>AE_DFF_LOW</type>
<position>526,2.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>239 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_DFF_LOW</type>
<position>514.5,3</position>
<input>
<ID>IN_0</ID>238 </input>
<output>
<ID>OUT_0</ID>240 </output>
<input>
<ID>clock</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_DFF_LOW</type>
<position>560.5,-8.5</position>
<input>
<ID>IN_0</ID>241 </input>
<output>
<ID>OUT_0</ID>244 </output>
<input>
<ID>clock</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_SMALL_INVERTER</type>
<position>523.5,20.5</position>
<input>
<ID>IN_0</ID>245 </input>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>321</ID>
<type>DE_TO</type>
<position>570,-6.5</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L6</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>515.5,28.5</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q6</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>490.5,2</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>324</ID>
<type>DA_FROM</type>
<position>490.5,-0.5</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>540,23</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>490.5,-5.5</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>327</ID>
<type>AI_XOR2</type>
<position>534,-1.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>AI_XOR2</type>
<position>550,-6.5</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_AND2</type>
<position>550,-15.5</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AA_AND2</type>
<position>534,-22.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AE_OR2</type>
<position>562.5,-19.5</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_AND2</type>
<position>522.5,12</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AA_AND2</type>
<position>511,11</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>245 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>351</ID>
<type>AE_DFF_LOW</type>
<position>616.5,3.5</position>
<input>
<ID>IN_0</ID>269 </input>
<output>
<ID>OUT_0</ID>271 </output>
<input>
<ID>clock</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>352</ID>
<type>AE_DFF_LOW</type>
<position>605,4</position>
<input>
<ID>IN_0</ID>270 </input>
<output>
<ID>OUT_0</ID>272 </output>
<input>
<ID>clock</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_DFF_LOW</type>
<position>651,-7.5</position>
<input>
<ID>IN_0</ID>273 </input>
<output>
<ID>OUT_0</ID>276 </output>
<input>
<ID>clock</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>354</ID>
<type>AE_SMALL_INVERTER</type>
<position>614,21.5</position>
<input>
<ID>IN_0</ID>277 </input>
<output>
<ID>OUT_0</ID>274 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>660.5,-5.5</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L7</lparam></gate>
<gate>
<ID>356</ID>
<type>DA_FROM</type>
<position>606,29.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q7</lparam></gate>
<gate>
<ID>357</ID>
<type>DA_FROM</type>
<position>581,3</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>581,0.5</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>630.5,24</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>581,-4.5</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>361</ID>
<type>AI_XOR2</type>
<position>624.5,-0.5</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>AI_XOR2</type>
<position>640.5,-5.5</position>
<input>
<ID>IN_0</ID>265 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>640.5,-14.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>AA_AND2</type>
<position>624.5,-21.5</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_OR2</type>
<position>653,-18.5</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>266 </input>
<output>
<ID>OUT</ID>300 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>366</ID>
<type>AA_AND2</type>
<position>613,13</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>269 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_AND2</type>
<position>601.5,12</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>277 </input>
<output>
<ID>OUT</ID>270 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>AE_DFF_LOW</type>
<position>704,5</position>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>303 </output>
<input>
<ID>clock</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>386</ID>
<type>AE_DFF_LOW</type>
<position>692.5,5.5</position>
<input>
<ID>IN_0</ID>302 </input>
<output>
<ID>OUT_0</ID>304 </output>
<input>
<ID>clock</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>387</ID>
<type>AE_DFF_LOW</type>
<position>738.5,-6</position>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>308 </output>
<input>
<ID>clock</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>388</ID>
<type>AE_SMALL_INVERTER</type>
<position>701.5,23</position>
<input>
<ID>IN_0</ID>309 </input>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>389</ID>
<type>DE_TO</type>
<position>748,-4</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L8</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>693.5,31</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q8</lparam></gate>
<gate>
<ID>391</ID>
<type>DA_FROM</type>
<position>668.5,4.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>392</ID>
<type>DA_FROM</type>
<position>668.5,2</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>718,25.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>394</ID>
<type>DA_FROM</type>
<position>668.5,-3</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>395</ID>
<type>AI_XOR2</type>
<position>712,1</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>297 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>AI_XOR2</type>
<position>728,-4</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>300 </input>
<output>
<ID>OUT</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_AND2</type>
<position>728,-13</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>297 </input>
<output>
<ID>OUT</ID>299 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_AND2</type>
<position>712,-20</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>298 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>AE_OR2</type>
<position>740.5,-17</position>
<input>
<ID>IN_0</ID>299 </input>
<input>
<ID>IN_1</ID>298 </input>
<output>
<ID>OUT</ID>313 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>AA_AND2</type>
<position>700.5,14.5</position>
<input>
<ID>IN_0</ID>306 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>AA_AND2</type>
<position>689,13.5</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>309 </input>
<output>
<ID>OUT</ID>302 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>DE_TO</type>
<position>753,-17</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CARRY</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_TOGGLE</type>
<position>-300,29</position>
<output>
<ID>OUT_0</ID>318 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_TOGGLE</type>
<position>-300,25.5</position>
<output>
<ID>OUT_0</ID>317 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_TOGGLE</type>
<position>-300,21.5</position>
<output>
<ID>OUT_0</ID>316 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>408</ID>
<type>GA_LED</type>
<position>-255.5,36.5</position>
<input>
<ID>N_in0</ID>314 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>-268,36.5</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CARRY</lparam></gate>
<gate>
<ID>412</ID>
<type>DE_TO</type>
<position>-293.5,33</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>413</ID>
<type>DE_TO</type>
<position>-293,29</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>414</ID>
<type>DE_TO</type>
<position>-293,25.5</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>415</ID>
<type>DE_TO</type>
<position>-293,21.5</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>638</ID>
<type>AE_DFF_LOW</type>
<position>-136,69</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>578 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>639</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,69</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>573 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>640</ID>
<type>AE_DFF_LOW</type>
<position>-90,69</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>572 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_DFF_LOW</type>
<position>-71,69</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>563 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>642</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,69</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>562 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>643</ID>
<type>AE_DFF_LOW</type>
<position>-27,69</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>553 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>644</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,69</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>545 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_DFF_LOW</type>
<position>14.5,69</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>543 </output>
<input>
<ID>clock</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>647</ID>
<type>BA_TRI_STATE</type>
<position>-129,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>578 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>648</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>573 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>649</ID>
<type>BA_TRI_STATE</type>
<position>-83,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>572 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>650</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>563 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>651</ID>
<type>BA_TRI_STATE</type>
<position>-41,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>562 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>652</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>553 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>653</ID>
<type>BA_TRI_STATE</type>
<position>2,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>545 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>654</ID>
<type>BA_TRI_STATE</type>
<position>22,63</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>543 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>655</ID>
<type>AE_DFF_LOW</type>
<position>-136,53.5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>579 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>656</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,53.5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>574 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>657</ID>
<type>AE_DFF_LOW</type>
<position>-90,53.5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>571 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>658</ID>
<type>AE_DFF_LOW</type>
<position>-71,53.5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>564 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>659</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,53.5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>561 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>660</ID>
<type>AE_DFF_LOW</type>
<position>-27,53.5</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>554 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>661</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,53.5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>546 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>662</ID>
<type>AE_DFF_LOW</type>
<position>14.5,53.5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>544 </output>
<input>
<ID>clock</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>663</ID>
<type>BA_TRI_STATE</type>
<position>-129,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>579 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>664</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>574 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>665</ID>
<type>BA_TRI_STATE</type>
<position>-83,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>571 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>666</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>564 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>667</ID>
<type>BA_TRI_STATE</type>
<position>-41,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>668</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>554 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>669</ID>
<type>BA_TRI_STATE</type>
<position>2,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>546 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>670</ID>
<type>BA_TRI_STATE</type>
<position>22,47.5</position>
<input>
<ID>ENABLE_0</ID>505 </input>
<input>
<ID>IN_0</ID>544 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>671</ID>
<type>AE_DFF_LOW</type>
<position>-136,37</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>582 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>672</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,37</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>575 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>673</ID>
<type>AE_DFF_LOW</type>
<position>-90,37</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>570 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>674</ID>
<type>AE_DFF_LOW</type>
<position>-71,37</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>565 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>675</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,37</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>560 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>676</ID>
<type>AE_DFF_LOW</type>
<position>-27,37</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>555 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>677</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,37</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>550 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>678</ID>
<type>AE_DFF_LOW</type>
<position>14.5,37</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>549 </output>
<input>
<ID>clock</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>679</ID>
<type>BA_TRI_STATE</type>
<position>-129,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>582 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>680</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>575 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>681</ID>
<type>BA_TRI_STATE</type>
<position>-83,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>570 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>682</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>565 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>683</ID>
<type>BA_TRI_STATE</type>
<position>-41,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>560 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>684</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>555 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>685</ID>
<type>BA_TRI_STATE</type>
<position>2,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>550 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>686</ID>
<type>BA_TRI_STATE</type>
<position>22,31</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>549 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_DFF_LOW</type>
<position>-136,21</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>581 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>688</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,21</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>576 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>689</ID>
<type>AE_DFF_LOW</type>
<position>-90,21</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>569 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_DFF_LOW</type>
<position>-71,21</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>566 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>691</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,21</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>559 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_DFF_LOW</type>
<position>-27,21</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>556 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>693</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,21</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>551 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>694</ID>
<type>AE_DFF_LOW</type>
<position>14.5,21</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>548 </output>
<input>
<ID>clock</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>695</ID>
<type>BA_TRI_STATE</type>
<position>-129,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>581 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>696</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>576 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>697</ID>
<type>BA_TRI_STATE</type>
<position>-83,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>569 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>698</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>566 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>699</ID>
<type>BA_TRI_STATE</type>
<position>-41,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>559 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>700</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>556 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>701</ID>
<type>BA_TRI_STATE</type>
<position>2,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>551 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>702</ID>
<type>BA_TRI_STATE</type>
<position>22,15</position>
<input>
<ID>ENABLE_0</ID>510 </input>
<input>
<ID>IN_0</ID>548 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>703</ID>
<type>AE_DFF_LOW</type>
<position>-136,5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>580 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>704</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>577 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>705</ID>
<type>AE_DFF_LOW</type>
<position>-90,5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>568 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>706</ID>
<type>AE_DFF_LOW</type>
<position>-71,5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>567 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>707</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>558 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>708</ID>
<type>AE_DFF_LOW</type>
<position>-27,5</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>557 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>709</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>552 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>710</ID>
<type>AE_DFF_LOW</type>
<position>14.5,5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>547 </output>
<input>
<ID>clock</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>711</ID>
<type>BA_TRI_STATE</type>
<position>-129,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>580 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>712</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>577 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>713</ID>
<type>BA_TRI_STATE</type>
<position>-83,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>568 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>714</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>567 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>715</ID>
<type>BA_TRI_STATE</type>
<position>-41,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>558 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>716</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>557 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>717</ID>
<type>BA_TRI_STATE</type>
<position>2,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>552 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>718</ID>
<type>BA_TRI_STATE</type>
<position>22,-1</position>
<input>
<ID>ENABLE_0</ID>512 </input>
<input>
<ID>IN_0</ID>547 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>719</ID>
<type>AE_DFF_LOW</type>
<position>-136,-11</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>583 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>720</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,-11</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>586 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>721</ID>
<type>AE_DFF_LOW</type>
<position>-90,-11</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>587 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>722</ID>
<type>AE_DFF_LOW</type>
<position>-71,-11</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>591 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>723</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,-11</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>596 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>724</ID>
<type>AE_DFF_LOW</type>
<position>-27,-11</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>597 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>725</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,-11</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>601 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>726</ID>
<type>AE_DFF_LOW</type>
<position>14.5,-11</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>603 </output>
<input>
<ID>clock</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>727</ID>
<type>BA_TRI_STATE</type>
<position>-129,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>583 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>728</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>586 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>729</ID>
<type>BA_TRI_STATE</type>
<position>-83,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>587 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>730</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>591 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>731</ID>
<type>BA_TRI_STATE</type>
<position>-41,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>596 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>732</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>597 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>733</ID>
<type>BA_TRI_STATE</type>
<position>2,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>601 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>734</ID>
<type>BA_TRI_STATE</type>
<position>22,-17</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>735</ID>
<type>AE_DFF_LOW</type>
<position>-136,-26</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>523 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>736</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,-26</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>585 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>737</ID>
<type>AE_DFF_LOW</type>
<position>-90,-26</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>590 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>738</ID>
<type>AE_DFF_LOW</type>
<position>-71,-26</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>593 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>739</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,-26</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>594 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>740</ID>
<type>AE_DFF_LOW</type>
<position>-27,-26</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>598 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>741</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,-26</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>600 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>742</ID>
<type>AE_DFF_LOW</type>
<position>14.5,-26</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>604 </output>
<input>
<ID>clock</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>743</ID>
<type>BA_TRI_STATE</type>
<position>-129,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>523 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>744</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>585 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>745</ID>
<type>BA_TRI_STATE</type>
<position>-83,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>590 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>746</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>593 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>747</ID>
<type>BA_TRI_STATE</type>
<position>-41,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>594 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>748</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>598 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>749</ID>
<type>BA_TRI_STATE</type>
<position>2,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>600 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>750</ID>
<type>BA_TRI_STATE</type>
<position>22,-32</position>
<input>
<ID>ENABLE_0</ID>522 </input>
<input>
<ID>IN_0</ID>604 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_DFF_LOW</type>
<position>-136,-41.5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>524 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>752</ID>
<type>AE_DFF_LOW</type>
<position>-113.5,-41.5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>584 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>753</ID>
<type>AE_DFF_LOW</type>
<position>-90,-41.5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>589 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>754</ID>
<type>AE_DFF_LOW</type>
<position>-71,-41.5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>592 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>755</ID>
<type>AE_DFF_LOW</type>
<position>-48.5,-41.5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>595 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>756</ID>
<type>AE_DFF_LOW</type>
<position>-27,-41.5</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>599 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>757</ID>
<type>AE_DFF_LOW</type>
<position>-5.5,-41.5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>602 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>758</ID>
<type>AE_DFF_LOW</type>
<position>14.5,-41.5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>605 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>759</ID>
<type>BA_TRI_STATE</type>
<position>-129,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>760</ID>
<type>BA_TRI_STATE</type>
<position>-105.5,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>584 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>761</ID>
<type>BA_TRI_STATE</type>
<position>-83,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>589 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>762</ID>
<type>BA_TRI_STATE</type>
<position>-62.5,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>592 </input>
<output>
<ID>OUT_0</ID>534 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>763</ID>
<type>BA_TRI_STATE</type>
<position>-41,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>595 </input>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>764</ID>
<type>BA_TRI_STATE</type>
<position>-19.5,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>599 </input>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>765</ID>
<type>BA_TRI_STATE</type>
<position>2,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>602 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>766</ID>
<type>BA_TRI_STATE</type>
<position>22,-47.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>605 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>768</ID>
<type>AA_AND2</type>
<position>-170.5,68</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>503 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-369,35.5,-363.5,35.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-276.5,61,-267,61</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-267 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-267,56.5,-267,61</points>
<intersection>56.5 7</intersection>
<intersection>61 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-267,56.5,-263.5,56.5</points>
<connection>
<GID>129</GID>
<name>IN_7</name></connection>
<intersection>-267 6</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,55.5,-268,58.5</points>
<intersection>55.5 1</intersection>
<intersection>58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268,55.5,-263.5,55.5</points>
<connection>
<GID>129</GID>
<name>IN_6</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-276.5,58.5,-268,58.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-270,54.5,-263.5,54.5</points>
<connection>
<GID>129</GID>
<name>IN_5</name></connection>
<intersection>-270 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-270,54.5,-270,56</points>
<intersection>54.5 1</intersection>
<intersection>56 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-276.5,56,-270,56</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-270 5</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-229.5,23.5,-229.5,69</points>
<intersection>23.5 2</intersection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-229.5,69,-173.5,69</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>-229.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,23.5,-229.5,23.5</points>
<connection>
<GID>786</GID>
<name>OUT_7</name></connection>
<intersection>-229.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,64,-178,69</points>
<intersection>64 4</intersection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,64,-165,64</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-276.5,53.5,-263.5,53.5</points>
<connection>
<GID>129</GID>
<name>IN_4</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227.5,22.5,-227.5,53.5</points>
<intersection>22.5 2</intersection>
<intersection>53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-227.5,53.5,-173.5,53.5</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<intersection>-227.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,22.5,-227.5,22.5</points>
<connection>
<GID>786</GID>
<name>OUT_6</name></connection>
<intersection>-227.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,48.5,-178,53.5</points>
<intersection>48.5 4</intersection>
<intersection>53.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,48.5,-165,48.5</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-270,51,-270,52.5</points>
<intersection>51 2</intersection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-270,52.5,-263.5,52.5</points>
<connection>
<GID>129</GID>
<name>IN_3</name></connection>
<intersection>-270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-276.5,51,-270,51</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-270 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224.5,21.5,-224.5,37</points>
<intersection>21.5 2</intersection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-224.5,37,-173.5,37</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>-224.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,21.5,-224.5,21.5</points>
<connection>
<GID>786</GID>
<name>OUT_5</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,32,-178,37</points>
<intersection>32 4</intersection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,32,-165,32</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-269,48,-269,51.5</points>
<intersection>48 2</intersection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-269,51.5,-263.5,51.5</points>
<connection>
<GID>129</GID>
<name>IN_2</name></connection>
<intersection>-269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-276.5,48,-269,48</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-269 0</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-240.5,21,-173.5,21</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>-240.5 6</intersection>
<intersection>-178 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,16,-178,21</points>
<intersection>16 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,16,-165,16</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-240.5,20.5,-240.5,21</points>
<connection>
<GID>786</GID>
<name>OUT_4</name></connection>
<intersection>21 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,45,-268,50.5</points>
<intersection>45 2</intersection>
<intersection>50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268,50.5,-263.5,50.5</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-276.5,45,-268,45</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224,5,-224,19.5</points>
<intersection>5 1</intersection>
<intersection>19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-224,5,-173.5,5</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>-224 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,19.5,-224,19.5</points>
<connection>
<GID>786</GID>
<name>OUT_3</name></connection>
<intersection>-224 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,0,-178,5</points>
<intersection>0 4</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,0,-165,0</points>
<connection>
<GID>778</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-267,42.5,-267,49.5</points>
<intersection>42.5 2</intersection>
<intersection>49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-267,49.5,-263.5,49.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-267 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-276.5,42.5,-267,42.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-267 0</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227.5,-11,-227.5,18.5</points>
<intersection>-11 1</intersection>
<intersection>18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-227.5,-11,-173.5,-11</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-227.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,18.5,-227.5,18.5</points>
<connection>
<GID>786</GID>
<name>OUT_2</name></connection>
<intersection>-227.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,-16,-178,-11</points>
<intersection>-16 4</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,-16,-165.5,-16</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230,-26,-230,17.5</points>
<intersection>-26 1</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230,-26,-173.5,-26</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>-230 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,17.5,-230,17.5</points>
<connection>
<GID>786</GID>
<name>OUT_1</name></connection>
<intersection>-230 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,-31,-178,-26</points>
<intersection>-31 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,-31,-165,-31</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233.5,-41.5,-233.5,16.5</points>
<intersection>-41.5 1</intersection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233.5,-41.5,-173.5,-41.5</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>-233.5 0</intersection>
<intersection>-178 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-240.5,16.5,-233.5,16.5</points>
<connection>
<GID>786</GID>
<name>OUT_0</name></connection>
<intersection>-233.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-178,-46.5,-178,-41.5</points>
<intersection>-46.5 4</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-178,-46.5,-165,-46.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>-178 3</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143,-71,-143,-67</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<connection>
<GID>812</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-119.5,-71,-119.5,-67</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<connection>
<GID>814</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97,-70,-97,-67</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<connection>
<GID>823</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-71,-76.5,-67</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<connection>
<GID>824</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-70.5,-55,-67</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<connection>
<GID>825</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-71,-33.5,-67</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<connection>
<GID>826</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-70.5,-12,-67</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<connection>
<GID>827</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-69.5,8,-67</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<connection>
<GID>828</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-158.5,-64,6,-64</points>
<connection>
<GID>797</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>802</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>801</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>800</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>799</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>798</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>796</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>795</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>829</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-123.5,96,-123.5,105.5</points>
<connection>
<GID>803</GID>
<name>OUT_0</name></connection>
<intersection>105.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-126,105.5,-123.5,105.5</points>
<connection>
<GID>835</GID>
<name>IN_0</name></connection>
<intersection>-123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,96,-100,105.5</points>
<connection>
<GID>804</GID>
<name>OUT_0</name></connection>
<intersection>105.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103,105.5,-100,105.5</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>-100 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,96,-78.5,105.5</points>
<connection>
<GID>805</GID>
<name>OUT_0</name></connection>
<intersection>105.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-80,105.5,-78.5,105.5</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,96,-57.5,106</points>
<connection>
<GID>806</GID>
<name>OUT_0</name></connection>
<intersection>106 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-59.5,106,-57.5,106</points>
<connection>
<GID>838</GID>
<name>IN_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,96,-36,106</points>
<connection>
<GID>807</GID>
<name>OUT_0</name></connection>
<intersection>106 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-38,106,-36,106</points>
<connection>
<GID>839</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,96,-14.5,106.5</points>
<connection>
<GID>808</GID>
<name>OUT_0</name></connection>
<intersection>106.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-16.5,106.5,-14.5,106.5</points>
<connection>
<GID>840</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,96,6,106</points>
<connection>
<GID>809</GID>
<name>OUT_0</name></connection>
<intersection>106 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>5,106,6,106</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,96,30.5,105.5</points>
<connection>
<GID>810</GID>
<name>OUT_0</name></connection>
<intersection>105.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>25,105.5,30.5,105.5</points>
<connection>
<GID>842</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-143,93.5,28.5,93.5</points>
<connection>
<GID>809</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>807</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>803</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>804</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>805</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>806</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>808</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>810</GID>
<name>ENABLE_0</name></connection>
<intersection>-143 34</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>-143,93,-143,93.5</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>93.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-187,-63.5,-187,67</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>-43.5 8</intersection>
<intersection>-28 7</intersection>
<intersection>-13 6</intersection>
<intersection>3 5</intersection>
<intersection>19 4</intersection>
<intersection>35 3</intersection>
<intersection>51.5 2</intersection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-187,67,-173.5,67</points>
<connection>
<GID>768</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-187,51.5,-173.5,51.5</points>
<connection>
<GID>771</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-187,35,-173.5,35</points>
<connection>
<GID>773</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-187,19,-173.5,19</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-187,3,-173.5,3</points>
<connection>
<GID>777</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-187,-13,-173.5,-13</points>
<connection>
<GID>779</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-187,-28,-173.5,-28</points>
<connection>
<GID>781</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-187,-43.5,-173.5,-43.5</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>-187 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-182,-48.5,-182,90.5</points>
<intersection>-48.5 1</intersection>
<intersection>-33 3</intersection>
<intersection>-18 5</intersection>
<intersection>-2 7</intersection>
<intersection>14 9</intersection>
<intersection>30 10</intersection>
<intersection>46.5 11</intersection>
<intersection>62 12</intersection>
<intersection>90.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-182,-48.5,-165,-48.5</points>
<connection>
<GID>784</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-182,-33,-165,-33</points>
<connection>
<GID>782</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-182,-18,-165.5,-18</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-182,-2,-165,-2</points>
<connection>
<GID>778</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-184,90.5,-182,90.5</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-182,14,-165,14</points>
<connection>
<GID>776</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-182,30,-165,30</points>
<connection>
<GID>774</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-182,46.5,-165,46.5</points>
<connection>
<GID>772</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-182,62,-165,62</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<intersection>-182 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,68,11.5,68</points>
<connection>
<GID>645</GID>
<name>clock</name></connection>
<connection>
<GID>644</GID>
<name>clock</name></connection>
<connection>
<GID>643</GID>
<name>clock</name></connection>
<connection>
<GID>642</GID>
<name>clock</name></connection>
<connection>
<GID>641</GID>
<name>clock</name></connection>
<connection>
<GID>640</GID>
<name>clock</name></connection>
<connection>
<GID>639</GID>
<name>clock</name></connection>
<connection>
<GID>638</GID>
<name>clock</name></connection>
<connection>
<GID>768</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,63,20,63</points>
<connection>
<GID>654</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>653</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>652</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>651</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>650</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>649</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>648</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>647</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>770</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,47.5,20,47.5</points>
<connection>
<GID>772</GID>
<name>OUT</name></connection>
<connection>
<GID>663</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>664</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>665</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>666</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>667</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>668</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>669</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>670</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,52.5,11.5,52.5</points>
<connection>
<GID>771</GID>
<name>OUT</name></connection>
<connection>
<GID>655</GID>
<name>clock</name></connection>
<connection>
<GID>656</GID>
<name>clock</name></connection>
<connection>
<GID>657</GID>
<name>clock</name></connection>
<connection>
<GID>658</GID>
<name>clock</name></connection>
<connection>
<GID>659</GID>
<name>clock</name></connection>
<connection>
<GID>660</GID>
<name>clock</name></connection>
<connection>
<GID>662</GID>
<name>clock</name></connection>
<connection>
<GID>661</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,36,11.5,36</points>
<connection>
<GID>678</GID>
<name>clock</name></connection>
<connection>
<GID>677</GID>
<name>clock</name></connection>
<connection>
<GID>676</GID>
<name>clock</name></connection>
<connection>
<GID>675</GID>
<name>clock</name></connection>
<connection>
<GID>674</GID>
<name>clock</name></connection>
<connection>
<GID>673</GID>
<name>clock</name></connection>
<connection>
<GID>672</GID>
<name>clock</name></connection>
<connection>
<GID>671</GID>
<name>clock</name></connection>
<connection>
<GID>773</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,31,20,31</points>
<connection>
<GID>686</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>685</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>684</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>683</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>682</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>681</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>679</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>774</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,20,11.5,20</points>
<connection>
<GID>775</GID>
<name>OUT</name></connection>
<connection>
<GID>687</GID>
<name>clock</name></connection>
<connection>
<GID>689</GID>
<name>clock</name></connection>
<connection>
<GID>690</GID>
<name>clock</name></connection>
<connection>
<GID>691</GID>
<name>clock</name></connection>
<connection>
<GID>692</GID>
<name>clock</name></connection>
<connection>
<GID>693</GID>
<name>clock</name></connection>
<connection>
<GID>694</GID>
<name>clock</name></connection>
<connection>
<GID>688</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,15,20,15</points>
<connection>
<GID>776</GID>
<name>OUT</name></connection>
<connection>
<GID>695</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>696</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>697</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>698</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>699</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>700</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>701</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>702</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,4,11.5,4</points>
<connection>
<GID>710</GID>
<name>clock</name></connection>
<connection>
<GID>709</GID>
<name>clock</name></connection>
<connection>
<GID>708</GID>
<name>clock</name></connection>
<connection>
<GID>707</GID>
<name>clock</name></connection>
<connection>
<GID>706</GID>
<name>clock</name></connection>
<connection>
<GID>705</GID>
<name>clock</name></connection>
<connection>
<GID>704</GID>
<name>clock</name></connection>
<connection>
<GID>777</GID>
<name>OUT</name></connection>
<connection>
<GID>703</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-159,-1,20,-1</points>
<connection>
<GID>718</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>717</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>716</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>715</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>714</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>713</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>712</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>778</GID>
<name>OUT</name></connection>
<connection>
<GID>711</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,-12,11.5,-12</points>
<connection>
<GID>779</GID>
<name>OUT</name></connection>
<connection>
<GID>719</GID>
<name>clock</name></connection>
<connection>
<GID>720</GID>
<name>clock</name></connection>
<connection>
<GID>721</GID>
<name>clock</name></connection>
<connection>
<GID>722</GID>
<name>clock</name></connection>
<connection>
<GID>723</GID>
<name>clock</name></connection>
<connection>
<GID>724</GID>
<name>clock</name></connection>
<connection>
<GID>725</GID>
<name>clock</name></connection>
<connection>
<GID>726</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159.5,-17,20,-17</points>
<connection>
<GID>780</GID>
<name>OUT</name></connection>
<connection>
<GID>727</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>728</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>729</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>730</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>731</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>732</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>733</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>734</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,-27,11.5,-27</points>
<connection>
<GID>735</GID>
<name>clock</name></connection>
<connection>
<GID>781</GID>
<name>OUT</name></connection>
<connection>
<GID>736</GID>
<name>clock</name></connection>
<connection>
<GID>737</GID>
<name>clock</name></connection>
<connection>
<GID>738</GID>
<name>clock</name></connection>
<connection>
<GID>739</GID>
<name>clock</name></connection>
<connection>
<GID>740</GID>
<name>clock</name></connection>
<connection>
<GID>742</GID>
<name>clock</name></connection>
<connection>
<GID>741</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167.5,-42.5,11.5,-42.5</points>
<connection>
<GID>783</GID>
<name>OUT</name></connection>
<connection>
<GID>751</GID>
<name>clock</name></connection>
<connection>
<GID>752</GID>
<name>clock</name></connection>
<connection>
<GID>753</GID>
<name>clock</name></connection>
<connection>
<GID>754</GID>
<name>clock</name></connection>
<connection>
<GID>755</GID>
<name>clock</name></connection>
<connection>
<GID>756</GID>
<name>clock</name></connection>
<connection>
<GID>757</GID>
<name>clock</name></connection>
<connection>
<GID>758</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,-47.5,20,-47.5</points>
<connection>
<GID>784</GID>
<name>OUT</name></connection>
<connection>
<GID>759</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>760</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>761</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>762</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>763</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>764</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>765</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>766</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-159,-32,20,-32</points>
<connection>
<GID>750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>749</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>748</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>745</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>746</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>744</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>743</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>782</GID>
<name>OUT</name></connection>
<connection>
<GID>747</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,-35,-132.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-24,-132.5,-24</points>
<connection>
<GID>735</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,-35,-129,-35</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,-50.5,-132,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-39.5,-132,-39.5</points>
<connection>
<GID>751</GID>
<name>OUT_0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132,-50.5,-129,-50.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143,-61.5,-143,71</points>
<connection>
<GID>795</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-143,71,-139,71</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-143,55.5,-139,55.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-143,39,-139,39</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-143,23,-139,23</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-143,7,-139,7</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-143,-9,-139,-9</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-143,-24,-139,-24</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-143,-39.5,-139,-39.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>-143 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-123.5,-45,-123.5,90.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 6</intersection>
<intersection>1.5 7</intersection>
<intersection>17.5 8</intersection>
<intersection>33.5 9</intersection>
<intersection>50 10</intersection>
<intersection>65.5 11</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-129,-45,-123.5,-45</points>
<connection>
<GID>759</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-129,-14.5,-123.5,-14.5</points>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-129,1.5,-123.5,1.5</points>
<connection>
<GID>711</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-129,17.5,-123.5,17.5</points>
<connection>
<GID>695</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-129,33.5,-123.5,33.5</points>
<connection>
<GID>679</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-129,50,-123.5,50</points>
<connection>
<GID>663</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-129,65.5,-123.5,65.5</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-129,-29.5,-123.5,-29.5</points>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection>
<intersection>-123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-119.5,-61.5,-119.5,71</points>
<connection>
<GID>796</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 7</intersection>
<intersection>-24 8</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-119.5,71,-116.5,71</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,55.5,-116.5,55.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-119.5,39,-116.5,39</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-119.5,23,-116.5,23</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-119.5,7,-116.5,7</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-119.5,-9,-116.5,-9</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-119.5,-39.5,-116.5,-39.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-119.5,-24,-116.5,-24</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>-119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-45,-100,90.5</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 9</intersection>
<intersection>33.5 8</intersection>
<intersection>50 6</intersection>
<intersection>65.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-105.5,-45,-100,-45</points>
<connection>
<GID>760</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-105.5,50,-100,50</points>
<connection>
<GID>664</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-105.5,65.5,-100,65.5</points>
<connection>
<GID>648</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-105.5,33.5,-100,33.5</points>
<connection>
<GID>680</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-105.5,17.5,-100,17.5</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-105.5,1.5,-100,1.5</points>
<connection>
<GID>712</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-105.5,-14.5,-100,-14.5</points>
<connection>
<GID>728</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-105.5,-29.5,-100,-29.5</points>
<connection>
<GID>744</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97,-61.5,-97,71</points>
<connection>
<GID>797</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-97,71,-93,71</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,55.5,-93,55.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-97,39,-93,39</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-97,23,-93,23</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-97,7,-93,7</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-97,-9,-93,-9</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-97,-24,-93,-24</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-97,-39.5,-93,-39.5</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>-97 0</intersection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,-45,-78.5,90.5</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 7</intersection>
<intersection>1.5 11</intersection>
<intersection>17.5 10</intersection>
<intersection>33.5 8</intersection>
<intersection>50 9</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-83,-45,-78.5,-45</points>
<connection>
<GID>761</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-83,65.5,-78.5,65.5</points>
<connection>
<GID>649</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-83,-14.5,-78.5,-14.5</points>
<connection>
<GID>729</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-83,33.5,-78.5,33.5</points>
<connection>
<GID>681</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-83,50,-78.5,50</points>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-83,17.5,-78.5,17.5</points>
<connection>
<GID>697</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-83,1.5,-78.5,1.5</points>
<connection>
<GID>713</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-83,-29.5,-78.5,-29.5</points>
<connection>
<GID>745</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-61.5,-76.5,71</points>
<connection>
<GID>798</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 2</intersection>
<intersection>55.5 3</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,71,-74,71</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76.5,39,-74,39</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-76.5,55.5,-74,55.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-76.5,23,-74,23</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-76.5,7,-74,7</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-76.5,-9,-74,-9</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-76.5,-24,-74,-24</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-76.5,-39.5,-74,-39.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-45,-57.5,90.5</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 8</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 11</intersection>
<intersection>33.5 9</intersection>
<intersection>50 6</intersection>
<intersection>65.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-62.5,-45,-57.5,-45</points>
<connection>
<GID>762</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-62.5,50,-57.5,50</points>
<connection>
<GID>666</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-62.5,65.5,-57.5,65.5</points>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-62.5,-14.5,-57.5,-14.5</points>
<connection>
<GID>730</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-62.5,33.5,-57.5,33.5</points>
<connection>
<GID>682</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-62.5,1.5,-57.5,1.5</points>
<connection>
<GID>714</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-62.5,17.5,-57.5,17.5</points>
<connection>
<GID>698</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-62.5,-29.5,-57.5,-29.5</points>
<connection>
<GID>746</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-61.5,-55,71</points>
<connection>
<GID>799</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 3</intersection>
<intersection>7 4</intersection>
<intersection>23 5</intersection>
<intersection>39 6</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,71,-51.5,71</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,55.5,-51.5,55.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55,-9,-51.5,-9</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-55,7,-51.5,7</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-55,23,-51.5,23</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-55,39,-51.5,39</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-55,-24,-51.5,-24</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-55,-39.5,-51.5,-39.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-45,-36,90.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 9</intersection>
<intersection>33.5 8</intersection>
<intersection>50 7</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-41,-45,-36,-45</points>
<connection>
<GID>763</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-41,65.5,-36,65.5</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-41,50,-36,50</points>
<connection>
<GID>667</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-41,33.5,-36,33.5</points>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-41,17.5,-36,17.5</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-41,1.5,-36,1.5</points>
<connection>
<GID>715</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-41,-14.5,-36,-14.5</points>
<connection>
<GID>731</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-41,-29.5,-36,-29.5</points>
<connection>
<GID>747</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-61.5,-33.5,71</points>
<connection>
<GID>800</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 3</intersection>
<intersection>7 4</intersection>
<intersection>23 5</intersection>
<intersection>39 6</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,71,-30,71</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,55.5,-30,55.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-33.5,-9,-30,-9</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-33.5,7,-30,7</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-33.5,23,-30,23</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-33.5,39,-30,39</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-33.5,-24,-30,-24</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-33.5,-39.5,-30,-39.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-45,-14.5,90.5</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 10</intersection>
<intersection>-14.5 9</intersection>
<intersection>1.5 8</intersection>
<intersection>17.5 7</intersection>
<intersection>33.5 6</intersection>
<intersection>50 5</intersection>
<intersection>65.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-45,-14.5,-45</points>
<connection>
<GID>764</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-19.5,65.5,-14.5,65.5</points>
<connection>
<GID>652</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-19.5,50,-14.5,50</points>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-19.5,33.5,-14.5,33.5</points>
<connection>
<GID>684</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-19.5,17.5,-14.5,17.5</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-19.5,1.5,-14.5,1.5</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-19.5,-14.5,-14.5,-14.5</points>
<connection>
<GID>732</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-19.5,-29.5,-14.5,-29.5</points>
<connection>
<GID>748</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-61.5,-12,71</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-24 7</intersection>
<intersection>-9 6</intersection>
<intersection>7 5</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,71,-8.5,71</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12,55.5,-8.5,55.5</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12,39,-8.5,39</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-12,23,-8.5,23</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12,7,-8.5,7</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-12,-9,-8.5,-9</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-12,-24,-8.5,-24</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-12,-39.5,-8.5,-39.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-45,6,90.5</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>-45 5</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 9</intersection>
<intersection>33.5 8</intersection>
<intersection>50 7</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>2,-45,6,-45</points>
<connection>
<GID>765</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>2,65.5,6,65.5</points>
<connection>
<GID>653</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>2,50,6,50</points>
<connection>
<GID>669</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>2,33.5,6,33.5</points>
<connection>
<GID>685</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>2,17.5,6,17.5</points>
<connection>
<GID>701</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>2,1.5,6,1.5</points>
<connection>
<GID>717</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>2,-14.5,6,-14.5</points>
<connection>
<GID>733</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>2,-29.5,6,-29.5</points>
<connection>
<GID>749</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-61.5,8,71</points>
<connection>
<GID>802</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 7</intersection>
<intersection>-24 5</intersection>
<intersection>-9 6</intersection>
<intersection>7 8</intersection>
<intersection>23 4</intersection>
<intersection>39 3</intersection>
<intersection>55.5 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,71,11.5,71</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,55.5,11.5,55.5</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,39,11.5,39</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8,23,11.5,23</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>8,-24,11.5,-24</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>8,-9,11.5,-9</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>8,-39.5,11.5,-39.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>8,7,11.5,7</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-45,30.5,90.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-45 3</intersection>
<intersection>-29.5 12</intersection>
<intersection>-14.5 11</intersection>
<intersection>1.5 10</intersection>
<intersection>17.5 8</intersection>
<intersection>33.5 9</intersection>
<intersection>50 7</intersection>
<intersection>65.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22,-45,30.5,-45</points>
<connection>
<GID>766</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>22,65.5,30.5,65.5</points>
<connection>
<GID>654</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22,50,30.5,50</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>22,17.5,30.5,17.5</points>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22,33.5,30.5,33.5</points>
<connection>
<GID>686</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>22,1.5,30.5,1.5</points>
<connection>
<GID>718</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>22,-14.5,30.5,-14.5</points>
<connection>
<GID>734</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>22,-29.5,30.5,-29.5</points>
<connection>
<GID>750</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-16,102.5,-1</points>
<intersection>-16 4</intersection>
<intersection>-5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-5,107.5,-5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-1,102.5,-1</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102.5,-16,107.5,-16</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,60,19,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,71,19,71</points>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,60,22,60</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-22,108.5,-20</points>
<intersection>-22 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-20,120,-20</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-22,108.5,-22</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,44.5,18.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,55.5,18.5,55.5</points>
<connection>
<GID>662</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,44.5,22,44.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-18,116.5,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-15,116.5,-15</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-18,120,-18</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,60,-2,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,71,-2,71</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,60,2,60</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-14,105.5,-7</points>
<intersection>-14 2</intersection>
<intersection>-10.5 4</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-7,107.5,-7</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-14,107.5,-14</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>72,-10.5,105.5,-10.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,44.5,-2,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,55.5,-2,55.5</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,44.5,2,44.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,5,83,9.5</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>83,5,83.5,5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-4,18,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,7,18,7</points>
<connection>
<GID>710</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-4,22,-4</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,5.5,71.5,8.5</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>71.5,5.5,72,5.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,12,18.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,23,18.5,23</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,12,22,12</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-21,90.5,5</points>
<intersection>-21 3</intersection>
<intersection>0 1</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,0,91.5,0</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>90.5,-21,91.5,-21</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,5,90.5,5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,28,18.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,39,18.5,39</points>
<connection>
<GID>678</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,28,22,28</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-23,80.5,5.5</points>
<intersection>-23 4</intersection>
<intersection>-2 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,5.5,80.5,5.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-2,91.5,-2</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>80.5,-23,91.5,-23</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,28,-1.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,39,-1.5,39</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,28,2,28</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-6,118,-6</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,12,-1.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,23,-1.5,23</points>
<connection>
<GID>693</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,12,2,12</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,15.5,84,19</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-4,-2,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,7,-2,7</points>
<connection>
<GID>709</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-4,2,-4</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>72.5,15.5,82,15.5</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<intersection>72.5 5</intersection>
<intersection>76 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>72.5,14.5,72.5,15.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>76,15.5,76,27</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,60,-23,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,71,-23,71</points>
<connection>
<GID>643</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,60,-19.5,60</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-6,128.5,-6</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,44.5,-23,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,55.5,-23,55.5</points>
<connection>
<GID>660</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,44.5,-19.5,44.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,14.5,70.5,23.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,23.5,98.5,23.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection>
<intersection>84 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>84,23,84,23.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,28,-22.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,39,-22.5,39</points>
<connection>
<GID>676</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,28,-19.5,28</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,2.5,72,2.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<connection>
<GID>231</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,12,-22,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,23,-22,23</points>
<connection>
<GID>692</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22,12,-19.5,12</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,0,68,2</points>
<intersection>0 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,2,83.5,2</points>
<connection>
<GID>230</GID>
<name>clock</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,0,68,0</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-4,-23,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,7,-23,7</points>
<connection>
<GID>708</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-4,-19.5,-4</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-9,85.5,-5</points>
<intersection>-9 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-9,118,-9</points>
<connection>
<GID>232</GID>
<name>clock</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-5,85.5,-5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-4,-44,7</points>
<intersection>-4 2</intersection>
<intersection>7 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-44,-4,-41,-4</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-45.5,7,-44,7</points>
<connection>
<GID>707</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-16,191,-1</points>
<intersection>-16 4</intersection>
<intersection>-5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-5,196,-5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-1,191,-1</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>191,-16,196,-16</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,12,-44.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,23,-44.5,23</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,12,-41,12</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-22,197,-20</points>
<intersection>-22 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,-20,208.5,-20</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-22,197,-22</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,28,-44.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,39,-44.5,39</points>
<connection>
<GID>675</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,28,-41,28</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-18,205,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202,-15,205,-15</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>205,-18,208.5,-18</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,44.5,-44.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,55.5,-44.5,55.5</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,44.5,-41,44.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-14,194,-7</points>
<intersection>-14 2</intersection>
<intersection>-11.5 5</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,-7,196,-7</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194,-14,196,-14</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>126,-11.5,194,-11.5</points>
<intersection>126 6</intersection>
<intersection>194 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>126,-19,126,-11.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>-11.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,60,-44,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,71,-44,71</points>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44,60,-41,60</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,5,171.5,9.5</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>171.5,5,172,5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,60,-65.5,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,71,-65.5,71</points>
<connection>
<GID>641</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,60,-62.5,60</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,5.5,160,8.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>160,5.5,160.5,5.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,44.5,-66,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,55.5,-66,55.5</points>
<connection>
<GID>658</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,44.5,-62.5,44.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-21,179,5</points>
<intersection>-21 3</intersection>
<intersection>0 1</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179,0,180,0</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>179,-21,180,-21</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>178,5,179,5</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>179 0</intersection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,28,-66,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,39,-66,39</points>
<connection>
<GID>674</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,28,-62.5,28</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-23,169,5.5</points>
<intersection>-23 4</intersection>
<intersection>-2 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,5.5,169,5.5</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-2,180,-2</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>169,-23,180,-23</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,12,-66,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,23,-66,23</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,12,-62.5,12</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-6,206.5,-6</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,-4,-66,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,7,-66,7</points>
<connection>
<GID>706</GID>
<name>OUT_0</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,-4,-62.5,-4</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,15.5,172.5,19</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,-4,-86.5,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,7,-86.5,7</points>
<connection>
<GID>705</GID>
<name>OUT_0</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-4,-83,-4</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>-86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>161,15.5,170.5,15.5</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>161 5</intersection>
<intersection>164.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>161,14.5,161,15.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>164.5,15.5,164.5,27</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,12,-87,23</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87,12,-83,12</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,-6,217,-6</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,28,-86,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,39,-86,39</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,28,-83,28</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,14.5,159,23.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159,23.5,187,23.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection>
<intersection>172.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>172.5,23,172.5,23.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,44.5,-86.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,55.5,-86.5,55.5</points>
<connection>
<GID>657</GID>
<name>OUT_0</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,44.5,-83,44.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>-86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,2.5,160.5,2.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>249</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,60,-86,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,71,-86,71</points>
<connection>
<GID>640</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,60,-83,60</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,0,156.5,2</points>
<intersection>0 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,2,172,2</points>
<connection>
<GID>248</GID>
<name>clock</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141.5,0,156.5,0</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,60,-109.5,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,71,-109.5,71</points>
<connection>
<GID>639</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,60,-105.5,60</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-9,174,-5</points>
<intersection>-9 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,-9,206.5,-9</points>
<connection>
<GID>250</GID>
<name>clock</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141.5,-5,174,-5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,44.5,-109.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,55.5,-109.5,55.5</points>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,44.5,-105.5,44.5</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-16,281.5,-1</points>
<intersection>-16 4</intersection>
<intersection>-5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-5,286.5,-5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276.5,-1,281.5,-1</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>281.5,-16,286.5,-16</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,28,-109,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,39,-109,39</points>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109,28,-105.5,28</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-22,287.5,-20</points>
<intersection>-22 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-20,299,-20</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>287.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276.5,-22,287.5,-22</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>287.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,12,-109.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,23,-109.5,23</points>
<connection>
<GID>688</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,12,-105.5,12</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-18,295.5,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-15,295.5,-15</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,-18,299,-18</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-4,-109.5,7</points>
<intersection>-4 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,7,-109.5,7</points>
<connection>
<GID>704</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,-4,-105.5,-4</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-14,284.5,-7</points>
<intersection>-14 2</intersection>
<intersection>-12 3</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-7,286.5,-7</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>284.5,-14,286.5,-14</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>214.5,-12,284.5,-12</points>
<intersection>214.5 4</intersection>
<intersection>284.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>214.5,-19,214.5,-12</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-12 3</intersection></vsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,60,-132,71</points>
<intersection>60 2</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,71,-132,71</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132,60,-129,60</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,5,262,9.5</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>262,5,262.5,5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131.5,44.5,-131.5,55.5</points>
<intersection>44.5 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,55.5,-131.5,55.5</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>-131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-131.5,44.5,-129,44.5</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>-131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,5.5,250.5,8.5</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>250.5,5.5,251,5.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-133,-4,-133,7</points>
<connection>
<GID>703</GID>
<name>OUT_0</name></connection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-133,-4,-129,-4</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>-133 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-21,269.5,5</points>
<intersection>-21 3</intersection>
<intersection>0 1</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,0,270.5,0</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>269.5,-21,270.5,-21</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>268.5,5,269.5,5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,12,-132.5,23</points>
<intersection>12 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,23,-132.5,23</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,12,-129,12</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-23,259.5,5.5</points>
<intersection>-23 4</intersection>
<intersection>-2 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,5.5,259.5,5.5</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-2,270.5,-2</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>259.5,-23,270.5,-23</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>259.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,28,-132.5,39</points>
<intersection>28 2</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,39,-132.5,39</points>
<connection>
<GID>671</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,28,-129,28</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-6,297,-6</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<connection>
<GID>268</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,-20,-132,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-9,-132,-9</points>
<connection>
<GID>719</GID>
<name>OUT_0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132,-20,-129,-20</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,15.5,263,19</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-50.5,-109.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-39.5,-109.5,-39.5</points>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,-50.5,-105.5,-50.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>251.5,15.5,261,15.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>251.5 5</intersection>
<intersection>255 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>251.5,14.5,251.5,15.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>255,15.5,255,27</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-35,-110,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-24,-110,-24</points>
<connection>
<GID>736</GID>
<name>OUT_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-110,-35,-105.5,-35</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>303,-6,307.5,-6</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-20,-109.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-9,-109.5,-9</points>
<connection>
<GID>720</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-109.5,-20,-105.5,-20</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,14.5,249.5,23.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,23.5,277.5,23.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection>
<intersection>263 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>263,23,263,23.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,-20,-86,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,-9,-86,-9</points>
<connection>
<GID>721</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-20,-83,-20</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>232,2.5,251,2.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<connection>
<GID>267</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,0,247,2</points>
<intersection>0 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,2,262.5,2</points>
<connection>
<GID>266</GID>
<name>clock</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>232,0,247,0</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,-50.5,-86,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,-39.5,-86,-39.5</points>
<connection>
<GID>753</GID>
<name>OUT_0</name></connection>
<intersection>-86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-86,-50.5,-83,-50.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>-86 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-9,264.5,-5</points>
<intersection>-9 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-9,297,-9</points>
<connection>
<GID>268</GID>
<name>clock</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>232,-5,264.5,-5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,-35,-87,-24</points>
<connection>
<GID>737</GID>
<name>OUT_0</name></connection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87,-35,-83,-35</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-16,369,-1</points>
<intersection>-16 4</intersection>
<intersection>-5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369,-5,374,-5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>364,-1,369,-1</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>369,-16,374,-16</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-20,-66.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-9,-66.5,-9</points>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,-20,-62.5,-20</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375,-22,375,-20</points>
<intersection>-22 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375,-20,386.5,-20</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>375 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>364,-22,375,-22</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>375 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-50.5,-67,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-39.5,-67,-39.5</points>
<connection>
<GID>754</GID>
<name>OUT_0</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-67,-50.5,-62.5,-50.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383,-18,383,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-15,383,-15</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>383 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>383,-18,386.5,-18</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>383 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-35,-66.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-24,-66.5,-24</points>
<connection>
<GID>738</GID>
<name>OUT_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,-35,-62.5,-35</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-14,372,-7</points>
<intersection>-14 2</intersection>
<intersection>-12.5 3</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372,-7,374,-7</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,-14,374,-14</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>305,-12.5,372,-12.5</points>
<intersection>305 4</intersection>
<intersection>372 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>305,-19,305,-12.5</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>-12.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-35,-44.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-24,-44.5,-24</points>
<connection>
<GID>739</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-35,-41,-35</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,5,349.5,9.5</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>349.5,5,350,5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-50.5,-44.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-39.5,-44.5,-39.5</points>
<connection>
<GID>755</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-50.5,-41,-50.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338,5.5,338,8.5</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>338,5.5,338.5,5.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>338 0</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-20,-44.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-9,-44.5,-9</points>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-20,-41,-20</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-21,357,5</points>
<intersection>-21 3</intersection>
<intersection>0 1</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,0,358,0</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-21,358,-21</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>356,5,357,5</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-20,-23.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-9,-23.5,-9</points>
<connection>
<GID>724</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-20,-19.5,-20</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,-23,347,5.5</points>
<intersection>-23 4</intersection>
<intersection>-2 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,5.5,347,5.5</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>347 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347,-2,358,-2</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>347 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>347,-23,358,-23</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>347 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-35,-23,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-24,-23,-24</points>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-35,-19.5,-35</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>380,-6,384.5,-6</points>
<connection>
<GID>294</GID>
<name>OUT</name></connection>
<connection>
<GID>285</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-50.5,-23.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-39.5,-23.5,-39.5</points>
<connection>
<GID>756</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-50.5,-19.5,-50.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350.5,15.5,350.5,19</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-35,-1,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-24,-1,-24</points>
<connection>
<GID>741</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-35,2,-35</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>339,15.5,348.5,15.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>339 5</intersection>
<intersection>342.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>339,14.5,339,15.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>342.5,15.5,342.5,27</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-20,-1.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-9,-1.5,-9</points>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-20,2,-20</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>390.5,-6,395,-6</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-50.5,-1,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-39.5,-1,-39.5</points>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-50.5,2,-50.5</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,14.5,337,23.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>337,23.5,365,23.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>337 0</intersection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,23,350.5,23.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-20,18.5,-9</points>
<intersection>-20 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-9,18.5,-9</points>
<connection>
<GID>726</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-20,22,-20</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>319.5,2.5,338.5,2.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<connection>
<GID>284</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-35,18.5,-24</points>
<intersection>-35 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-24,18.5,-24</points>
<connection>
<GID>742</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-35,22,-35</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,0,334.5,2</points>
<intersection>0 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334.5,2,350,2</points>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<intersection>334.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>319.5,0,334.5,0</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>334.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-50.5,18.5,-39.5</points>
<intersection>-50.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-39.5,18.5,-39.5</points>
<connection>
<GID>758</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-50.5,22,-50.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-9,352,-5</points>
<intersection>-9 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-9,384.5,-9</points>
<connection>
<GID>285</GID>
<name>clock</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>319.5,-5,352,-5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-368,29,-365,29</points>
<connection>
<GID>846</GID>
<name>OUT_0</name></connection>
<connection>
<GID>869</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-16,456,-1</points>
<intersection>-16 4</intersection>
<intersection>-5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456,-5,461,-5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451,-1,456,-1</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>456,-16,461,-16</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>456 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-368,21.5,-364,21.5</points>
<connection>
<GID>847</GID>
<name>OUT_0</name></connection>
<connection>
<GID>871</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462,-22,462,-20</points>
<intersection>-22 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>462,-20,473.5,-20</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451,-22,462,-22</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>462 0</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-368,14.5,-364,14.5</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<connection>
<GID>848</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-18,470,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-15,470,-15</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<intersection>470 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>470,-18,473.5,-18</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>470 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-352,-1.5,-352,4</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<connection>
<GID>849</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-14,459,-7</points>
<intersection>-14 2</intersection>
<intersection>-12 3</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459,-7,461,-7</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>459 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>459,-14,461,-14</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>459 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>392.5,-12,459,-12</points>
<intersection>392.5 4</intersection>
<intersection>459 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>392.5,-19,392.5,-12</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>-12 3</intersection></vsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-344,-1.5,-344,4</points>
<connection>
<GID>874</GID>
<name>IN_0</name></connection>
<connection>
<GID>850</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,5,436.5,9.5</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>436.5,5,437,5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-337,-1,-337,4</points>
<connection>
<GID>851</GID>
<name>OUT_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425,5.5,425,8.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>425,5.5,425.5,5.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>425 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-331,-0.5,-331,4</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<connection>
<GID>852</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,-21,444,5</points>
<intersection>-21 3</intersection>
<intersection>0 1</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444,0,445,0</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>444,-21,445,-21</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>443,5,444,5</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-325,-1.5,-325,4.5</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<connection>
<GID>853</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434,-23,434,5.5</points>
<intersection>-23 4</intersection>
<intersection>-2 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,5.5,434,5.5</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>434,-2,445,-2</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>434,-23,445,-23</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>434 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-319,-1.5,-319,4</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<connection>
<GID>854</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>467,-6,471.5,-6</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<connection>
<GID>302</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-313,-1,-313,4</points>
<connection>
<GID>855</GID>
<name>OUT_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437.5,15.5,437.5,19</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-306,-1,-306,4</points>
<connection>
<GID>856</GID>
<name>OUT_0</name></connection>
<connection>
<GID>880</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>426,15.5,435.5,15.5</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>426 5</intersection>
<intersection>429.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>426,14.5,426,15.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>429.5,15.5,429.5,27</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-355,44,-355,52</points>
<connection>
<GID>858</GID>
<name>N_in3</name></connection>
<connection>
<GID>882</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-6,482,-6</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<connection>
<GID>304</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-346.5,44,-346.5,51.5</points>
<connection>
<GID>861</GID>
<name>N_in3</name></connection>
<connection>
<GID>883</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424,14.5,424,23.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424,23.5,452,23.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>424 0</intersection>
<intersection>437.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>437.5,23,437.5,23.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-339,44,-339,51.5</points>
<connection>
<GID>862</GID>
<name>N_in3</name></connection>
<connection>
<GID>884</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406.5,2.5,425.5,2.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<connection>
<GID>301</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-333,44,-333,52</points>
<connection>
<GID>863</GID>
<name>N_in3</name></connection>
<connection>
<GID>885</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,0,421.5,2</points>
<intersection>0 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>421.5,2,437,2</points>
<connection>
<GID>300</GID>
<name>clock</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>406.5,0,421.5,0</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-326.5,44,-326.5,52</points>
<connection>
<GID>864</GID>
<name>N_in3</name></connection>
<connection>
<GID>886</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>439,-9,439,-5</points>
<intersection>-9 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>439,-9,471.5,-9</points>
<connection>
<GID>302</GID>
<name>clock</name></connection>
<intersection>439 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>406.5,-5,439,-5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>439 0</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-320.5,44,-320.5,52</points>
<connection>
<GID>865</GID>
<name>N_in3</name></connection>
<connection>
<GID>887</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542,-16.5,542,-1.5</points>
<intersection>-16.5 4</intersection>
<intersection>-5.5 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>542,-5.5,547,-5.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>537,-1.5,542,-1.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>542,-16.5,547,-16.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>542 0</intersection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-313.5,44,-313.5,52</points>
<connection>
<GID>866</GID>
<name>N_in3</name></connection>
<connection>
<GID>888</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>548,-22.5,548,-20.5</points>
<intersection>-22.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>548,-20.5,559.5,-20.5</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>548 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>537,-22.5,548,-22.5</points>
<connection>
<GID>330</GID>
<name>OUT</name></connection>
<intersection>548 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-308,44,-308,52</points>
<connection>
<GID>867</GID>
<name>N_in3</name></connection>
<connection>
<GID>889</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>556,-18.5,556,-15.5</points>
<intersection>-18.5 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>553,-15.5,556,-15.5</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>556 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>556,-18.5,559.5,-18.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>556 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-270,23.5,-246.5,23.5</points>
<connection>
<GID>786</GID>
<name>ENABLE</name></connection>
<connection>
<GID>794</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>545,-14.5,545,-7.5</points>
<intersection>-14.5 2</intersection>
<intersection>-12.5 3</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>545,-7.5,547,-7.5</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>545 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>545,-14.5,547,-14.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>545 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>479.5,-12.5,545,-12.5</points>
<intersection>479.5 4</intersection>
<intersection>545 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>479.5,-19,479.5,-12.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>-12.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-261.5,19,-246.5,19</points>
<connection>
<GID>788</GID>
<name>OUT_0</name></connection>
<intersection>-246.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-246.5,18.5,-246.5,19</points>
<connection>
<GID>786</GID>
<name>IN_2</name></connection>
<intersection>19 1</intersection></vsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>522.5,4.5,522.5,9</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>4.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>522.5,4.5,523,4.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>522.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,5,511,8</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<intersection>5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>511,5,511.5,5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-254,14.5,-254,17.5</points>
<intersection>14.5 2</intersection>
<intersection>17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-254,17.5,-246.5,17.5</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>-254 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261.5,14.5,-254,14.5</points>
<connection>
<GID>790</GID>
<name>OUT_0</name></connection>
<intersection>-254 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,-21.5,530,4.5</points>
<intersection>-21.5 3</intersection>
<intersection>-0.5 1</intersection>
<intersection>4.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-0.5,531,-0.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>530,-21.5,531,-21.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>529,4.5,530,4.5</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<intersection>530 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-252.5,11.5,-252.5,16.5</points>
<intersection>11.5 2</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-252.5,16.5,-246.5,16.5</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>-252.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-261.5,11.5,-252.5,11.5</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<intersection>-252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520,-23.5,520,5</points>
<intersection>-23.5 4</intersection>
<intersection>-2.5 2</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517.5,5,520,5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>520 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520,-2.5,531,-2.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>520 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>520,-23.5,531,-23.5</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<intersection>520 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>553,-6.5,557.5,-6.5</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<connection>
<GID>319</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>523.5,15,523.5,18.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>512,15,521.5,15</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>512 5</intersection>
<intersection>515.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>512,14,512,15</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>515.5,15,515.5,26.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>563.5,-6.5,568,-6.5</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<connection>
<GID>321</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,14,510,23</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,23,538,23</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection>
<intersection>523.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>523.5,22.5,523.5,23</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>23 1</intersection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>492.5,2,511.5,2</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507.5,-0.5,507.5,1.5</points>
<intersection>-0.5 2</intersection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507.5,1.5,523,1.5</points>
<connection>
<GID>317</GID>
<name>clock</name></connection>
<intersection>507.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,-0.5,507.5,-0.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>507.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525,-9.5,525,-5.5</points>
<intersection>-9.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,-9.5,557.5,-9.5</points>
<connection>
<GID>319</GID>
<name>clock</name></connection>
<intersection>525 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,-5.5,525,-5.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>525 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>632.5,-15.5,632.5,-0.5</points>
<intersection>-15.5 4</intersection>
<intersection>-4.5 1</intersection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>632.5,-4.5,637.5,-4.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>632.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>627.5,-0.5,632.5,-0.5</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>632.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>632.5,-15.5,637.5,-15.5</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>632.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638.5,-21.5,638.5,-19.5</points>
<intersection>-21.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>638.5,-19.5,650,-19.5</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>638.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>627.5,-21.5,638.5,-21.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>638.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>646.5,-17.5,646.5,-14.5</points>
<intersection>-17.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643.5,-14.5,646.5,-14.5</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>646.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>646.5,-17.5,650,-17.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>646.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>635.5,-13.5,635.5,-6.5</points>
<intersection>-13.5 2</intersection>
<intersection>-12 3</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>635.5,-6.5,637.5,-6.5</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>635.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>635.5,-13.5,637.5,-13.5</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>635.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>565.5,-12,635.5,-12</points>
<intersection>565.5 4</intersection>
<intersection>635.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>565.5,-19.5,565.5,-12</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>-12 3</intersection></vsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>613,5.5,613,10</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>5.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>613,5.5,613.5,5.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>613 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>601.5,6,601.5,9</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>601.5,6,602,6</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>601.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>620.5,-20.5,620.5,5.5</points>
<intersection>-20.5 3</intersection>
<intersection>0.5 1</intersection>
<intersection>5.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>620.5,0.5,621.5,0.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>620.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>620.5,-20.5,621.5,-20.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>620.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>619.5,5.5,620.5,5.5</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>620.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>610.5,-22.5,610.5,6</points>
<intersection>-22.5 4</intersection>
<intersection>-1.5 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>608,6,610.5,6</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<intersection>610.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>610.5,-1.5,621.5,-1.5</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<intersection>610.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>610.5,-22.5,621.5,-22.5</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>610.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>643.5,-5.5,648,-5.5</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<connection>
<GID>353</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>614,16,614,19.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>602.5,16,612,16</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>602.5 5</intersection>
<intersection>606 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>602.5,15,602.5,16</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>606,16,606,27.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></vsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>654,-5.5,658.5,-5.5</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<connection>
<GID>355</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600.5,15,600.5,24</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>600.5,24,628.5,24</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>600.5 0</intersection>
<intersection>614 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>614,23.5,614,24</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583,3,602,3</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<connection>
<GID>352</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>598,0.5,598,2.5</points>
<intersection>0.5 2</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>598,2.5,613.5,2.5</points>
<connection>
<GID>351</GID>
<name>clock</name></connection>
<intersection>598 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583,0.5,598,0.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>598 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>615.5,-8.5,615.5,-4.5</points>
<intersection>-8.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>615.5,-8.5,648,-8.5</points>
<connection>
<GID>353</GID>
<name>clock</name></connection>
<intersection>615.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583,-4.5,615.5,-4.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>615.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>720,-14,720,1</points>
<intersection>-14 4</intersection>
<intersection>-3 1</intersection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>720,-3,725,-3</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>720 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>715,1,720,1</points>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<intersection>720 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>720,-14,725,-14</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>720 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>726,-20,726,-18</points>
<intersection>-20 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>726,-18,737.5,-18</points>
<connection>
<GID>399</GID>
<name>IN_1</name></connection>
<intersection>726 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>715,-20,726,-20</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<intersection>726 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>734,-16,734,-13</points>
<intersection>-16 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>731,-13,734,-13</points>
<connection>
<GID>397</GID>
<name>OUT</name></connection>
<intersection>734 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>734,-16,737.5,-16</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>734 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>723,-12,723,-5</points>
<intersection>-12 2</intersection>
<intersection>-11 3</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>723,-5,725,-5</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>723 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>723,-12,725,-12</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>723 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>656,-11,723,-11</points>
<intersection>656 4</intersection>
<intersection>723 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>656,-18.5,656,-11</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>-11 3</intersection></vsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>700.5,7,700.5,11.5</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>7 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>700.5,7,701,7</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>700.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,7.5,689,10.5</points>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>689,7.5,689.5,7.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>689 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>708,-19,708,7</points>
<intersection>-19 3</intersection>
<intersection>2 1</intersection>
<intersection>7 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>708,2,709,2</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<intersection>708 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>708,-19,709,-19</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>708 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>707,7,708,7</points>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<intersection>708 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698,-21,698,7.5</points>
<intersection>-21 4</intersection>
<intersection>0 2</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>695.5,7.5,698,7.5</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<intersection>698 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>698,0,709,0</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<intersection>698 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>698,-21,709,-21</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<intersection>698 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>731,-4,735.5,-4</points>
<connection>
<GID>396</GID>
<name>OUT</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>701.5,17.5,701.5,21</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<connection>
<GID>400</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>690,17.5,699.5,17.5</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>690 5</intersection>
<intersection>693.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>690,16.5,690,17.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>17.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>693.5,17.5,693.5,29</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>17.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>741.5,-4,746,-4</points>
<connection>
<GID>387</GID>
<name>OUT_0</name></connection>
<connection>
<GID>389</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>688,16.5,688,25.5</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<intersection>25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>688,25.5,716,25.5</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>688 0</intersection>
<intersection>701.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>701.5,25,701.5,25.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>670.5,4.5,689.5,4.5</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<connection>
<GID>386</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>685.5,2,685.5,4</points>
<intersection>2 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>685.5,4,701,4</points>
<connection>
<GID>385</GID>
<name>clock</name></connection>
<intersection>685.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>670.5,2,685.5,2</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>685.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>703,-7,703,-3</points>
<intersection>-7 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>703,-7,735.5,-7</points>
<connection>
<GID>387</GID>
<name>clock</name></connection>
<intersection>703 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>670.5,-3,703,-3</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>703 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>743.5,-17,751,-17</points>
<connection>
<GID>399</GID>
<name>OUT</name></connection>
<connection>
<GID>403</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-266,36.5,-256.5,36.5</points>
<connection>
<GID>408</GID>
<name>N_in0</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,33,-295.5,33</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<connection>
<GID>412</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,21.5,-295,21.5</points>
<connection>
<GID>406</GID>
<name>OUT_0</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,25.5,-295,25.5</points>
<connection>
<GID>405</GID>
<name>OUT_0</name></connection>
<connection>
<GID>414</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,29,-295,29</points>
<connection>
<GID>404</GID>
<name>OUT_0</name></connection>
<connection>
<GID>413</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>684.485,106.519,1317.1,-206.171</PageViewport>
<gate>
<ID>197</ID>
<type>AE_DFF_LOW</type>
<position>783.5,-11</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>131 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_DFF_LOW</type>
<position>772,-10.5</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>132 </output>
<input>
<ID>clock</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_DFF_LOW</type>
<position>818,-22</position>
<input>
<ID>IN_0</ID>138 </input>
<output>
<ID>OUT_0</ID>146 </output>
<input>
<ID>clock</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>214</ID>
<type>AE_SMALL_INVERTER</type>
<position>781,7</position>
<input>
<ID>IN_0</ID>147 </input>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>DE_TO</type>
<position>827.5,-20</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L1</lparam></gate>
<gate>
<ID>220</ID>
<type>DA_FROM</type>
<position>773,15</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>748,-11.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>748,-14</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>797.5,9.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>748,-19</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP</lparam></gate>
<gate>
<ID>507</ID>
<type>AE_DFF_LOW</type>
<position>482,1.5</position>
<input>
<ID>IN_0</ID>389 </input>
<output>
<ID>OUT_0</ID>398 </output>
<input>
<ID>clock</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>509</ID>
<type>AE_DFF_LOW</type>
<position>516.5,2</position>
<input>
<ID>IN_0</ID>390 </input>
<output>
<ID>OUT_0</ID>399 </output>
<input>
<ID>clock</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>511</ID>
<type>AE_DFF_LOW</type>
<position>546.5,2</position>
<input>
<ID>IN_0</ID>391 </input>
<output>
<ID>OUT_0</ID>400 </output>
<input>
<ID>clock</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>898</ID>
<type>GA_LED</type>
<position>506.5,57</position>
<input>
<ID>N_in2</ID>647 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>513</ID>
<type>AE_DFF_LOW</type>
<position>578,2.5</position>
<input>
<ID>IN_0</ID>392 </input>
<output>
<ID>OUT_0</ID>401 </output>
<input>
<ID>clock</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>899</ID>
<type>GA_LED</type>
<position>539,57</position>
<input>
<ID>N_in2</ID>648 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>900</ID>
<type>GA_LED</type>
<position>569.5,57</position>
<input>
<ID>N_in2</ID>649 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>AE_DFF_LOW</type>
<position>481.5,-22</position>
<input>
<ID>IN_0</ID>389 </input>
<output>
<ID>OUT_0</ID>402 </output>
<input>
<ID>clock</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>901</ID>
<type>GA_LED</type>
<position>601,57</position>
<input>
<ID>N_in2</ID>650 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>AE_DFF_LOW</type>
<position>515.5,-21.5</position>
<input>
<ID>IN_0</ID>390 </input>
<output>
<ID>OUT_0</ID>403 </output>
<input>
<ID>clock</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>519</ID>
<type>AE_DFF_LOW</type>
<position>546,-21.5</position>
<input>
<ID>IN_0</ID>391 </input>
<output>
<ID>OUT_0</ID>404 </output>
<input>
<ID>clock</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>521</ID>
<type>AE_DFF_LOW</type>
<position>578,-22</position>
<input>
<ID>IN_0</ID>392 </input>
<output>
<ID>OUT_0</ID>405 </output>
<input>
<ID>clock</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>523</ID>
<type>AA_AND2</type>
<position>452,2.5</position>
<input>
<ID>IN_0</ID>365 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>369 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>525</ID>
<type>AA_AND2</type>
<position>458.5,-3.5</position>
<input>
<ID>IN_0</ID>365 </input>
<input>
<ID>IN_1</ID>652 </input>
<output>
<ID>OUT</ID>406 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND2</type>
<position>451.5,-16.5</position>
<input>
<ID>IN_0</ID>366 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>529</ID>
<type>AA_AND2</type>
<position>460,-24</position>
<input>
<ID>IN_0</ID>366 </input>
<input>
<ID>IN_1</ID>652 </input>
<output>
<ID>OUT</ID>407 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>924</ID>
<type>AA_TOGGLE</type>
<position>462,22</position>
<output>
<ID>OUT_0</ID>651 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>926</ID>
<type>AA_TOGGLE</type>
<position>452,19</position>
<output>
<ID>OUT_0</ID>652 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>542</ID>
<type>BA_TRI_STATE</type>
<position>494.5,-8.5</position>
<input>
<ID>ENABLE_0</ID>406 </input>
<input>
<ID>IN_0</ID>398 </input>
<output>
<ID>OUT_0</ID>393 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>543</ID>
<type>BA_TRI_STATE</type>
<position>499.5,-33</position>
<input>
<ID>ENABLE_0</ID>407 </input>
<input>
<ID>IN_0</ID>402 </input>
<output>
<ID>OUT_0</ID>393 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>544</ID>
<type>BA_TRI_STATE</type>
<position>536,-8</position>
<input>
<ID>ENABLE_0</ID>406 </input>
<input>
<ID>IN_0</ID>399 </input>
<output>
<ID>OUT_0</ID>394 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>545</ID>
<type>BA_TRI_STATE</type>
<position>534.5,-34</position>
<input>
<ID>ENABLE_0</ID>407 </input>
<input>
<ID>IN_0</ID>403 </input>
<output>
<ID>OUT_0</ID>394 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>546</ID>
<type>BA_TRI_STATE</type>
<position>566.5,-8</position>
<input>
<ID>ENABLE_0</ID>406 </input>
<input>
<ID>IN_0</ID>400 </input>
<output>
<ID>OUT_0</ID>396 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>547</ID>
<type>BA_TRI_STATE</type>
<position>566,-34.5</position>
<input>
<ID>ENABLE_0</ID>407 </input>
<input>
<ID>IN_0</ID>404 </input>
<output>
<ID>OUT_0</ID>396 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>548</ID>
<type>BA_TRI_STATE</type>
<position>598,-7.5</position>
<input>
<ID>ENABLE_0</ID>406 </input>
<input>
<ID>IN_0</ID>401 </input>
<output>
<ID>OUT_0</ID>397 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>549</ID>
<type>BA_TRI_STATE</type>
<position>598,-33</position>
<input>
<ID>ENABLE_0</ID>407 </input>
<input>
<ID>IN_0</ID>405 </input>
<output>
<ID>OUT_0</ID>397 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>551</ID>
<type>BA_TRI_STATE</type>
<position>507,22</position>
<input>
<ID>ENABLE_0</ID>651 </input>
<input>
<ID>IN_0</ID>393 </input>
<output>
<ID>OUT_0</ID>647 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>552</ID>
<type>BA_TRI_STATE</type>
<position>539,22</position>
<input>
<ID>ENABLE_0</ID>651 </input>
<input>
<ID>IN_0</ID>394 </input>
<output>
<ID>OUT_0</ID>648 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AI_XOR2</type>
<position>791.5,-15</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>553</ID>
<type>BA_TRI_STATE</type>
<position>570,22</position>
<input>
<ID>ENABLE_0</ID>651 </input>
<input>
<ID>IN_0</ID>396 </input>
<output>
<ID>OUT_0</ID>649 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>168</ID>
<type>AI_XOR2</type>
<position>807.5,-20</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>554</ID>
<type>BA_TRI_STATE</type>
<position>601.5,22</position>
<input>
<ID>ENABLE_0</ID>651 </input>
<input>
<ID>IN_0</ID>397 </input>
<output>
<ID>OUT_0</ID>650 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND2</type>
<position>807.5,-29</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>BA_TRI_STATE</type>
<position>476.5,-46.5</position>
<input>
<ID>ENABLE_0</ID>388 </input>
<input>
<ID>IN_0</ID>356 </input>
<output>
<ID>OUT_0</ID>389 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>791.5,-36</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>BA_TRI_STATE</type>
<position>507,-46</position>
<input>
<ID>ENABLE_0</ID>388 </input>
<input>
<ID>IN_0</ID>357 </input>
<output>
<ID>OUT_0</ID>390 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>171</ID>
<type>AE_OR2</type>
<position>820,-33</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>557</ID>
<type>BA_TRI_STATE</type>
<position>540.5,-46.5</position>
<input>
<ID>ENABLE_0</ID>388 </input>
<input>
<ID>IN_0</ID>358 </input>
<output>
<ID>OUT_0</ID>391 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>558</ID>
<type>BA_TRI_STATE</type>
<position>571,-45.5</position>
<input>
<ID>ENABLE_0</ID>388 </input>
<input>
<ID>IN_0</ID>359 </input>
<output>
<ID>OUT_0</ID>392 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_TOGGLE</type>
<position>767,-24.5</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>560</ID>
<type>AA_INVERTER</type>
<position>434.5,-7</position>
<input>
<ID>IN_0</ID>365 </input>
<output>
<ID>OUT_0</ID>366 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>562</ID>
<type>AA_TOGGLE</type>
<position>425.5,0.5</position>
<output>
<ID>OUT_0</ID>365 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>566</ID>
<type>AA_TOGGLE</type>
<position>441,-42.5</position>
<output>
<ID>OUT_0</ID>367 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>780,-1.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_TOGGLE</type>
<position>460.5,-46.5</position>
<output>
<ID>OUT_0</ID>388 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND2</type>
<position>768.5,-2.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>570</ID>
<type>AA_TOGGLE</type>
<position>475.5,-60</position>
<output>
<ID>OUT_0</ID>356 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>571</ID>
<type>AA_TOGGLE</type>
<position>507,-59.5</position>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_TOGGLE</type>
<position>538.5,-58.5</position>
<output>
<ID>OUT_0</ID>358 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>573</ID>
<type>AA_TOGGLE</type>
<position>571,-58</position>
<output>
<ID>OUT_0</ID>359 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462.5,-46.5,569,-46.5</points>
<connection>
<GID>557</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>555</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>568</GID>
<name>OUT_0</name></connection>
<intersection>505 3</intersection>
<intersection>569 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>505,-46.5,505,-46</points>
<connection>
<GID>556</GID>
<name>ENABLE_0</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>569,-46.5,569,-45.5</points>
<connection>
<GID>558</GID>
<name>ENABLE_0</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>476.5,-44,476.5,3.5</points>
<connection>
<GID>555</GID>
<name>OUT_0</name></connection>
<intersection>-20 2</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>476.5,3.5,479,3.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>476.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>476.5,-20,478.5,-20</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>476.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,-43.5,507,4</points>
<connection>
<GID>556</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507,4,513.5,4</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507,-19.5,512.5,-19.5</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>507 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-44,540.5,4</points>
<connection>
<GID>557</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540.5,4,543.5,4</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-19.5,543,-19.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571,-43,571,4.5</points>
<connection>
<GID>558</GID>
<name>OUT_0</name></connection>
<intersection>-20 2</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571,4.5,575,4.5</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>571 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>571,-20,575,-20</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>571 0</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503.5,-30.5,503.5,19</points>
<intersection>-30.5 4</intersection>
<intersection>-5.5 5</intersection>
<intersection>19 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>503.5,19,507,19</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>503.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>499.5,-30.5,503.5,-30.5</points>
<connection>
<GID>543</GID>
<name>OUT_0</name></connection>
<intersection>503.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>494.5,-5.5,503.5,-5.5</points>
<intersection>494.5 6</intersection>
<intersection>503.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>494.5,-6,494.5,-5.5</points>
<connection>
<GID>542</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,-31.5,539,19</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>-31.5 3</intersection>
<intersection>-5.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>534.5,-31.5,539,-31.5</points>
<connection>
<GID>545</GID>
<name>OUT_0</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>536,-5.5,539,-5.5</points>
<connection>
<GID>544</GID>
<name>OUT_0</name></connection>
<intersection>539 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570,-32,570,19</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>-32 3</intersection>
<intersection>-5.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>566,-32,570,-32</points>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection>
<intersection>570 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>566.5,-5.5,570,-5.5</points>
<connection>
<GID>546</GID>
<name>OUT_0</name></connection>
<intersection>570 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>601.5,-5.5,601.5,19</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-5.5 2</intersection>
<intersection>-5 4</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>602,-30.5,602,-5.5</points>
<intersection>-30.5 3</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>601.5,-5.5,602,-5.5</points>
<intersection>601.5 0</intersection>
<intersection>602 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>598,-30.5,602,-30.5</points>
<connection>
<GID>549</GID>
<name>OUT_0</name></connection>
<intersection>602 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>598,-5,601.5,-5</points>
<connection>
<GID>548</GID>
<name>OUT_0</name></connection>
<intersection>601.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490,-11.5,490,3.5</points>
<intersection>-11.5 2</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>485,3.5,490,3.5</points>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>490,-11.5,494.5,-11.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>529.5,-11,529.5,4</points>
<intersection>-11 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>519.5,4,529.5,4</points>
<connection>
<GID>509</GID>
<name>OUT_0</name></connection>
<intersection>529.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529.5,-11,536,-11</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>529.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>560.5,-11,560.5,4</points>
<intersection>-11 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>549.5,4,560.5,4</points>
<connection>
<GID>511</GID>
<name>OUT_0</name></connection>
<intersection>560.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>560.5,-11,566.5,-11</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>560.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-10.5,589.5,4.5</points>
<intersection>-10.5 2</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581,4.5,589.5,4.5</points>
<connection>
<GID>513</GID>
<name>OUT_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,-10.5,598,-10.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,-36,492.5,-20</points>
<intersection>-36 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484.5,-20,492.5,-20</points>
<connection>
<GID>515</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,-36,499.5,-36</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,-37,524.5,-19.5</points>
<intersection>-37 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>518.5,-19.5,524.5,-19.5</points>
<connection>
<GID>517</GID>
<name>OUT_0</name></connection>
<intersection>524.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>524.5,-37,534.5,-37</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>524.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>554.5,-37.5,554.5,-19.5</points>
<intersection>-37.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>549,-19.5,554.5,-19.5</points>
<connection>
<GID>519</GID>
<name>OUT_0</name></connection>
<intersection>554.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>554.5,-37.5,566,-37.5</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>554.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-36,589.5,-20</points>
<intersection>-36 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581,-20,589.5,-20</points>
<connection>
<GID>521</GID>
<name>OUT_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,-36,598,-36</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477,-8.5,477,-3.5</points>
<intersection>-8.5 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-8.5,534,-8.5</points>
<connection>
<GID>542</GID>
<name>ENABLE_0</name></connection>
<intersection>477 0</intersection>
<intersection>534 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>461.5,-3.5,477,-3.5</points>
<connection>
<GID>525</GID>
<name>OUT</name></connection>
<intersection>477 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>534,-8.5,534,-8</points>
<connection>
<GID>544</GID>
<name>ENABLE_0</name></connection>
<intersection>-8.5 1</intersection>
<intersection>-8 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>534,-8,596,-8</points>
<connection>
<GID>546</GID>
<name>ENABLE_0</name></connection>
<intersection>534 3</intersection>
<intersection>596 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>596,-8,596,-7.5</points>
<connection>
<GID>548</GID>
<name>ENABLE_0</name></connection>
<intersection>-8 4</intersection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>480,-33,480,-24</points>
<intersection>-33 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-33,532.5,-33</points>
<connection>
<GID>543</GID>
<name>ENABLE_0</name></connection>
<intersection>480 0</intersection>
<intersection>532.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>463,-24,480,-24</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<intersection>480 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>532.5,-34.5,532.5,-33</points>
<connection>
<GID>545</GID>
<name>ENABLE_0</name></connection>
<intersection>-34.5 4</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>532.5,-34.5,596,-34.5</points>
<connection>
<GID>547</GID>
<name>ENABLE_0</name></connection>
<intersection>532.5 3</intersection>
<intersection>596 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>596,-34.5,596,-33</points>
<connection>
<GID>549</GID>
<name>ENABLE_0</name></connection>
<intersection>-34.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506.5,40,506.5,56</points>
<connection>
<GID>898</GID>
<name>N_in2</name></connection>
<intersection>40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>507,24.5,507,40</points>
<connection>
<GID>551</GID>
<name>OUT_0</name></connection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>506.5,40,507,40</points>
<intersection>506.5 0</intersection>
<intersection>507 1</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,24.5,539,56</points>
<connection>
<GID>899</GID>
<name>N_in2</name></connection>
<connection>
<GID>552</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,40,569.5,56</points>
<connection>
<GID>900</GID>
<name>N_in2</name></connection>
<intersection>40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>570,24.5,570,40</points>
<connection>
<GID>553</GID>
<name>OUT_0</name></connection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>569.5,40,570,40</points>
<intersection>569.5 0</intersection>
<intersection>570 1</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>601,40,601,56</points>
<connection>
<GID>901</GID>
<name>N_in2</name></connection>
<intersection>40 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>601.5,24.5,601.5,40</points>
<connection>
<GID>554</GID>
<name>OUT_0</name></connection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>601,40,601.5,40</points>
<intersection>601 0</intersection>
<intersection>601.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>464,22,599.5,22</points>
<connection>
<GID>554</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>553</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>552</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>551</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>924</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-25,456,19</points>
<intersection>-25 3</intersection>
<intersection>-4.5 1</intersection>
<intersection>19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455.5,-4.5,456,-4.5</points>
<connection>
<GID>525</GID>
<name>IN_1</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>454,19,456,19</points>
<connection>
<GID>926</GID>
<name>OUT_0</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>456,-25,457,-25</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>456 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>799.5,-30,799.5,-15</points>
<intersection>-30 4</intersection>
<intersection>-19 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>799.5,-19,804.5,-19</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>799.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>794.5,-15,799.5,-15</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>799.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>799.5,-30,804.5,-30</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>799.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>805.5,-36,805.5,-34</points>
<intersection>-36 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>805.5,-34,817,-34</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>805.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>794.5,-36,805.5,-36</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>805.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>813.5,-32,813.5,-29</points>
<intersection>-32 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>810.5,-29,813.5,-29</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>813.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>813.5,-32,817,-32</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>813.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>802.5,-28,802.5,-21</points>
<intersection>-28 2</intersection>
<intersection>-24.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>802.5,-21,804.5,-21</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>802.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>802.5,-28,804.5,-28</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>802.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>769,-24.5,802.5,-24.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>802.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>780,-9,780,-4.5</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>-9 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>780,-9,780.5,-9</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>780 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>768.5,-8.5,768.5,-5.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>768.5,-8.5,769,-8.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>768.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>787.5,-35,787.5,-9</points>
<intersection>-35 3</intersection>
<intersection>-14 1</intersection>
<intersection>-9 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>787.5,-14,788.5,-14</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>787.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>787.5,-35,788.5,-35</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>787.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>786.5,-9,787.5,-9</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>787.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>777.5,-37,777.5,-8.5</points>
<intersection>-37 4</intersection>
<intersection>-16 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>775,-8.5,777.5,-8.5</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>777.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>777.5,-16,788.5,-16</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>777.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>777.5,-37,788.5,-37</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>777.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>810.5,-20,815,-20</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>781,1.5,781,5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>769.5,1.5,779,1.5</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>769.5 5</intersection>
<intersection>773 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>769.5,0.5,769.5,1.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>1.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>773,1.5,773,13</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>1.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>821,-20,825.5,-20</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<connection>
<GID>218</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>767.5,0.5,767.5,9.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>767.5,9.5,795.5,9.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>767.5 0</intersection>
<intersection>781 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>781,9,781,9.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>750,-11.5,769,-11.5</points>
<connection>
<GID>199</GID>
<name>clock</name></connection>
<connection>
<GID>222</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>765,-14,765,-12</points>
<intersection>-14 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>765,-12,780.5,-12</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>765 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>750,-14,765,-14</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>765 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>782.5,-23,782.5,-19</points>
<intersection>-23 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>782.5,-23,815,-23</points>
<connection>
<GID>206</GID>
<name>clock</name></connection>
<intersection>782.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>750,-19,782.5,-19</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>782.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>476.5,-53.5,476.5,-49.5</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>475.5,-58,475.5,-53.5</points>
<connection>
<GID>570</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>475.5,-53.5,476.5,-53.5</points>
<intersection>475.5 1</intersection>
<intersection>476.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,-57.5,507,-49</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<connection>
<GID>571</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-56.5,540.5,-49.5</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>-56.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>538.5,-56.5,540.5,-56.5</points>
<connection>
<GID>572</GID>
<name>OUT_0</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571,-56,571,-48.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<connection>
<GID>573</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-4,434.5,3.5</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>0.5 5</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434.5,3.5,449,3.5</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection>
<intersection>448 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>448,-2.5,448,3.5</points>
<intersection>-2.5 4</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>448,-2.5,455.5,-2.5</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>448 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>427.5,0.5,434.5,0.5</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-15.5,434.5,-10</points>
<connection>
<GID>560</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-15.5,448.5,-15.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection>
<intersection>447.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>447.5,-23,447.5,-15.5</points>
<intersection>-23 3</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>447.5,-23,457,-23</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>447.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,-42.5,445.5,1.5</points>
<intersection>-42.5 2</intersection>
<intersection>-17.5 1</intersection>
<intersection>1.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,-17.5,448.5,-17.5</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443,-42.5,445.5,-42.5</points>
<connection>
<GID>566</GID>
<name>OUT_0</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>445.5,1.5,449,1.5</points>
<connection>
<GID>523</GID>
<name>IN_1</name></connection>
<intersection>445.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,0.5,467,2.5</points>
<intersection>0.5 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,0.5,513.5,0.5</points>
<connection>
<GID>507</GID>
<name>clock</name></connection>
<intersection>467 0</intersection>
<intersection>513.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>455,2.5,467,2.5</points>
<connection>
<GID>523</GID>
<name>OUT</name></connection>
<intersection>467 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>513.5,0.5,513.5,1</points>
<connection>
<GID>509</GID>
<name>clock</name></connection>
<intersection>0.5 1</intersection>
<intersection>1 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>513.5,1,575,1</points>
<connection>
<GID>511</GID>
<name>clock</name></connection>
<intersection>513.5 3</intersection>
<intersection>575 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>575,1,575,1.5</points>
<connection>
<GID>513</GID>
<name>clock</name></connection>
<intersection>1 4</intersection></vsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466.5,-23,466.5,-16.5</points>
<intersection>-23 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>466.5,-23,512.5,-23</points>
<connection>
<GID>515</GID>
<name>clock</name></connection>
<intersection>466.5 0</intersection>
<intersection>512.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>454.5,-16.5,466.5,-16.5</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<intersection>466.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>512.5,-23,512.5,-22.5</points>
<connection>
<GID>517</GID>
<name>clock</name></connection>
<intersection>-23 1</intersection>
<intersection>-22.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>512.5,-22.5,575,-22.5</points>
<connection>
<GID>519</GID>
<name>clock</name></connection>
<intersection>512.5 3</intersection>
<intersection>575 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>575,-23,575,-22.5</points>
<connection>
<GID>521</GID>
<name>clock</name></connection>
<intersection>-22.5 4</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>33.2304,600.093,1257.23,-4.90692</PageViewport></page 2>
<page 3>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 3>
<page 4>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 4>
<page 5>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 5>
<page 6>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 6>
<page 7>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 7>
<page 8>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 8>
<page 9>
<PageViewport>-0.00025201,384.093,1224,-220.907</PageViewport></page 9></circuit>