<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-47.1487,503.125,1176.85,-101.875</PageViewport>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW</type>
<position>108.5,31</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>66.5,29</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_AND2</type>
<position>67,4</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>68,-23</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>67.5,-47</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_DFF_LOW</type>
<position>120,31</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_INVERTER</type>
<position>52,-0.5</position>
<input>
<ID>IN_0</ID>100 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_INVERTER</type>
<position>40,-29</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_DFF_LOW</type>
<position>132,31</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>56 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>146,31</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>57 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_DFF_LOW</type>
<position>157,31</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_DFF_LOW</type>
<position>184,30</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>61 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_DFF_LOW</type>
<position>212,29.5</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>63 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_DFF_LOW</type>
<position>108.5,5</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_DFF_LOW</type>
<position>120.5,5</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_DFF_LOW</type>
<position>96,31</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_DFF_LOW</type>
<position>94.5,5</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_DFF_LOW</type>
<position>94.5,-21</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_DFF_LOW</type>
<position>95,-47</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_DFF_LOW</type>
<position>132.5,5</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_DFF_LOW</type>
<position>146.5,5</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_DFF_LOW</type>
<position>157,5.5</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>192,8.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>71 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>210.5,4.5</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>72 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_DFF_LOW</type>
<position>109,-21</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>119.5,-20.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>32.5,-22.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>134,-20.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>39.5,9.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_DFF_LOW</type>
<position>145.5,-21</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_DFF_LOW</type>
<position>158.5,-21</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>169,-20.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-21.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_DFF_LOW</type>
<position>109.5,-47</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_DFF_LOW</type>
<position>122,-47</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_DFF_LOW</type>
<position>132.5,-47</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_DFF_LOW</type>
<position>145.5,-47.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>158.5,-47.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_DFF_LOW</type>
<position>169.5,-47.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-47</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>79,28</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>40.5,-66</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>BA_TRI_STATE</type>
<position>231,1.5</position>
<input>
<ID>ENABLE_0</ID>64 </input>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>79.5,3</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>78,-33.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>BA_TRI_STATE</type>
<position>231,22.5</position>
<input>
<ID>ENABLE_0</ID>13 </input>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_TRI_STATE</type>
<position>101,-66.5</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>79,-53.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>58,-53.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>BA_TRI_STATE</type>
<position>89,-66</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>BA_TRI_STATE</type>
<position>199.5,23</position>
<input>
<ID>ENABLE_0</ID>16 </input>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>55</ID>
<type>BA_TRI_STATE</type>
<position>114.5,-66</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>56</ID>
<type>BA_TRI_STATE</type>
<position>100,40</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>57</ID>
<type>BA_TRI_STATE</type>
<position>127.5,-66</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_TRI_STATE</type>
<position>137.5,-66</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_TRI_STATE</type>
<position>113,40</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>61</ID>
<type>BA_TRI_STATE</type>
<position>151.5,-66</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_TRI_STATE</type>
<position>201.5,0</position>
<input>
<ID>ENABLE_0</ID>15 </input>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>63</ID>
<type>BA_TRI_STATE</type>
<position>124.5,40</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_TRI_STATE</type>
<position>179.5,-66</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_TRI_STATE</type>
<position>136.5,40</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>67</ID>
<type>BA_TRI_STATE</type>
<position>205,-68.5</position>
<input>
<ID>ENABLE_0</ID>21 </input>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>90,-77.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>100.5,-77</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>114.5,-78</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>127.5,-77</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>137.5,-77.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>151.5,-76.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>163,-76.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>174,-76.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>77</ID>
<type>BA_TRI_STATE</type>
<position>150,40</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>79</ID>
<type>BA_TRI_STATE</type>
<position>161.5,40</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>81</ID>
<type>BA_TRI_STATE</type>
<position>202.5,39</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>83</ID>
<type>BA_TRI_STATE</type>
<position>231,41</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>33,39</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>100,53</position>
<input>
<ID>N_in2</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>113,53</position>
<input>
<ID>N_in2</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>GA_LED</type>
<position>124.5,53</position>
<input>
<ID>N_in2</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>136.5,53</position>
<input>
<ID>N_in2</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>150,52.5</position>
<input>
<ID>N_in1</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>GA_LED</type>
<position>161.5,52.5</position>
<input>
<ID>N_in2</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>171.5,52.5</position>
<input>
<ID>N_in2</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>183.5,52.5</position>
<input>
<ID>N_in1</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>97.5,23.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>BA_TRI_STATE</type>
<position>81,19</position>
<input>
<ID>ENABLE_0</ID>7 </input>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND2</type>
<position>110.5,23.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>122,23</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>BA_TRI_STATE</type>
<position>81,-7.5</position>
<input>
<ID>ENABLE_0</ID>6 </input>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>134.5,23</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>147.5,23</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>159.5,23.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>191,23</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>219.5,25.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>96,-4</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND2</type>
<position>110.5,-4</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>121.5,-3.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>133,-3</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>148,-4</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND2</type>
<position>160,-4</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_AND2</type>
<position>194,0</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_AND2</type>
<position>218.5,-6</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,3.5,207.5,3.5</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>82.5 32</intersection>
<intersection>91.5 26</intersection>
<intersection>105.5 27</intersection>
<intersection>117.5 28</intersection>
<intersection>129.5 29</intersection>
<intersection>143.5 30</intersection>
<intersection>154 7</intersection>
<intersection>188 31</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>154,3.5,154,4.5</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>91.5,3.5,91.5,4</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>105.5,3.5,105.5,4</points>
<connection>
<GID>15</GID>
<name>clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>117.5,3.5,117.5,4</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>129.5,3.5,129.5,4</points>
<connection>
<GID>21</GID>
<name>clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>143.5,3.5,143.5,4</points>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>188,3.5,188,7.5</points>
<intersection>3.5 1</intersection>
<intersection>7.5 33</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>82.5,3,82.5,3.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>188,7.5,189,7.5</points>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<intersection>188 31</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-52.5,73,-47</points>
<intersection>-52.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-52.5,76,-52.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-47,73,-47</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-53.5,76,-53.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>73 4</intersection>
<intersection>76 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>73,-53.5,73,27</points>
<intersection>-53.5 1</intersection>
<intersection>-34.5 7</intersection>
<intersection>2 6</intersection>
<intersection>27 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>73,27,76,27</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>73 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>73,2,76.5,2</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>73 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>73,-34.5,75,-34.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>73 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>76,-54.5,76,-53.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-32.5,73,-23</points>
<intersection>-32.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-32.5,75,-32.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-23,73,-23</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,4,81,4</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>81 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81,-5.5,81,4</points>
<connection>
<GID>110</GID>
<name>ENABLE_0</name></connection>
<intersection>4 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,29,81,29</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>81 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>81,21,81,29</points>
<connection>
<GID>106</GID>
<name>ENABLE_0</name></connection>
<intersection>29 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-33.5,177.5,-33.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>91.5 4</intersection>
<intersection>106 5</intersection>
<intersection>131 7</intersection>
<intersection>142.5 8</intersection>
<intersection>155.5 9</intersection>
<intersection>177.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177.5,-33.5,177.5,-22.5</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>91.5,-33.5,91.5,-22</points>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>106,-33.5,106,-21.5</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection>
<intersection>-21.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>106,-21.5,116.5,-21.5</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>106 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>131,-33.5,131,-21.5</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>142.5,-33.5,142.5,-22</points>
<connection>
<GID>31</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>155.5,-33.5,155.5,-21.5</points>
<connection>
<GID>32</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection>
<intersection>-21.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>155.5,-21.5,166,-21.5</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>155.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-53.5,177.5,-53.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>92 4</intersection>
<intersection>106.5 5</intersection>
<intersection>119 6</intersection>
<intersection>129.5 7</intersection>
<intersection>142.5 8</intersection>
<intersection>155.5 9</intersection>
<intersection>166.5 10</intersection>
<intersection>177.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177.5,-53.5,177.5,-48</points>
<connection>
<GID>41</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>92,-53.5,92,-48</points>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>106.5,-53.5,106.5,-48</points>
<connection>
<GID>35</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>119,-53.5,119,-48</points>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>129.5,-53.5,129.5,-48</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>142.5,-53.5,142.5,-48.5</points>
<connection>
<GID>38</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>155.5,-53.5,155.5,-48.5</points>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>166.5,-53.5,166.5,-48.5</points>
<connection>
<GID>40</GID>
<name>clock</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,22.5,226,25.5</points>
<intersection>22.5 2</intersection>
<intersection>25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,25.5,226,25.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>226,22.5,229,22.5</points>
<connection>
<GID>48</GID>
<name>ENABLE_0</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234,4,234,38</points>
<intersection>4 9</intersection>
<intersection>25 8</intersection>
<intersection>38 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>231,25,234,25</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>234 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>231,4,234,4</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>234 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>231,38,234,38</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>234 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>197,0,199.5,0</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,23,197.5,23</points>
<connection>
<GID>54</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,30.5,202.5,36</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>30.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>202,2.5,202,30.5</points>
<intersection>2.5 3</intersection>
<intersection>25.5 4</intersection>
<intersection>30.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>202,30.5,202.5,30.5</points>
<intersection>202 1</intersection>
<intersection>202.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>201.5,2.5,202,2.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>202 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199.5,25.5,202,25.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>202 1</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,28,84.5,30</points>
<intersection>28 2</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,30,181,30</points>
<connection>
<GID>11</GID>
<name>clock</name></connection>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<connection>
<GID>9</GID>
<name>clock</name></connection>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<connection>
<GID>17</GID>
<name>clock</name></connection>
<intersection>84.5 0</intersection>
<intersection>181 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,28,84.5,28</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>181,28.5,181,30</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>28.5 9</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>181,28.5,209,28.5</points>
<connection>
<GID>13</GID>
<name>clock</name></connection>
<intersection>181 8</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-59.5,170.5,-59.5</points>
<intersection>86 4</intersection>
<intersection>98.5 5</intersection>
<intersection>111.5 6</intersection>
<intersection>123 7</intersection>
<intersection>135.5 8</intersection>
<intersection>148 9</intersection>
<intersection>158.5 10</intersection>
<intersection>170.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>170.5,-59.5,170.5,-59</points>
<intersection>-59.5 1</intersection>
<intersection>-59 17</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>86,-66,86,-59.5</points>
<intersection>-66 11</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>98.5,-66.5,98.5,-59.5</points>
<intersection>-66.5 21</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>111.5,-66,111.5,-59.5</points>
<intersection>-66 13</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>123,-66,123,-59.5</points>
<intersection>-66 14</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>135.5,-66,135.5,-59.5</points>
<connection>
<GID>59</GID>
<name>ENABLE_0</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>148,-66,148,-59.5</points>
<intersection>-66 15</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>158.5,-66,158.5,-59.5</points>
<intersection>-66 16</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>42.5,-66,87,-66</points>
<connection>
<GID>53</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>86 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>111.5,-66,112.5,-66</points>
<connection>
<GID>55</GID>
<name>ENABLE_0</name></connection>
<intersection>111.5 6</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>123,-66,125.5,-66</points>
<connection>
<GID>57</GID>
<name>ENABLE_0</name></connection>
<intersection>123 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>148,-66,149.5,-66</points>
<connection>
<GID>61</GID>
<name>ENABLE_0</name></connection>
<intersection>148 9</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>158.5,-66,177.5,-66</points>
<connection>
<GID>65</GID>
<name>ENABLE_0</name></connection>
<intersection>158.5 10</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>170.5,-59,203,-59</points>
<intersection>170.5 3</intersection>
<intersection>203 25</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>98.5,-66.5,99,-66.5</points>
<connection>
<GID>49</GID>
<name>ENABLE_0</name></connection>
<intersection>98.5 5</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>203,-68.5,203,-59</points>
<connection>
<GID>67</GID>
<name>ENABLE_0</name></connection>
<intersection>-59 17</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-75.5,90,-69</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-69 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>89,-69,90,-69</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-76,101,-69.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-76 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>100.5,-76,101,-76</points>
<intersection>100.5 14</intersection>
<intersection>101 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>100.5,-76,100.5,-75</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-76 13</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-76,114.5,-69</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-75,127.5,-69</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-75.5,137.5,-69</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-74.5,151.5,-69</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,39,66.5,40</points>
<intersection>39 2</intersection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,40,229,40</points>
<connection>
<GID>79</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>77</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>66</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>63</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>60</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>56</GID>
<name>ENABLE_0</name></connection>
<intersection>66.5 0</intersection>
<intersection>74 8</intersection>
<intersection>200.5 12</intersection>
<intersection>229 13</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,39,66.5,39</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>74,-7.5,74,40</points>
<intersection>-7.5 10</intersection>
<intersection>19 11</intersection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>74,-7.5,78,-7.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>74 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>74,19,78,19</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>74 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>200.5,39,200.5,40</points>
<connection>
<GID>81</GID>
<name>ENABLE_0</name></connection>
<intersection>40 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>229,40,229,41</points>
<connection>
<GID>83</GID>
<name>ENABLE_0</name></connection>
<intersection>40 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-74.5,179.5,-69</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-74.5,179.5,-74.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-74.5,205,-74.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>205 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>205,-74.5,205,-71.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,42.5,100,52</points>
<connection>
<GID>87</GID>
<name>N_in2</name></connection>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,42.5,113,52</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>89</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,19,89,22.5</points>
<intersection>19 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,22.5,119,22.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>89 0</intersection>
<intersection>119 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,19,89,19</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>89 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>119,22,119,22.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>22 5</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>119,22,216.5,22</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>119 4</intersection>
<intersection>156.5 7</intersection>
<intersection>216.5 10</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>156.5,22,156.5,22.5</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>22 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>216.5,22,216.5,24.5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>22 5</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-7.5,88,-5</points>
<intersection>-7.5 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-5,118.5,-5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>88 0</intersection>
<intersection>118.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-7.5,88,-7.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>118.5,-5,118.5,-4</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-5 1</intersection>
<intersection>-4 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>118.5,-4,145,-4</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>118.5 4</intersection>
<intersection>145 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>145,-5,145,-4</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-5 7</intersection>
<intersection>-4 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>145,-5,157,-5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>145 6</intersection>
<intersection>156.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>156.5,-12.5,156.5,-5</points>
<intersection>-12.5 10</intersection>
<intersection>-5 7</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>203,-12.5,203,-7</points>
<intersection>-12.5 10</intersection>
<intersection>-7 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>156.5,-12.5,203,-12.5</points>
<intersection>156.5 8</intersection>
<intersection>191 12</intersection>
<intersection>203 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>203,-7,215.5,-7</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>203 9</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>191,-12.5,191,-1</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>-12.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,42.5,124.5,52</points>
<connection>
<GID>91</GID>
<name>N_in2</name></connection>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,42.5,136.5,52</points>
<connection>
<GID>93</GID>
<name>N_in2</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,42.5,150,52.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,52.5,151,52.5</points>
<connection>
<GID>95</GID>
<name>N_in1</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,42.5,161.5,51.5</points>
<connection>
<GID>97</GID>
<name>N_in2</name></connection>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,47,171.5,51.5</points>
<connection>
<GID>99</GID>
<name>N_in2</name></connection>
<intersection>47 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>202.5,41.5,202.5,47</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>47 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>171.5,47,202.5,47</points>
<intersection>171.5 0</intersection>
<intersection>202.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-63.5,88,33</points>
<intersection>-63.5 5</intersection>
<intersection>-45 4</intersection>
<intersection>-19 3</intersection>
<intersection>7 2</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,33,93,33</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88,7,91.5,7</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>88,-19,91.5,-19</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>88,-45,92,-45</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>88,-63.5,89,-63.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-64,102,33</points>
<intersection>-64 8</intersection>
<intersection>-45 4</intersection>
<intersection>-19 3</intersection>
<intersection>7 2</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,33,105.5,33</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,7,105.5,7</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,-19,106,-19</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102,-45,106.5,-45</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>101,-64,102,-64</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-63.5,116,33</points>
<intersection>-63.5 9</intersection>
<intersection>-45 6</intersection>
<intersection>-18.5 5</intersection>
<intersection>7 3</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,33,117,33</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>116,7,117.5,7</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>116,-18.5,116.5,-18.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>116,-45,119,-45</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114.5,-63.5,116,-63.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-63.5,127.5,33</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-45 4</intersection>
<intersection>-18.5 3</intersection>
<intersection>7 2</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,33,129,33</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,7,129.5,7</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>127.5,-18.5,131,-18.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>127.5,-45,129.5,-45</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-63.5,139.5,33</points>
<intersection>-63.5 6</intersection>
<intersection>-45.5 4</intersection>
<intersection>-19 3</intersection>
<intersection>7 2</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,33,143,33</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,7,143.5,7</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>139.5,-19,142.5,-19</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>139.5,-45.5,142.5,-45.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>137.5,-63.5,139.5,-63.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-63.5,151.5,33</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>-45.5 4</intersection>
<intersection>-19 3</intersection>
<intersection>7.5 2</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,33,154,33</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>151.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151.5,7.5,154,7.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>151.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>151.5,-19,155.5,-19</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>151.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>151.5,-45.5,155.5,-45.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>151.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-63.5,179.5,32</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-45.5 4</intersection>
<intersection>-18.5 3</intersection>
<intersection>10.5 2</intersection>
<intersection>32 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>179.5,10.5,189,10.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>166,-18.5,179.5,-18.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>166.5,-45.5,179.5,-45.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>179.5,32,181,32</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-66,205,31.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>-45 6</intersection>
<intersection>-19.5 5</intersection>
<intersection>6.5 4</intersection>
<intersection>31.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>205,6.5,207.5,6.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>177.5,-19.5,205,-19.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>177.5,-45,205,-45</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205,31.5,209,31.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231,43.5,231,52.5</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,52.5,231,52.5</points>
<connection>
<GID>103</GID>
<name>N_in1</name></connection>
<intersection>231 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,24.5,96.5,33</points>
<intersection>24.5 1</intersection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94.5,24.5,96.5,24.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,33,99,33</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-4,100,37</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-4 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,23.5,100.5,23.5</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-4,100,-4</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,24.5,109.5,33</points>
<intersection>24.5 1</intersection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,24.5,109.5,24.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,33,111.5,33</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,23.5,113,37</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,23.5,113.5,23.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>113 0</intersection>
<intersection>113.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>113.5,-4,113.5,23.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,24,121,33</points>
<intersection>24 1</intersection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,24,121,24</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,33,123,33</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-3.5,124.5,37</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,23,125,23</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-3,136.5,37</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-3 2</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,23,137.5,23</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>136,-3,136.5,-3</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,24,133,33</points>
<intersection>24 1</intersection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,24,133,24</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,33,135,33</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,24,146.5,33</points>
<intersection>24 1</intersection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,24,146.5,24</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,33,149,33</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,23,150,37</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,23,151,23</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>150 0</intersection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-4,151,23</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>23 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,24.5,158,33</points>
<intersection>24.5 1</intersection>
<intersection>33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,24.5,158,24.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>158,33,160,33</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,23.5,161.5,37</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,23.5,163,23.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>161.5 0</intersection>
<intersection>163 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>163,-4,163,23.5</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,20,188,32</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection>
<intersection>32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>187,32,188,32</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188,20,199.5,20</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>188 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,19,216,31.5</points>
<intersection>19 3</intersection>
<intersection>26.5 1</intersection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,26.5,216.5,26.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>215,31.5,216,31.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>216,19,231,19</points>
<intersection>216 0</intersection>
<intersection>231 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>231,19,231,19.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-6,225,1.5</points>
<intersection>-6 2</intersection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1.5,229,1.5</points>
<connection>
<GID>44</GID>
<name>ENABLE_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>221.5,-6,225,-6</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-3,92,7</points>
<intersection>-3 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-3,93,-3</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,7,97.5,7</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3,109.5,7</points>
<intersection>-3 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-3,109.5,-3</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,7,111.5,7</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-2.5,121,7</points>
<intersection>-2.5 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-2.5,121,-2.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,7,123.5,7</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-2,132.5,7</points>
<intersection>-2 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-2,132.5,-2</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,7,135.5,7</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-3,147,7</points>
<intersection>-3 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-3,147,-3</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147,7,149.5,7</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>147 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-3,158.5,7.5</points>
<intersection>-3 1</intersection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-3,158.5,-3</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>158.5,7.5,160,7.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-3,194,4.5</points>
<intersection>-3 4</intersection>
<intersection>1 1</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,1,194,1</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194,4.5,196,4.5</points>
<intersection>194 0</intersection>
<intersection>196 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>196,4.5,196,10.5</points>
<intersection>4.5 2</intersection>
<intersection>10.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>194,-3,201.5,-3</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>195,10.5,196,10.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>196 3</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-2,214,6.5</points>
<intersection>-2 1</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214,-2,231,-2</points>
<intersection>214 0</intersection>
<intersection>215.5 5</intersection>
<intersection>231 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,6.5,214,6.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>214 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>231,-2,231,-1.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>215.5,-5,215.5,-2</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-46,52,-3.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-46 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-22,65,-22</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52,-46,64.5,-46</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,2.5,52,30</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>5 3</intersection>
<intersection>9.5 1</intersection>
<intersection>30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,9.5,52,9.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,30,63.5,30</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,5,64,5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-26,40,-24</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-24,65,-24</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>34.5 5</intersection>
<intersection>40 0</intersection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58,-24,58,28</points>
<intersection>-24 1</intersection>
<intersection>28 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>58,28,63.5,28</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>34.5,-24,34.5,-22.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-48,40,3</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-48 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-48,64.5,-48</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,3,64,3</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-319.327,74.0241,-101.482,-33.6529</PageViewport>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>32,-5066</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>BA_TRI_STATE</type>
<position>42.5,-5066</position>
<input>
<ID>ENABLE_0</ID>8 </input>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>112,278</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>AE_DFF_LOW</type>
<position>28,284.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>172 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>252</ID>
<type>BA_TRI_STATE</type>
<position>52.5,278</position>
<input>
<ID>ENABLE_0</ID>171 </input>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>38,278</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_DFF_LOW</type>
<position>101.5,284.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>174 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>255</ID>
<type>BA_TRI_STATE</type>
<position>126,278</position>
<input>
<ID>ENABLE_0</ID>173 </input>
<input>
<ID>IN_0</ID>174 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>270,276</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>AE_DFF_LOW</type>
<position>186,284.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>176 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>258</ID>
<type>BA_TRI_STATE</type>
<position>210.5,276</position>
<input>
<ID>ENABLE_0</ID>175 </input>
<input>
<ID>IN_0</ID>176 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_AND2</type>
<position>196,276</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_DFF_LOW</type>
<position>260.5,284.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>178 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>261</ID>
<type>BA_TRI_STATE</type>
<position>284,276</position>
<input>
<ID>ENABLE_0</ID>177 </input>
<input>
<ID>IN_0</ID>178 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>435,274.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_DFF_LOW</type>
<position>351,284.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>180 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>264</ID>
<type>BA_TRI_STATE</type>
<position>375.5,274.5</position>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>361,274.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_DFF_LOW</type>
<position>424.5,284.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>182 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>267</ID>
<type>BA_TRI_STATE</type>
<position>449,274.5</position>
<input>
<ID>ENABLE_0</ID>181 </input>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>593,272.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_DFF_LOW</type>
<position>509,284.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>184 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>270</ID>
<type>BA_TRI_STATE</type>
<position>533.5,272.5</position>
<input>
<ID>ENABLE_0</ID>183 </input>
<input>
<ID>IN_0</ID>184 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND2</type>
<position>519,272.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>AE_DFF_LOW</type>
<position>582.5,284.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>186 </output>
<input>
<ID>clock</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>273</ID>
<type>BA_TRI_STATE</type>
<position>607,272.5</position>
<input>
<ID>ENABLE_0</ID>185 </input>
<input>
<ID>IN_0</ID>186 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_AND2</type>
<position>-3.5,283.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>BA_TRI_STATE</type>
<position>-25,264.5</position>
<input>
<ID>ENABLE_0</ID>169 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>109,368</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AE_DFF_LOW</type>
<position>25,374.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>191 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>278</ID>
<type>BA_TRI_STATE</type>
<position>49.5,368</position>
<input>
<ID>ENABLE_0</ID>190 </input>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_AND2</type>
<position>35,368</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AE_DFF_LOW</type>
<position>98.5,374.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>193 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>281</ID>
<type>BA_TRI_STATE</type>
<position>123,368</position>
<input>
<ID>ENABLE_0</ID>192 </input>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_AND2</type>
<position>267,366</position>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>AE_DFF_LOW</type>
<position>183,374.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>195 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>284</ID>
<type>BA_TRI_STATE</type>
<position>207.5,366</position>
<input>
<ID>ENABLE_0</ID>194 </input>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>285</ID>
<type>AA_AND2</type>
<position>193,366</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_DFF_LOW</type>
<position>257.5,374.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>197 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>287</ID>
<type>BA_TRI_STATE</type>
<position>281,366</position>
<input>
<ID>ENABLE_0</ID>196 </input>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_AND2</type>
<position>432,364.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_DFF_LOW</type>
<position>348,374.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>199 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>290</ID>
<type>BA_TRI_STATE</type>
<position>372.5,364.5</position>
<input>
<ID>ENABLE_0</ID>198 </input>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_AND2</type>
<position>358,364.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_DFF_LOW</type>
<position>421.5,374.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>201 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>293</ID>
<type>BA_TRI_STATE</type>
<position>446,364.5</position>
<input>
<ID>ENABLE_0</ID>200 </input>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_AND2</type>
<position>590,362.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>AE_DFF_LOW</type>
<position>506,374.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>203 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>296</ID>
<type>BA_TRI_STATE</type>
<position>530.5,362.5</position>
<input>
<ID>ENABLE_0</ID>202 </input>
<input>
<ID>IN_0</ID>203 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_AND2</type>
<position>516,362.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>AE_DFF_LOW</type>
<position>579.5,374.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>205 </output>
<input>
<ID>clock</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>299</ID>
<type>BA_TRI_STATE</type>
<position>604,362.5</position>
<input>
<ID>ENABLE_0</ID>204 </input>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND2</type>
<position>-6.5,373.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>BA_TRI_STATE</type>
<position>-28,354.5</position>
<input>
<ID>ENABLE_0</ID>188 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>189 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND2</type>
<position>116,110</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_DFF_LOW</type>
<position>32,116.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>210 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>304</ID>
<type>BA_TRI_STATE</type>
<position>56.5,110</position>
<input>
<ID>ENABLE_0</ID>209 </input>
<input>
<ID>IN_0</ID>210 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_AND2</type>
<position>42,110</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>105.5,116.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>212 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>BA_TRI_STATE</type>
<position>130,110</position>
<input>
<ID>ENABLE_0</ID>211 </input>
<input>
<ID>IN_0</ID>212 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_AND2</type>
<position>274,108</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_DFF_LOW</type>
<position>190,116.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>214 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>310</ID>
<type>BA_TRI_STATE</type>
<position>214.5,108</position>
<input>
<ID>ENABLE_0</ID>213 </input>
<input>
<ID>IN_0</ID>214 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_AND2</type>
<position>200,108</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>312</ID>
<type>AE_DFF_LOW</type>
<position>264.5,116.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>216 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>313</ID>
<type>BA_TRI_STATE</type>
<position>288,108</position>
<input>
<ID>ENABLE_0</ID>215 </input>
<input>
<ID>IN_0</ID>216 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>439,106.5</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AE_DFF_LOW</type>
<position>355,116.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>218 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>316</ID>
<type>BA_TRI_STATE</type>
<position>386,106</position>
<input>
<ID>ENABLE_0</ID>217 </input>
<input>
<ID>IN_0</ID>218 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_AND2</type>
<position>365,106.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_DFF_LOW</type>
<position>428.5,116.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>220 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>319</ID>
<type>BA_TRI_STATE</type>
<position>453,106.5</position>
<input>
<ID>ENABLE_0</ID>219 </input>
<input>
<ID>IN_0</ID>220 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>597,104.5</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AE_DFF_LOW</type>
<position>513,116.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>222 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>322</ID>
<type>BA_TRI_STATE</type>
<position>537.5,104.5</position>
<input>
<ID>ENABLE_0</ID>221 </input>
<input>
<ID>IN_0</ID>222 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>323</ID>
<type>AA_AND2</type>
<position>523,104.5</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_DFF_LOW</type>
<position>586.5,116.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>224 </output>
<input>
<ID>clock</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>325</ID>
<type>BA_TRI_STATE</type>
<position>611,104.5</position>
<input>
<ID>ENABLE_0</ID>223 </input>
<input>
<ID>IN_0</ID>224 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>326</ID>
<type>AA_AND2</type>
<position>0.5,115.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>BA_TRI_STATE</type>
<position>-21,96.5</position>
<input>
<ID>ENABLE_0</ID>207 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>208 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>113,200</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AE_DFF_LOW</type>
<position>29,206.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>229 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>330</ID>
<type>BA_TRI_STATE</type>
<position>53.5,200</position>
<input>
<ID>ENABLE_0</ID>228 </input>
<input>
<ID>IN_0</ID>229 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_AND2</type>
<position>39,200</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_DFF_LOW</type>
<position>102.5,206.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>231 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>333</ID>
<type>BA_TRI_STATE</type>
<position>127,200</position>
<input>
<ID>ENABLE_0</ID>230 </input>
<input>
<ID>IN_0</ID>231 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_AND2</type>
<position>271,198</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_DFF_LOW</type>
<position>187,206.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>233 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>336</ID>
<type>BA_TRI_STATE</type>
<position>211.5,198</position>
<input>
<ID>ENABLE_0</ID>232 </input>
<input>
<ID>IN_0</ID>233 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_AND2</type>
<position>197,198</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_DFF_LOW</type>
<position>261.5,206.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>235 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>339</ID>
<type>BA_TRI_STATE</type>
<position>285,198</position>
<input>
<ID>ENABLE_0</ID>234 </input>
<input>
<ID>IN_0</ID>235 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>436,196.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AE_DFF_LOW</type>
<position>352,206.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>237 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>342</ID>
<type>BA_TRI_STATE</type>
<position>376.5,196.5</position>
<input>
<ID>ENABLE_0</ID>236 </input>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_AND2</type>
<position>362,196.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_DFF_LOW</type>
<position>425.5,206.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>239 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>345</ID>
<type>BA_TRI_STATE</type>
<position>450,196.5</position>
<input>
<ID>ENABLE_0</ID>238 </input>
<input>
<ID>IN_0</ID>239 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>346</ID>
<type>AA_AND2</type>
<position>594,194.5</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>AE_DFF_LOW</type>
<position>510,206.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>241 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>348</ID>
<type>BA_TRI_STATE</type>
<position>534.5,194.5</position>
<input>
<ID>ENABLE_0</ID>240 </input>
<input>
<ID>IN_0</ID>241 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_AND2</type>
<position>520,194.5</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_DFF_LOW</type>
<position>583.5,206.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>243 </output>
<input>
<ID>clock</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>351</ID>
<type>BA_TRI_STATE</type>
<position>608,194.5</position>
<input>
<ID>ENABLE_0</ID>242 </input>
<input>
<ID>IN_0</ID>243 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND2</type>
<position>-2.5,205.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>BA_TRI_STATE</type>
<position>-24,186.5</position>
<input>
<ID>ENABLE_0</ID>226 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>114,-98</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AE_DFF_LOW</type>
<position>30,-91.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>248 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>356</ID>
<type>BA_TRI_STATE</type>
<position>54.5,-98</position>
<input>
<ID>ENABLE_0</ID>247 </input>
<input>
<ID>IN_0</ID>248 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_AND2</type>
<position>40,-98</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-91.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>250 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>359</ID>
<type>BA_TRI_STATE</type>
<position>128,-98</position>
<input>
<ID>ENABLE_0</ID>249 </input>
<input>
<ID>IN_0</ID>250 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_AND2</type>
<position>272,-100</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AE_DFF_LOW</type>
<position>188,-91.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>252 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>362</ID>
<type>BA_TRI_STATE</type>
<position>212.5,-100</position>
<input>
<ID>ENABLE_0</ID>251 </input>
<input>
<ID>IN_0</ID>252 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>198,-100</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-91.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>254 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>365</ID>
<type>BA_TRI_STATE</type>
<position>286,-100</position>
<input>
<ID>ENABLE_0</ID>253 </input>
<input>
<ID>IN_0</ID>254 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>366</ID>
<type>AA_AND2</type>
<position>437,-101.5</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AE_DFF_LOW</type>
<position>353,-91.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>256 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>368</ID>
<type>BA_TRI_STATE</type>
<position>377.5,-101.5</position>
<input>
<ID>ENABLE_0</ID>255 </input>
<input>
<ID>IN_0</ID>256 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_AND2</type>
<position>363,-101.5</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>AE_DFF_LOW</type>
<position>426.5,-91.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>258 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>371</ID>
<type>BA_TRI_STATE</type>
<position>451,-101.5</position>
<input>
<ID>ENABLE_0</ID>257 </input>
<input>
<ID>IN_0</ID>258 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>595,-103.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AE_DFF_LOW</type>
<position>511,-91.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>260 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>374</ID>
<type>BA_TRI_STATE</type>
<position>535.5,-103.5</position>
<input>
<ID>ENABLE_0</ID>259 </input>
<input>
<ID>IN_0</ID>260 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_AND2</type>
<position>521,-103.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>AE_DFF_LOW</type>
<position>584.5,-91.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>262 </output>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>377</ID>
<type>BA_TRI_STATE</type>
<position>609,-103.5</position>
<input>
<ID>ENABLE_0</ID>261 </input>
<input>
<ID>IN_0</ID>262 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_AND2</type>
<position>-1.5,-92.5</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>BA_TRI_STATE</type>
<position>-23,-111.5</position>
<input>
<ID>ENABLE_0</ID>245 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>246 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_AND2</type>
<position>111,-8</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AE_DFF_LOW</type>
<position>27,-1.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>267 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>382</ID>
<type>BA_TRI_STATE</type>
<position>51.5,-8</position>
<input>
<ID>ENABLE_0</ID>266 </input>
<input>
<ID>IN_0</ID>267 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_AND2</type>
<position>37,-8</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-1.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>269 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>385</ID>
<type>BA_TRI_STATE</type>
<position>125,-8</position>
<input>
<ID>ENABLE_0</ID>268 </input>
<input>
<ID>IN_0</ID>269 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>386</ID>
<type>AA_AND2</type>
<position>269,-10</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>272 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>387</ID>
<type>AE_DFF_LOW</type>
<position>185,-1.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>271 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>388</ID>
<type>BA_TRI_STATE</type>
<position>209.5,-10</position>
<input>
<ID>ENABLE_0</ID>270 </input>
<input>
<ID>IN_0</ID>271 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>389</ID>
<type>AA_AND2</type>
<position>195,-10</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-1.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>273 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>391</ID>
<type>BA_TRI_STATE</type>
<position>283,-10</position>
<input>
<ID>ENABLE_0</ID>272 </input>
<input>
<ID>IN_0</ID>273 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>392</ID>
<type>AA_AND2</type>
<position>434,-11.5</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>AE_DFF_LOW</type>
<position>350,-1.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>275 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>394</ID>
<type>BA_TRI_STATE</type>
<position>374.5,-11.5</position>
<input>
<ID>ENABLE_0</ID>274 </input>
<input>
<ID>IN_0</ID>275 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_AND2</type>
<position>360,-11.5</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>AE_DFF_LOW</type>
<position>423.5,-1.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>277 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>397</ID>
<type>BA_TRI_STATE</type>
<position>448,-11.5</position>
<input>
<ID>ENABLE_0</ID>276 </input>
<input>
<ID>IN_0</ID>277 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_AND2</type>
<position>592,-13.5</position>
<input>
<ID>IN_0</ID>281 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>AE_DFF_LOW</type>
<position>508,-1.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>279 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>400</ID>
<type>BA_TRI_STATE</type>
<position>532.5,-13.5</position>
<input>
<ID>ENABLE_0</ID>278 </input>
<input>
<ID>IN_0</ID>279 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>401</ID>
<type>AA_AND2</type>
<position>518,-13.5</position>
<input>
<ID>IN_0</ID>279 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>278 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>AE_DFF_LOW</type>
<position>581.5,-1.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>281 </output>
<input>
<ID>clock</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>403</ID>
<type>BA_TRI_STATE</type>
<position>606,-13.5</position>
<input>
<ID>ENABLE_0</ID>280 </input>
<input>
<ID>IN_0</ID>281 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>-4.5,-2.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>282 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>BA_TRI_STATE</type>
<position>-26,-21.5</position>
<input>
<ID>ENABLE_0</ID>264 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>265 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>118,-266</position>
<input>
<ID>IN_0</ID>288 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AE_DFF_LOW</type>
<position>34,-259.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>286 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>408</ID>
<type>BA_TRI_STATE</type>
<position>58.5,-266</position>
<input>
<ID>ENABLE_0</ID>285 </input>
<input>
<ID>IN_0</ID>286 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND2</type>
<position>44,-266</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>285 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_DFF_LOW</type>
<position>107.5,-259.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>288 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>411</ID>
<type>BA_TRI_STATE</type>
<position>132,-266</position>
<input>
<ID>ENABLE_0</ID>287 </input>
<input>
<ID>IN_0</ID>288 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_AND2</type>
<position>276,-268</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>291 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>413</ID>
<type>AE_DFF_LOW</type>
<position>192,-259.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>290 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>414</ID>
<type>BA_TRI_STATE</type>
<position>216.5,-268</position>
<input>
<ID>ENABLE_0</ID>289 </input>
<input>
<ID>IN_0</ID>290 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>415</ID>
<type>AA_AND2</type>
<position>202,-268</position>
<input>
<ID>IN_0</ID>290 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>289 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>AE_DFF_LOW</type>
<position>266.5,-259.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>292 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>417</ID>
<type>BA_TRI_STATE</type>
<position>290,-268</position>
<input>
<ID>ENABLE_0</ID>291 </input>
<input>
<ID>IN_0</ID>292 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_AND2</type>
<position>441,-269.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>295 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>AE_DFF_LOW</type>
<position>357,-259.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>294 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>420</ID>
<type>BA_TRI_STATE</type>
<position>381.5,-269.5</position>
<input>
<ID>ENABLE_0</ID>293 </input>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>421</ID>
<type>AA_AND2</type>
<position>367,-269.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>422</ID>
<type>AE_DFF_LOW</type>
<position>430.5,-259.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>296 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>423</ID>
<type>BA_TRI_STATE</type>
<position>455,-269.5</position>
<input>
<ID>ENABLE_0</ID>295 </input>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>424</ID>
<type>AA_AND2</type>
<position>599,-271.5</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>299 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>AE_DFF_LOW</type>
<position>515,-259.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>298 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>426</ID>
<type>BA_TRI_STATE</type>
<position>539.5,-271.5</position>
<input>
<ID>ENABLE_0</ID>297 </input>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>427</ID>
<type>AA_AND2</type>
<position>525,-271.5</position>
<input>
<ID>IN_0</ID>298 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>297 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>428</ID>
<type>AE_DFF_LOW</type>
<position>588.5,-259.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>300 </output>
<input>
<ID>clock</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>429</ID>
<type>BA_TRI_STATE</type>
<position>613,-271.5</position>
<input>
<ID>ENABLE_0</ID>299 </input>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>430</ID>
<type>AA_AND2</type>
<position>2.5,-260.5</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>431</ID>
<type>BA_TRI_STATE</type>
<position>-19,-279.5</position>
<input>
<ID>ENABLE_0</ID>283 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>284 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>432</ID>
<type>AA_AND2</type>
<position>115,-176</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>306 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>AE_DFF_LOW</type>
<position>31,-169.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>305 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>434</ID>
<type>BA_TRI_STATE</type>
<position>55.5,-176</position>
<input>
<ID>ENABLE_0</ID>304 </input>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>435</ID>
<type>AA_AND2</type>
<position>41,-176</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>304 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>AE_DFF_LOW</type>
<position>104.5,-169.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>307 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>437</ID>
<type>BA_TRI_STATE</type>
<position>129,-176</position>
<input>
<ID>ENABLE_0</ID>306 </input>
<input>
<ID>IN_0</ID>307 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>438</ID>
<type>AA_AND2</type>
<position>273,-178</position>
<input>
<ID>IN_0</ID>311 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>439</ID>
<type>AE_DFF_LOW</type>
<position>189,-169.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>309 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>440</ID>
<type>BA_TRI_STATE</type>
<position>213.5,-178</position>
<input>
<ID>ENABLE_0</ID>308 </input>
<input>
<ID>IN_0</ID>309 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>441</ID>
<type>AA_AND2</type>
<position>199,-178</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>442</ID>
<type>AE_DFF_LOW</type>
<position>263.5,-169.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>311 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>443</ID>
<type>BA_TRI_STATE</type>
<position>287,-178</position>
<input>
<ID>ENABLE_0</ID>310 </input>
<input>
<ID>IN_0</ID>311 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>444</ID>
<type>AA_AND2</type>
<position>438,-179.5</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>445</ID>
<type>AE_DFF_LOW</type>
<position>354,-169.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>313 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>446</ID>
<type>BA_TRI_STATE</type>
<position>378.5,-179.5</position>
<input>
<ID>ENABLE_0</ID>312 </input>
<input>
<ID>IN_0</ID>313 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>447</ID>
<type>AA_AND2</type>
<position>364,-179.5</position>
<input>
<ID>IN_0</ID>313 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>448</ID>
<type>AE_DFF_LOW</type>
<position>427.5,-169.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>315 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>449</ID>
<type>BA_TRI_STATE</type>
<position>452,-179.5</position>
<input>
<ID>ENABLE_0</ID>314 </input>
<input>
<ID>IN_0</ID>315 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_AND2</type>
<position>596,-181.5</position>
<input>
<ID>IN_0</ID>319 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>318 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>451</ID>
<type>AE_DFF_LOW</type>
<position>512,-169.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>317 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>452</ID>
<type>BA_TRI_STATE</type>
<position>536.5,-181.5</position>
<input>
<ID>ENABLE_0</ID>1463 </input>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_AND2</type>
<position>522,-181.5</position>
<input>
<ID>IN_0</ID>317 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>1463 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>AE_DFF_LOW</type>
<position>585.5,-169.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>319 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>455</ID>
<type>BA_TRI_STATE</type>
<position>610,-181.5</position>
<input>
<ID>ENABLE_0</ID>318 </input>
<input>
<ID>IN_0</ID>319 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>456</ID>
<type>AA_AND2</type>
<position>-0.5,-170.5</position>
<input>
<ID>IN_0</ID>302 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>457</ID>
<type>BA_TRI_STATE</type>
<position>-22,-189.5</position>
<input>
<ID>ENABLE_0</ID>302 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>303 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>459</ID>
<type>BE_DECODER_3x8</type>
<position>-119.5,39</position>
<input>
<ID>ENABLE</ID>1393 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>283 </output>
<output>
<ID>OUT_1</ID>302 </output>
<output>
<ID>OUT_2</ID>245 </output>
<output>
<ID>OUT_3</ID>264 </output>
<output>
<ID>OUT_4</ID>207 </output>
<output>
<ID>OUT_5</ID>226 </output>
<output>
<ID>OUT_6</ID>169 </output>
<output>
<ID>OUT_7</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>460</ID>
<type>AA_AND2</type>
<position>195,-835.5</position>
<input>
<ID>IN_0</ID>423 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>461</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-827</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>425 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>462</ID>
<type>BA_TRI_STATE</type>
<position>283,-835.5</position>
<input>
<ID>ENABLE_0</ID>424 </input>
<input>
<ID>IN_0</ID>425 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_AND2</type>
<position>434,-837</position>
<input>
<ID>IN_0</ID>429 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>AE_DFF_LOW</type>
<position>350,-827</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>427 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>465</ID>
<type>BA_TRI_STATE</type>
<position>374.5,-837</position>
<input>
<ID>ENABLE_0</ID>426 </input>
<input>
<ID>IN_0</ID>427 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>466</ID>
<type>AA_AND2</type>
<position>360,-837</position>
<input>
<ID>IN_0</ID>427 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>426 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>467</ID>
<type>AE_DFF_LOW</type>
<position>423.5,-827</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>429 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>468</ID>
<type>BA_TRI_STATE</type>
<position>448,-837</position>
<input>
<ID>ENABLE_0</ID>428 </input>
<input>
<ID>IN_0</ID>429 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_AND2</type>
<position>592,-839</position>
<input>
<ID>IN_0</ID>433 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>470</ID>
<type>AE_DFF_LOW</type>
<position>508,-827</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>431 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>471</ID>
<type>BA_TRI_STATE</type>
<position>532.5,-839</position>
<input>
<ID>ENABLE_0</ID>430 </input>
<input>
<ID>IN_0</ID>431 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_AND2</type>
<position>518,-839</position>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>473</ID>
<type>AE_DFF_LOW</type>
<position>581.5,-827</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>433 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>474</ID>
<type>BA_TRI_STATE</type>
<position>606,-839</position>
<input>
<ID>ENABLE_0</ID>432 </input>
<input>
<ID>IN_0</ID>433 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_AND2</type>
<position>-4.5,-828</position>
<input>
<ID>IN_0</ID>416 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>476</ID>
<type>BA_TRI_STATE</type>
<position>-26,-847</position>
<input>
<ID>ENABLE_0</ID>416 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>417 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>477</ID>
<type>AA_AND2</type>
<position>118,-1091.5</position>
<input>
<ID>IN_0</ID>440 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>AE_DFF_LOW</type>
<position>34,-1085</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>438 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>479</ID>
<type>BA_TRI_STATE</type>
<position>58.5,-1091.5</position>
<input>
<ID>ENABLE_0</ID>437 </input>
<input>
<ID>IN_0</ID>438 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_AND2</type>
<position>44,-1091.5</position>
<input>
<ID>IN_0</ID>438 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>481</ID>
<type>AE_DFF_LOW</type>
<position>107.5,-1085</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>440 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>482</ID>
<type>BA_TRI_STATE</type>
<position>132,-1091.5</position>
<input>
<ID>ENABLE_0</ID>439 </input>
<input>
<ID>IN_0</ID>440 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>483</ID>
<type>AA_AND2</type>
<position>276,-1093.5</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>443 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>484</ID>
<type>AE_DFF_LOW</type>
<position>192,-1085</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>442 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>485</ID>
<type>BA_TRI_STATE</type>
<position>216.5,-1093.5</position>
<input>
<ID>ENABLE_0</ID>441 </input>
<input>
<ID>IN_0</ID>442 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>486</ID>
<type>AA_AND2</type>
<position>202,-1093.5</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>441 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_DFF_LOW</type>
<position>266.5,-1085</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>444 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>488</ID>
<type>BA_TRI_STATE</type>
<position>290,-1093.5</position>
<input>
<ID>ENABLE_0</ID>443 </input>
<input>
<ID>IN_0</ID>444 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>489</ID>
<type>AA_AND2</type>
<position>441,-1095</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>447 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>490</ID>
<type>AE_DFF_LOW</type>
<position>357,-1085</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>446 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>491</ID>
<type>BA_TRI_STATE</type>
<position>381.5,-1095</position>
<input>
<ID>ENABLE_0</ID>445 </input>
<input>
<ID>IN_0</ID>446 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_AND2</type>
<position>367,-1095</position>
<input>
<ID>IN_0</ID>446 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>493</ID>
<type>AE_DFF_LOW</type>
<position>430.5,-1085</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>448 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>494</ID>
<type>BA_TRI_STATE</type>
<position>455,-1095</position>
<input>
<ID>ENABLE_0</ID>447 </input>
<input>
<ID>IN_0</ID>448 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>495</ID>
<type>AA_AND2</type>
<position>599,-1097</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>496</ID>
<type>AE_DFF_LOW</type>
<position>515,-1085</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>450 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>497</ID>
<type>BA_TRI_STATE</type>
<position>539.5,-1097</position>
<input>
<ID>ENABLE_0</ID>449 </input>
<input>
<ID>IN_0</ID>450 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>498</ID>
<type>AA_AND2</type>
<position>525,-1097</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>499</ID>
<type>AE_DFF_LOW</type>
<position>588.5,-1085</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>452 </output>
<input>
<ID>clock</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>500</ID>
<type>BA_TRI_STATE</type>
<position>613,-1097</position>
<input>
<ID>ENABLE_0</ID>451 </input>
<input>
<ID>IN_0</ID>452 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>501</ID>
<type>AA_AND2</type>
<position>2.5,-1086</position>
<input>
<ID>IN_0</ID>435 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>BA_TRI_STATE</type>
<position>-19,-1105</position>
<input>
<ID>ENABLE_0</ID>435 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>436 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>503</ID>
<type>AA_AND2</type>
<position>115,-1001.5</position>
<input>
<ID>IN_0</ID>459 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>458 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>AE_DFF_LOW</type>
<position>31,-995</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>457 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>505</ID>
<type>BA_TRI_STATE</type>
<position>55.5,-1001.5</position>
<input>
<ID>ENABLE_0</ID>456 </input>
<input>
<ID>IN_0</ID>457 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_AND2</type>
<position>41,-1001.5</position>
<input>
<ID>IN_0</ID>457 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>456 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>507</ID>
<type>AE_DFF_LOW</type>
<position>104.5,-995</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>459 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>508</ID>
<type>BA_TRI_STATE</type>
<position>129,-1001.5</position>
<input>
<ID>ENABLE_0</ID>458 </input>
<input>
<ID>IN_0</ID>459 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_AND2</type>
<position>273,-1003.5</position>
<input>
<ID>IN_0</ID>463 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AE_DFF_LOW</type>
<position>189,-995</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>461 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>511</ID>
<type>BA_TRI_STATE</type>
<position>213.5,-1003.5</position>
<input>
<ID>ENABLE_0</ID>460 </input>
<input>
<ID>IN_0</ID>461 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_AND2</type>
<position>199,-1003.5</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AE_DFF_LOW</type>
<position>263.5,-995</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>463 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>514</ID>
<type>BA_TRI_STATE</type>
<position>287,-1003.5</position>
<input>
<ID>ENABLE_0</ID>462 </input>
<input>
<ID>IN_0</ID>463 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_AND2</type>
<position>438,-1005</position>
<input>
<ID>IN_0</ID>467 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AE_DFF_LOW</type>
<position>354,-995</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>465 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>517</ID>
<type>BA_TRI_STATE</type>
<position>378.5,-1005</position>
<input>
<ID>ENABLE_0</ID>464 </input>
<input>
<ID>IN_0</ID>465 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>518</ID>
<type>AA_AND2</type>
<position>364,-1005</position>
<input>
<ID>IN_0</ID>465 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>464 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>519</ID>
<type>AE_DFF_LOW</type>
<position>427.5,-995</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>467 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>520</ID>
<type>BA_TRI_STATE</type>
<position>452,-1005</position>
<input>
<ID>ENABLE_0</ID>466 </input>
<input>
<ID>IN_0</ID>467 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>521</ID>
<type>AA_AND2</type>
<position>596,-1007</position>
<input>
<ID>IN_0</ID>471 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>470 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>522</ID>
<type>AE_DFF_LOW</type>
<position>512,-995</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>469 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>523</ID>
<type>BA_TRI_STATE</type>
<position>536.5,-1007</position>
<input>
<ID>ENABLE_0</ID>468 </input>
<input>
<ID>IN_0</ID>469 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>524</ID>
<type>AA_AND2</type>
<position>522,-1007</position>
<input>
<ID>IN_0</ID>469 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>525</ID>
<type>AE_DFF_LOW</type>
<position>585.5,-995</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>471 </output>
<input>
<ID>clock</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>526</ID>
<type>BA_TRI_STATE</type>
<position>610,-1007</position>
<input>
<ID>ENABLE_0</ID>470 </input>
<input>
<ID>IN_0</ID>471 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND2</type>
<position>-0.5,-996</position>
<input>
<ID>IN_0</ID>454 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>BA_TRI_STATE</type>
<position>-22,-1015</position>
<input>
<ID>ENABLE_0</ID>454 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>455 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>529</ID>
<type>BE_DECODER_3x8</type>
<position>-119.5,-786.5</position>
<input>
<ID>ENABLE</ID>1394 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>435 </output>
<output>
<ID>OUT_1</ID>454 </output>
<output>
<ID>OUT_2</ID>397 </output>
<output>
<ID>OUT_3</ID>416 </output>
<output>
<ID>OUT_4</ID>359 </output>
<output>
<ID>OUT_5</ID>378 </output>
<output>
<ID>OUT_6</ID>321 </output>
<output>
<ID>OUT_7</ID>340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>530</ID>
<type>AA_AND2</type>
<position>112,-547.5</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>AE_DFF_LOW</type>
<position>28,-541</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>324 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>532</ID>
<type>BA_TRI_STATE</type>
<position>52.5,-547.5</position>
<input>
<ID>ENABLE_0</ID>323 </input>
<input>
<ID>IN_0</ID>324 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>533</ID>
<type>AA_AND2</type>
<position>38,-547.5</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>534</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-541</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>326 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>535</ID>
<type>BA_TRI_STATE</type>
<position>126,-547.5</position>
<input>
<ID>ENABLE_0</ID>325 </input>
<input>
<ID>IN_0</ID>326 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>536</ID>
<type>AA_AND2</type>
<position>270,-549.5</position>
<input>
<ID>IN_0</ID>330 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>537</ID>
<type>AE_DFF_LOW</type>
<position>186,-541</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>328 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>538</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-549.5</position>
<input>
<ID>ENABLE_0</ID>327 </input>
<input>
<ID>IN_0</ID>328 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>539</ID>
<type>AA_AND2</type>
<position>196,-549.5</position>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>327 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>540</ID>
<type>AE_DFF_LOW</type>
<position>260.5,-541</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>330 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>541</ID>
<type>BA_TRI_STATE</type>
<position>284,-549.5</position>
<input>
<ID>ENABLE_0</ID>329 </input>
<input>
<ID>IN_0</ID>330 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>542</ID>
<type>AA_AND2</type>
<position>435,-551</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>333 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>543</ID>
<type>AE_DFF_LOW</type>
<position>351,-541</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>332 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>544</ID>
<type>BA_TRI_STATE</type>
<position>375.5,-551</position>
<input>
<ID>ENABLE_0</ID>331 </input>
<input>
<ID>IN_0</ID>332 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>545</ID>
<type>AA_AND2</type>
<position>361,-551</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>331 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>546</ID>
<type>AE_DFF_LOW</type>
<position>424.5,-541</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>334 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>547</ID>
<type>BA_TRI_STATE</type>
<position>449,-551</position>
<input>
<ID>ENABLE_0</ID>333 </input>
<input>
<ID>IN_0</ID>334 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>548</ID>
<type>AA_AND2</type>
<position>593,-553</position>
<input>
<ID>IN_0</ID>338 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>549</ID>
<type>AE_DFF_LOW</type>
<position>509,-541</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>336 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>550</ID>
<type>BA_TRI_STATE</type>
<position>533.5,-553</position>
<input>
<ID>ENABLE_0</ID>335 </input>
<input>
<ID>IN_0</ID>336 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>551</ID>
<type>AA_AND2</type>
<position>519,-553</position>
<input>
<ID>IN_0</ID>336 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>552</ID>
<type>AE_DFF_LOW</type>
<position>582.5,-541</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>338 </output>
<input>
<ID>clock</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>553</ID>
<type>BA_TRI_STATE</type>
<position>607,-553</position>
<input>
<ID>ENABLE_0</ID>337 </input>
<input>
<ID>IN_0</ID>338 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>554</ID>
<type>AA_AND2</type>
<position>-3.5,-542</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>339 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>BA_TRI_STATE</type>
<position>-25,-561</position>
<input>
<ID>ENABLE_0</ID>321 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>322 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>556</ID>
<type>AA_AND2</type>
<position>109,-457.5</position>
<input>
<ID>IN_0</ID>345 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>344 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>557</ID>
<type>AE_DFF_LOW</type>
<position>25,-451</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>343 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>558</ID>
<type>BA_TRI_STATE</type>
<position>49.5,-457.5</position>
<input>
<ID>ENABLE_0</ID>342 </input>
<input>
<ID>IN_0</ID>343 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>559</ID>
<type>AA_AND2</type>
<position>35,-457.5</position>
<input>
<ID>IN_0</ID>343 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>560</ID>
<type>AE_DFF_LOW</type>
<position>98.5,-451</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>345 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>561</ID>
<type>BA_TRI_STATE</type>
<position>123,-457.5</position>
<input>
<ID>ENABLE_0</ID>344 </input>
<input>
<ID>IN_0</ID>345 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>562</ID>
<type>AA_AND2</type>
<position>267,-459.5</position>
<input>
<ID>IN_0</ID>349 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>348 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>563</ID>
<type>AE_DFF_LOW</type>
<position>183,-451</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>347 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>564</ID>
<type>BA_TRI_STATE</type>
<position>207.5,-459.5</position>
<input>
<ID>ENABLE_0</ID>346 </input>
<input>
<ID>IN_0</ID>347 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_AND2</type>
<position>193,-459.5</position>
<input>
<ID>IN_0</ID>347 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>346 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>566</ID>
<type>AE_DFF_LOW</type>
<position>257.5,-451</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>349 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>567</ID>
<type>BA_TRI_STATE</type>
<position>281,-459.5</position>
<input>
<ID>ENABLE_0</ID>348 </input>
<input>
<ID>IN_0</ID>349 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_AND2</type>
<position>432,-461</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>352 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>569</ID>
<type>AE_DFF_LOW</type>
<position>348,-451</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>351 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>570</ID>
<type>BA_TRI_STATE</type>
<position>372.5,-461</position>
<input>
<ID>ENABLE_0</ID>350 </input>
<input>
<ID>IN_0</ID>351 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>571</ID>
<type>AA_AND2</type>
<position>358,-461</position>
<input>
<ID>IN_0</ID>351 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>AE_DFF_LOW</type>
<position>421.5,-451</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>353 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>573</ID>
<type>BA_TRI_STATE</type>
<position>446,-461</position>
<input>
<ID>ENABLE_0</ID>352 </input>
<input>
<ID>IN_0</ID>353 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>574</ID>
<type>AA_AND2</type>
<position>590,-463</position>
<input>
<ID>IN_0</ID>357 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>356 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>575</ID>
<type>AE_DFF_LOW</type>
<position>506,-451</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>355 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>576</ID>
<type>BA_TRI_STATE</type>
<position>530.5,-463</position>
<input>
<ID>ENABLE_0</ID>354 </input>
<input>
<ID>IN_0</ID>355 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>577</ID>
<type>AA_AND2</type>
<position>516,-463</position>
<input>
<ID>IN_0</ID>355 </input>
<input>
<ID>IN_1</ID>341 </input>
<output>
<ID>OUT</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>AE_DFF_LOW</type>
<position>579.5,-451</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>357 </output>
<input>
<ID>clock</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>579</ID>
<type>BA_TRI_STATE</type>
<position>604,-463</position>
<input>
<ID>ENABLE_0</ID>356 </input>
<input>
<ID>IN_0</ID>357 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>580</ID>
<type>AA_AND2</type>
<position>-6.5,-452</position>
<input>
<ID>IN_0</ID>340 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>581</ID>
<type>BA_TRI_STATE</type>
<position>-28,-471</position>
<input>
<ID>ENABLE_0</ID>340 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>341 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>582</ID>
<type>AA_AND2</type>
<position>116,-715.5</position>
<input>
<ID>IN_0</ID>364 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>583</ID>
<type>AE_DFF_LOW</type>
<position>32,-709</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>362 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>584</ID>
<type>BA_TRI_STATE</type>
<position>56.5,-715.5</position>
<input>
<ID>ENABLE_0</ID>361 </input>
<input>
<ID>IN_0</ID>362 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_AND2</type>
<position>42,-715.5</position>
<input>
<ID>IN_0</ID>362 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>361 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>586</ID>
<type>AE_DFF_LOW</type>
<position>105.5,-709</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>364 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>587</ID>
<type>BA_TRI_STATE</type>
<position>130,-715.5</position>
<input>
<ID>ENABLE_0</ID>363 </input>
<input>
<ID>IN_0</ID>364 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>588</ID>
<type>AA_AND2</type>
<position>274,-717.5</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>589</ID>
<type>AE_DFF_LOW</type>
<position>190,-709</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>366 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>590</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-717.5</position>
<input>
<ID>ENABLE_0</ID>365 </input>
<input>
<ID>IN_0</ID>366 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>591</ID>
<type>AA_AND2</type>
<position>200,-717.5</position>
<input>
<ID>IN_0</ID>366 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>592</ID>
<type>AE_DFF_LOW</type>
<position>264.5,-709</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>368 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>593</ID>
<type>BA_TRI_STATE</type>
<position>288,-717.5</position>
<input>
<ID>ENABLE_0</ID>367 </input>
<input>
<ID>IN_0</ID>368 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>594</ID>
<type>AA_AND2</type>
<position>439,-719</position>
<input>
<ID>IN_0</ID>372 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>371 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>595</ID>
<type>AE_DFF_LOW</type>
<position>355,-709</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>370 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>596</ID>
<type>BA_TRI_STATE</type>
<position>379.5,-719</position>
<input>
<ID>ENABLE_0</ID>369 </input>
<input>
<ID>IN_0</ID>370 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>597</ID>
<type>AA_AND2</type>
<position>365,-719</position>
<input>
<ID>IN_0</ID>370 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>369 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>AE_DFF_LOW</type>
<position>428.5,-709</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>372 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>599</ID>
<type>BA_TRI_STATE</type>
<position>453,-719</position>
<input>
<ID>ENABLE_0</ID>371 </input>
<input>
<ID>IN_0</ID>372 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_AND2</type>
<position>597,-721</position>
<input>
<ID>IN_0</ID>376 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>375 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AE_DFF_LOW</type>
<position>513,-709</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>374 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>602</ID>
<type>BA_TRI_STATE</type>
<position>537.5,-721</position>
<input>
<ID>ENABLE_0</ID>373 </input>
<input>
<ID>IN_0</ID>374 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_AND2</type>
<position>523,-721</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>373 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>604</ID>
<type>AE_DFF_LOW</type>
<position>586.5,-709</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>376 </output>
<input>
<ID>clock</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>605</ID>
<type>BA_TRI_STATE</type>
<position>611,-721</position>
<input>
<ID>ENABLE_0</ID>375 </input>
<input>
<ID>IN_0</ID>376 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>606</ID>
<type>AA_AND2</type>
<position>0.5,-710</position>
<input>
<ID>IN_0</ID>359 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>377 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>607</ID>
<type>BA_TRI_STATE</type>
<position>-21,-729</position>
<input>
<ID>ENABLE_0</ID>359 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>360 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_AND2</type>
<position>113,-625.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>609</ID>
<type>AE_DFF_LOW</type>
<position>29,-619</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>381 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>610</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-625.5</position>
<input>
<ID>ENABLE_0</ID>380 </input>
<input>
<ID>IN_0</ID>381 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>611</ID>
<type>AA_AND2</type>
<position>39,-625.5</position>
<input>
<ID>IN_0</ID>381 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>612</ID>
<type>AE_DFF_LOW</type>
<position>102.5,-619</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>383 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>613</ID>
<type>BA_TRI_STATE</type>
<position>127,-625.5</position>
<input>
<ID>ENABLE_0</ID>382 </input>
<input>
<ID>IN_0</ID>383 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>614</ID>
<type>AA_AND2</type>
<position>271,-627.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AE_DFF_LOW</type>
<position>187,-619</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>385 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>616</ID>
<type>BA_TRI_STATE</type>
<position>211.5,-627.5</position>
<input>
<ID>ENABLE_0</ID>384 </input>
<input>
<ID>IN_0</ID>385 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>617</ID>
<type>AA_AND2</type>
<position>197,-627.5</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>384 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>AE_DFF_LOW</type>
<position>261.5,-619</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>387 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>619</ID>
<type>BA_TRI_STATE</type>
<position>285,-627.5</position>
<input>
<ID>ENABLE_0</ID>386 </input>
<input>
<ID>IN_0</ID>387 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>620</ID>
<type>AA_AND2</type>
<position>436,-629</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>390 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>621</ID>
<type>AE_DFF_LOW</type>
<position>352,-619</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>389 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>622</ID>
<type>BA_TRI_STATE</type>
<position>376.5,-629</position>
<input>
<ID>ENABLE_0</ID>388 </input>
<input>
<ID>IN_0</ID>389 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>623</ID>
<type>AA_AND2</type>
<position>362,-629</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>388 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>624</ID>
<type>AE_DFF_LOW</type>
<position>425.5,-619</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>391 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>625</ID>
<type>BA_TRI_STATE</type>
<position>450,-629</position>
<input>
<ID>ENABLE_0</ID>390 </input>
<input>
<ID>IN_0</ID>391 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>626</ID>
<type>AA_AND2</type>
<position>594,-631</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>627</ID>
<type>AE_DFF_LOW</type>
<position>510,-619</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>393 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>628</ID>
<type>BA_TRI_STATE</type>
<position>534.5,-631</position>
<input>
<ID>ENABLE_0</ID>392 </input>
<input>
<ID>IN_0</ID>393 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>629</ID>
<type>AA_AND2</type>
<position>520,-631</position>
<input>
<ID>IN_0</ID>393 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>630</ID>
<type>AE_DFF_LOW</type>
<position>583.5,-619</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>395 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>631</ID>
<type>BA_TRI_STATE</type>
<position>608,-631</position>
<input>
<ID>ENABLE_0</ID>394 </input>
<input>
<ID>IN_0</ID>395 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>632</ID>
<type>AA_AND2</type>
<position>-2.5,-620</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>633</ID>
<type>BA_TRI_STATE</type>
<position>-24,-639</position>
<input>
<ID>ENABLE_0</ID>378 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>379 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>634</ID>
<type>AA_AND2</type>
<position>114,-923.5</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>635</ID>
<type>AE_DFF_LOW</type>
<position>30,-917</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>400 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>636</ID>
<type>BA_TRI_STATE</type>
<position>54.5,-923.5</position>
<input>
<ID>ENABLE_0</ID>399 </input>
<input>
<ID>IN_0</ID>400 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>637</ID>
<type>AA_AND2</type>
<position>40,-923.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>638</ID>
<type>AE_DFF_LOW</type>
<position>103.5,-917</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>402 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>639</ID>
<type>BA_TRI_STATE</type>
<position>129,-923.5</position>
<input>
<ID>ENABLE_0</ID>401 </input>
<input>
<ID>IN_0</ID>402 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>640</ID>
<type>AA_AND2</type>
<position>272,-925.5</position>
<input>
<ID>IN_0</ID>406 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>405 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_DFF_LOW</type>
<position>188,-917</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>404 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>642</ID>
<type>BA_TRI_STATE</type>
<position>212.5,-925.5</position>
<input>
<ID>ENABLE_0</ID>403 </input>
<input>
<ID>IN_0</ID>404 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>643</ID>
<type>AA_AND2</type>
<position>198,-925.5</position>
<input>
<ID>IN_0</ID>404 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>403 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>644</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-917</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>406 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>645</ID>
<type>BA_TRI_STATE</type>
<position>286,-925.5</position>
<input>
<ID>ENABLE_0</ID>405 </input>
<input>
<ID>IN_0</ID>406 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>646</ID>
<type>AA_AND2</type>
<position>437,-927</position>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>647</ID>
<type>AE_DFF_LOW</type>
<position>353,-917</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>408 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>648</ID>
<type>BA_TRI_STATE</type>
<position>377.5,-927</position>
<input>
<ID>ENABLE_0</ID>407 </input>
<input>
<ID>IN_0</ID>408 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>649</ID>
<type>AA_AND2</type>
<position>363,-927</position>
<input>
<ID>IN_0</ID>408 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>407 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>650</ID>
<type>AE_DFF_LOW</type>
<position>426.5,-917</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>410 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>651</ID>
<type>BA_TRI_STATE</type>
<position>451,-927</position>
<input>
<ID>ENABLE_0</ID>409 </input>
<input>
<ID>IN_0</ID>410 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>652</ID>
<type>AA_AND2</type>
<position>595,-929</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>653</ID>
<type>AE_DFF_LOW</type>
<position>511,-917</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>412 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>654</ID>
<type>BA_TRI_STATE</type>
<position>535.5,-929</position>
<input>
<ID>ENABLE_0</ID>411 </input>
<input>
<ID>IN_0</ID>412 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>655</ID>
<type>AA_AND2</type>
<position>521,-929</position>
<input>
<ID>IN_0</ID>412 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>656</ID>
<type>AE_DFF_LOW</type>
<position>584.5,-917</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>414 </output>
<input>
<ID>clock</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>657</ID>
<type>BA_TRI_STATE</type>
<position>609,-929</position>
<input>
<ID>ENABLE_0</ID>413 </input>
<input>
<ID>IN_0</ID>414 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>658</ID>
<type>AA_AND2</type>
<position>-1.5,-918</position>
<input>
<ID>IN_0</ID>397 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>659</ID>
<type>BA_TRI_STATE</type>
<position>-23,-937</position>
<input>
<ID>ENABLE_0</ID>397 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>398 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>660</ID>
<type>AA_AND2</type>
<position>111,-833.5</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>661</ID>
<type>AE_DFF_LOW</type>
<position>27,-827</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>419 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>662</ID>
<type>BA_TRI_STATE</type>
<position>51.5,-833.5</position>
<input>
<ID>ENABLE_0</ID>418 </input>
<input>
<ID>IN_0</ID>419 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>663</ID>
<type>AA_AND2</type>
<position>37,-833.5</position>
<input>
<ID>IN_0</ID>419 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>664</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-827</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>421 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>665</ID>
<type>BA_TRI_STATE</type>
<position>125,-833.5</position>
<input>
<ID>ENABLE_0</ID>420 </input>
<input>
<ID>IN_0</ID>421 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>666</ID>
<type>AA_AND2</type>
<position>269,-835.5</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>667</ID>
<type>AE_DFF_LOW</type>
<position>185,-827</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>423 </output>
<input>
<ID>clock</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>668</ID>
<type>BA_TRI_STATE</type>
<position>209.5,-835.5</position>
<input>
<ID>ENABLE_0</ID>422 </input>
<input>
<ID>IN_0</ID>423 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>669</ID>
<type>AA_AND2</type>
<position>192.5,-1760</position>
<input>
<ID>IN_0</ID>575 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>574 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>AE_DFF_LOW</type>
<position>257,-1751.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>577 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>671</ID>
<type>BA_TRI_STATE</type>
<position>280.5,-1760</position>
<input>
<ID>ENABLE_0</ID>576 </input>
<input>
<ID>IN_0</ID>577 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>672</ID>
<type>AA_AND2</type>
<position>431.5,-1761.5</position>
<input>
<ID>IN_0</ID>581 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>673</ID>
<type>AE_DFF_LOW</type>
<position>347.5,-1751.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>579 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>674</ID>
<type>BA_TRI_STATE</type>
<position>372,-1761.5</position>
<input>
<ID>ENABLE_0</ID>578 </input>
<input>
<ID>IN_0</ID>579 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_AND2</type>
<position>357.5,-1761.5</position>
<input>
<ID>IN_0</ID>579 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>578 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>676</ID>
<type>AE_DFF_LOW</type>
<position>421,-1751.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>581 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>677</ID>
<type>BA_TRI_STATE</type>
<position>445.5,-1761.5</position>
<input>
<ID>ENABLE_0</ID>580 </input>
<input>
<ID>IN_0</ID>581 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>678</ID>
<type>AA_AND2</type>
<position>589.5,-1763.5</position>
<input>
<ID>IN_0</ID>585 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>679</ID>
<type>AE_DFF_LOW</type>
<position>505.5,-1751.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>583 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>680</ID>
<type>BA_TRI_STATE</type>
<position>530,-1763.5</position>
<input>
<ID>ENABLE_0</ID>582 </input>
<input>
<ID>IN_0</ID>583 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>681</ID>
<type>AA_AND2</type>
<position>515.5,-1763.5</position>
<input>
<ID>IN_0</ID>583 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>582 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>682</ID>
<type>AE_DFF_LOW</type>
<position>579,-1751.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>585 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>683</ID>
<type>BA_TRI_STATE</type>
<position>603.5,-1763.5</position>
<input>
<ID>ENABLE_0</ID>584 </input>
<input>
<ID>IN_0</ID>585 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>684</ID>
<type>AA_AND2</type>
<position>-7,-1752.5</position>
<input>
<ID>IN_0</ID>568 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>685</ID>
<type>BA_TRI_STATE</type>
<position>-28.5,-1771.5</position>
<input>
<ID>ENABLE_0</ID>568 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>569 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>686</ID>
<type>AA_AND2</type>
<position>115.5,-2016</position>
<input>
<ID>IN_0</ID>592 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_DFF_LOW</type>
<position>31.5,-2009.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>590 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>688</ID>
<type>BA_TRI_STATE</type>
<position>56,-2016</position>
<input>
<ID>ENABLE_0</ID>589 </input>
<input>
<ID>IN_0</ID>590 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>689</ID>
<type>AA_AND2</type>
<position>41.5,-2016</position>
<input>
<ID>IN_0</ID>590 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>589 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_DFF_LOW</type>
<position>105,-2009.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>592 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>691</ID>
<type>BA_TRI_STATE</type>
<position>129.5,-2016</position>
<input>
<ID>ENABLE_0</ID>591 </input>
<input>
<ID>IN_0</ID>592 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>692</ID>
<type>AA_AND2</type>
<position>273.5,-2018</position>
<input>
<ID>IN_0</ID>596 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>693</ID>
<type>AE_DFF_LOW</type>
<position>189.5,-2009.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>594 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>694</ID>
<type>BA_TRI_STATE</type>
<position>214,-2018</position>
<input>
<ID>ENABLE_0</ID>593 </input>
<input>
<ID>IN_0</ID>594 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>695</ID>
<type>AA_AND2</type>
<position>199.5,-2018</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>696</ID>
<type>AE_DFF_LOW</type>
<position>264,-2009.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>596 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>697</ID>
<type>BA_TRI_STATE</type>
<position>287.5,-2018</position>
<input>
<ID>ENABLE_0</ID>595 </input>
<input>
<ID>IN_0</ID>596 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>698</ID>
<type>AA_AND2</type>
<position>438.5,-2019.5</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>699</ID>
<type>AE_DFF_LOW</type>
<position>354.5,-2009.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>598 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>700</ID>
<type>BA_TRI_STATE</type>
<position>379,-2019.5</position>
<input>
<ID>ENABLE_0</ID>597 </input>
<input>
<ID>IN_0</ID>598 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_AND2</type>
<position>364.5,-2019.5</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>702</ID>
<type>AE_DFF_LOW</type>
<position>428,-2009.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>600 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>703</ID>
<type>BA_TRI_STATE</type>
<position>452.5,-2019.5</position>
<input>
<ID>ENABLE_0</ID>599 </input>
<input>
<ID>IN_0</ID>600 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>704</ID>
<type>AA_AND2</type>
<position>596.5,-2021.5</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>603 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>705</ID>
<type>AE_DFF_LOW</type>
<position>512.5,-2009.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>602 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>706</ID>
<type>BA_TRI_STATE</type>
<position>537,-2021.5</position>
<input>
<ID>ENABLE_0</ID>601 </input>
<input>
<ID>IN_0</ID>602 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>707</ID>
<type>AA_AND2</type>
<position>522.5,-2021.5</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>588 </input>
<output>
<ID>OUT</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>708</ID>
<type>AE_DFF_LOW</type>
<position>586,-2009.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>604 </output>
<input>
<ID>clock</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>709</ID>
<type>BA_TRI_STATE</type>
<position>610.5,-2021.5</position>
<input>
<ID>ENABLE_0</ID>603 </input>
<input>
<ID>IN_0</ID>604 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>710</ID>
<type>AA_AND2</type>
<position>0,-2010.5</position>
<input>
<ID>IN_0</ID>587 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>605 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>711</ID>
<type>BA_TRI_STATE</type>
<position>-21.5,-2029.5</position>
<input>
<ID>ENABLE_0</ID>587 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>588 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>712</ID>
<type>AA_AND2</type>
<position>112.5,-1926</position>
<input>
<ID>IN_0</ID>611 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>610 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>713</ID>
<type>AE_DFF_LOW</type>
<position>28.5,-1919.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>609 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>714</ID>
<type>BA_TRI_STATE</type>
<position>53,-1926</position>
<input>
<ID>ENABLE_0</ID>608 </input>
<input>
<ID>IN_0</ID>609 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>715</ID>
<type>AA_AND2</type>
<position>38.5,-1926</position>
<input>
<ID>IN_0</ID>609 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>716</ID>
<type>AE_DFF_LOW</type>
<position>102,-1919.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>611 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>717</ID>
<type>BA_TRI_STATE</type>
<position>126.5,-1926</position>
<input>
<ID>ENABLE_0</ID>610 </input>
<input>
<ID>IN_0</ID>611 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>718</ID>
<type>AA_AND2</type>
<position>270.5,-1928</position>
<input>
<ID>IN_0</ID>615 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>614 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>719</ID>
<type>AE_DFF_LOW</type>
<position>186.5,-1919.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>613 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>720</ID>
<type>BA_TRI_STATE</type>
<position>211,-1928</position>
<input>
<ID>ENABLE_0</ID>612 </input>
<input>
<ID>IN_0</ID>613 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>721</ID>
<type>AA_AND2</type>
<position>196.5,-1928</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>722</ID>
<type>AE_DFF_LOW</type>
<position>261,-1919.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>615 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>723</ID>
<type>BA_TRI_STATE</type>
<position>284.5,-1928</position>
<input>
<ID>ENABLE_0</ID>614 </input>
<input>
<ID>IN_0</ID>615 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>724</ID>
<type>AA_AND2</type>
<position>435.5,-1929.5</position>
<input>
<ID>IN_0</ID>619 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>618 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>725</ID>
<type>AE_DFF_LOW</type>
<position>351.5,-1919.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>617 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>726</ID>
<type>BA_TRI_STATE</type>
<position>376,-1929.5</position>
<input>
<ID>ENABLE_0</ID>616 </input>
<input>
<ID>IN_0</ID>617 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>727</ID>
<type>AA_AND2</type>
<position>361.5,-1929.5</position>
<input>
<ID>IN_0</ID>617 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>616 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>728</ID>
<type>AE_DFF_LOW</type>
<position>425,-1919.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>619 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>729</ID>
<type>BA_TRI_STATE</type>
<position>449.5,-1929.5</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>619 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>730</ID>
<type>AA_AND2</type>
<position>593.5,-1931.5</position>
<input>
<ID>IN_0</ID>623 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>622 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>731</ID>
<type>AE_DFF_LOW</type>
<position>509.5,-1919.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>621 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>732</ID>
<type>BA_TRI_STATE</type>
<position>534,-1931.5</position>
<input>
<ID>ENABLE_0</ID>620 </input>
<input>
<ID>IN_0</ID>621 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>733</ID>
<type>AA_AND2</type>
<position>519.5,-1931.5</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>620 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>734</ID>
<type>AE_DFF_LOW</type>
<position>583,-1919.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>623 </output>
<input>
<ID>clock</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>735</ID>
<type>BA_TRI_STATE</type>
<position>607.5,-1931.5</position>
<input>
<ID>ENABLE_0</ID>622 </input>
<input>
<ID>IN_0</ID>623 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>736</ID>
<type>AA_AND2</type>
<position>-3,-1920.5</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>624 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>737</ID>
<type>BA_TRI_STATE</type>
<position>-24.5,-1939.5</position>
<input>
<ID>ENABLE_0</ID>606 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>607 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>738</ID>
<type>BE_DECODER_3x8</type>
<position>-122,-1711</position>
<input>
<ID>ENABLE</ID>1395 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>587 </output>
<output>
<ID>OUT_1</ID>606 </output>
<output>
<ID>OUT_2</ID>549 </output>
<output>
<ID>OUT_3</ID>568 </output>
<output>
<ID>OUT_4</ID>511 </output>
<output>
<ID>OUT_5</ID>530 </output>
<output>
<ID>OUT_6</ID>473 </output>
<output>
<ID>OUT_7</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>739</ID>
<type>AA_AND2</type>
<position>109.5,-1472</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>477 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>740</ID>
<type>AE_DFF_LOW</type>
<position>25.5,-1465.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>476 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>741</ID>
<type>BA_TRI_STATE</type>
<position>50,-1472</position>
<input>
<ID>ENABLE_0</ID>475 </input>
<input>
<ID>IN_0</ID>476 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>742</ID>
<type>AA_AND2</type>
<position>35.5,-1472</position>
<input>
<ID>IN_0</ID>476 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>475 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>743</ID>
<type>AE_DFF_LOW</type>
<position>99,-1465.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>478 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>744</ID>
<type>BA_TRI_STATE</type>
<position>123.5,-1472</position>
<input>
<ID>ENABLE_0</ID>477 </input>
<input>
<ID>IN_0</ID>478 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>745</ID>
<type>AA_AND2</type>
<position>267.5,-1474</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>746</ID>
<type>AE_DFF_LOW</type>
<position>183.5,-1465.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>480 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>747</ID>
<type>BA_TRI_STATE</type>
<position>208,-1474</position>
<input>
<ID>ENABLE_0</ID>479 </input>
<input>
<ID>IN_0</ID>480 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>748</ID>
<type>AA_AND2</type>
<position>193.5,-1474</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>749</ID>
<type>AE_DFF_LOW</type>
<position>258,-1465.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>482 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>750</ID>
<type>BA_TRI_STATE</type>
<position>281.5,-1474</position>
<input>
<ID>ENABLE_0</ID>481 </input>
<input>
<ID>IN_0</ID>482 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>751</ID>
<type>AA_AND2</type>
<position>432.5,-1475.5</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>752</ID>
<type>AE_DFF_LOW</type>
<position>348.5,-1465.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>484 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>753</ID>
<type>BA_TRI_STATE</type>
<position>373,-1475.5</position>
<input>
<ID>ENABLE_0</ID>483 </input>
<input>
<ID>IN_0</ID>484 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>754</ID>
<type>AA_AND2</type>
<position>358.5,-1475.5</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>755</ID>
<type>AE_DFF_LOW</type>
<position>422,-1465.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>486 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>756</ID>
<type>BA_TRI_STATE</type>
<position>446.5,-1475.5</position>
<input>
<ID>ENABLE_0</ID>485 </input>
<input>
<ID>IN_0</ID>486 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>757</ID>
<type>AA_AND2</type>
<position>590.5,-1477.5</position>
<input>
<ID>IN_0</ID>490 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>489 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>758</ID>
<type>AE_DFF_LOW</type>
<position>506.5,-1465.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>488 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>759</ID>
<type>BA_TRI_STATE</type>
<position>531,-1477.5</position>
<input>
<ID>ENABLE_0</ID>487 </input>
<input>
<ID>IN_0</ID>488 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>760</ID>
<type>AA_AND2</type>
<position>516.5,-1477.5</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>AE_DFF_LOW</type>
<position>580,-1465.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>490 </output>
<input>
<ID>clock</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>762</ID>
<type>BA_TRI_STATE</type>
<position>604.5,-1477.5</position>
<input>
<ID>ENABLE_0</ID>489 </input>
<input>
<ID>IN_0</ID>490 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>763</ID>
<type>AA_AND2</type>
<position>-6,-1466.5</position>
<input>
<ID>IN_0</ID>473 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>491 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>764</ID>
<type>BA_TRI_STATE</type>
<position>-27.5,-1485.5</position>
<input>
<ID>ENABLE_0</ID>473 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>474 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_AND2</type>
<position>106.5,-1382</position>
<input>
<ID>IN_0</ID>497 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>766</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-1375.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>495 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>767</ID>
<type>BA_TRI_STATE</type>
<position>47,-1382</position>
<input>
<ID>ENABLE_0</ID>494 </input>
<input>
<ID>IN_0</ID>495 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>768</ID>
<type>AA_AND2</type>
<position>32.5,-1382</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>769</ID>
<type>AE_DFF_LOW</type>
<position>96,-1375.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>497 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>770</ID>
<type>BA_TRI_STATE</type>
<position>120.5,-1382</position>
<input>
<ID>ENABLE_0</ID>496 </input>
<input>
<ID>IN_0</ID>497 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>771</ID>
<type>AA_AND2</type>
<position>264.5,-1384</position>
<input>
<ID>IN_0</ID>501 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>500 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>772</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-1375.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>499 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>773</ID>
<type>BA_TRI_STATE</type>
<position>205,-1384</position>
<input>
<ID>ENABLE_0</ID>498 </input>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>774</ID>
<type>AA_AND2</type>
<position>190.5,-1384</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>498 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>775</ID>
<type>AE_DFF_LOW</type>
<position>255,-1375.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>501 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>776</ID>
<type>BA_TRI_STATE</type>
<position>278.5,-1384</position>
<input>
<ID>ENABLE_0</ID>500 </input>
<input>
<ID>IN_0</ID>501 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_AND2</type>
<position>429.5,-1385.5</position>
<input>
<ID>IN_0</ID>505 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>778</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-1375.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>503 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>779</ID>
<type>BA_TRI_STATE</type>
<position>370,-1385.5</position>
<input>
<ID>ENABLE_0</ID>502 </input>
<input>
<ID>IN_0</ID>503 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>780</ID>
<type>AA_AND2</type>
<position>355.5,-1385.5</position>
<input>
<ID>IN_0</ID>503 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>502 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>781</ID>
<type>AE_DFF_LOW</type>
<position>419,-1375.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>505 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>782</ID>
<type>BA_TRI_STATE</type>
<position>443.5,-1385.5</position>
<input>
<ID>ENABLE_0</ID>504 </input>
<input>
<ID>IN_0</ID>505 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>783</ID>
<type>AA_AND2</type>
<position>587.5,-1387.5</position>
<input>
<ID>IN_0</ID>509 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AE_DFF_LOW</type>
<position>503.5,-1375.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>507 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>785</ID>
<type>BA_TRI_STATE</type>
<position>528,-1387.5</position>
<input>
<ID>ENABLE_0</ID>506 </input>
<input>
<ID>IN_0</ID>507 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>786</ID>
<type>AA_AND2</type>
<position>513.5,-1387.5</position>
<input>
<ID>IN_0</ID>507 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>787</ID>
<type>AE_DFF_LOW</type>
<position>577,-1375.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>509 </output>
<input>
<ID>clock</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>788</ID>
<type>BA_TRI_STATE</type>
<position>601.5,-1387.5</position>
<input>
<ID>ENABLE_0</ID>508 </input>
<input>
<ID>IN_0</ID>509 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>789</ID>
<type>AA_AND2</type>
<position>-9,-1376.5</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>790</ID>
<type>BA_TRI_STATE</type>
<position>-26,-1396</position>
<input>
<ID>ENABLE_0</ID>492 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>493 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>791</ID>
<type>AA_AND2</type>
<position>113.5,-1640</position>
<input>
<ID>IN_0</ID>516 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>515 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>792</ID>
<type>AE_DFF_LOW</type>
<position>29.5,-1633.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>514 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>793</ID>
<type>BA_TRI_STATE</type>
<position>54,-1640</position>
<input>
<ID>ENABLE_0</ID>513 </input>
<input>
<ID>IN_0</ID>514 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>794</ID>
<type>AA_AND2</type>
<position>39.5,-1640</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>795</ID>
<type>AE_DFF_LOW</type>
<position>103,-1633.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>516 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>796</ID>
<type>BA_TRI_STATE</type>
<position>127.5,-1640</position>
<input>
<ID>ENABLE_0</ID>515 </input>
<input>
<ID>IN_0</ID>516 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>797</ID>
<type>AA_AND2</type>
<position>271.5,-1642</position>
<input>
<ID>IN_0</ID>520 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>519 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>798</ID>
<type>AE_DFF_LOW</type>
<position>187.5,-1633.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>518 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>799</ID>
<type>BA_TRI_STATE</type>
<position>212,-1642</position>
<input>
<ID>ENABLE_0</ID>517 </input>
<input>
<ID>IN_0</ID>518 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_AND2</type>
<position>197.5,-1642</position>
<input>
<ID>IN_0</ID>518 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>801</ID>
<type>AE_DFF_LOW</type>
<position>262,-1633.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>520 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>802</ID>
<type>BA_TRI_STATE</type>
<position>285.5,-1642</position>
<input>
<ID>ENABLE_0</ID>519 </input>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>803</ID>
<type>AA_AND2</type>
<position>436.5,-1643.5</position>
<input>
<ID>IN_0</ID>524 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>804</ID>
<type>AE_DFF_LOW</type>
<position>352.5,-1633.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>522 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>805</ID>
<type>BA_TRI_STATE</type>
<position>377,-1643.5</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>806</ID>
<type>AA_AND2</type>
<position>362.5,-1643.5</position>
<input>
<ID>IN_0</ID>522 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>521 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>807</ID>
<type>AE_DFF_LOW</type>
<position>426,-1633.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>524 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>808</ID>
<type>BA_TRI_STATE</type>
<position>450.5,-1643.5</position>
<input>
<ID>ENABLE_0</ID>523 </input>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>809</ID>
<type>AA_AND2</type>
<position>594.5,-1645.5</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>527 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>810</ID>
<type>AE_DFF_LOW</type>
<position>510.5,-1633.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>526 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>811</ID>
<type>BA_TRI_STATE</type>
<position>535,-1645.5</position>
<input>
<ID>ENABLE_0</ID>525 </input>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>812</ID>
<type>AA_AND2</type>
<position>520.5,-1645.5</position>
<input>
<ID>IN_0</ID>526 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>813</ID>
<type>AE_DFF_LOW</type>
<position>584,-1633.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>528 </output>
<input>
<ID>clock</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>814</ID>
<type>BA_TRI_STATE</type>
<position>608.5,-1645.5</position>
<input>
<ID>ENABLE_0</ID>527 </input>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>815</ID>
<type>AA_AND2</type>
<position>-2,-1634.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>1456 </input>
<output>
<ID>OUT</ID>529 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>816</ID>
<type>BA_TRI_STATE</type>
<position>-23.5,-1653.5</position>
<input>
<ID>ENABLE_0</ID>511 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>512 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>817</ID>
<type>AA_AND2</type>
<position>110.5,-1550</position>
<input>
<ID>IN_0</ID>535 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>534 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>818</ID>
<type>AE_DFF_LOW</type>
<position>26.5,-1543.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>533 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>819</ID>
<type>BA_TRI_STATE</type>
<position>51,-1550</position>
<input>
<ID>ENABLE_0</ID>532 </input>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>820</ID>
<type>AA_AND2</type>
<position>36.5,-1550</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>821</ID>
<type>AE_DFF_LOW</type>
<position>100,-1543.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>535 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>822</ID>
<type>BA_TRI_STATE</type>
<position>124.5,-1550</position>
<input>
<ID>ENABLE_0</ID>534 </input>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>823</ID>
<type>AA_AND2</type>
<position>268.5,-1552</position>
<input>
<ID>IN_0</ID>539 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>538 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>824</ID>
<type>AE_DFF_LOW</type>
<position>184.5,-1543.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>537 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>825</ID>
<type>BA_TRI_STATE</type>
<position>209,-1552</position>
<input>
<ID>ENABLE_0</ID>536 </input>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>826</ID>
<type>AA_AND2</type>
<position>194.5,-1552</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>536 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>827</ID>
<type>AE_DFF_LOW</type>
<position>259,-1543.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>539 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>828</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-1552</position>
<input>
<ID>ENABLE_0</ID>538 </input>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>829</ID>
<type>AA_AND2</type>
<position>433.5,-1553.5</position>
<input>
<ID>IN_0</ID>543 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>542 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>830</ID>
<type>AE_DFF_LOW</type>
<position>349.5,-1543.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>541 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>831</ID>
<type>BA_TRI_STATE</type>
<position>374,-1553.5</position>
<input>
<ID>ENABLE_0</ID>540 </input>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>832</ID>
<type>AA_AND2</type>
<position>359.5,-1553.5</position>
<input>
<ID>IN_0</ID>541 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>540 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>833</ID>
<type>AE_DFF_LOW</type>
<position>423,-1543.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>543 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>834</ID>
<type>BA_TRI_STATE</type>
<position>447.5,-1553.5</position>
<input>
<ID>ENABLE_0</ID>542 </input>
<input>
<ID>IN_0</ID>543 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>835</ID>
<type>AA_AND2</type>
<position>591.5,-1555.5</position>
<input>
<ID>IN_0</ID>547 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>836</ID>
<type>AE_DFF_LOW</type>
<position>507.5,-1543.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>545 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>837</ID>
<type>BA_TRI_STATE</type>
<position>532,-1555.5</position>
<input>
<ID>ENABLE_0</ID>544 </input>
<input>
<ID>IN_0</ID>545 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>838</ID>
<type>AA_AND2</type>
<position>517.5,-1555.5</position>
<input>
<ID>IN_0</ID>545 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>544 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>839</ID>
<type>AE_DFF_LOW</type>
<position>581,-1543.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>547 </output>
<input>
<ID>clock</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>840</ID>
<type>BA_TRI_STATE</type>
<position>605.5,-1555.5</position>
<input>
<ID>ENABLE_0</ID>546 </input>
<input>
<ID>IN_0</ID>547 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>841</ID>
<type>AA_AND2</type>
<position>-5,-1544.5</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>548 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>842</ID>
<type>BA_TRI_STATE</type>
<position>-26.5,-1563.5</position>
<input>
<ID>ENABLE_0</ID>530 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>531 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>843</ID>
<type>AA_AND2</type>
<position>111.5,-1848</position>
<input>
<ID>IN_0</ID>554 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>844</ID>
<type>AE_DFF_LOW</type>
<position>27.5,-1841.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>552 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>845</ID>
<type>BA_TRI_STATE</type>
<position>52,-1848</position>
<input>
<ID>ENABLE_0</ID>551 </input>
<input>
<ID>IN_0</ID>552 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>846</ID>
<type>AA_AND2</type>
<position>37.5,-1848</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>551 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>847</ID>
<type>AE_DFF_LOW</type>
<position>101,-1841.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>554 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>848</ID>
<type>BA_TRI_STATE</type>
<position>125.5,-1848</position>
<input>
<ID>ENABLE_0</ID>553 </input>
<input>
<ID>IN_0</ID>554 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>849</ID>
<type>AA_AND2</type>
<position>269.5,-1850</position>
<input>
<ID>IN_0</ID>558 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>557 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>850</ID>
<type>AE_DFF_LOW</type>
<position>185.5,-1841.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>556 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>851</ID>
<type>BA_TRI_STATE</type>
<position>210,-1850</position>
<input>
<ID>ENABLE_0</ID>555 </input>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>852</ID>
<type>AA_AND2</type>
<position>195.5,-1850</position>
<input>
<ID>IN_0</ID>556 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>853</ID>
<type>AE_DFF_LOW</type>
<position>260,-1841.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>558 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>854</ID>
<type>BA_TRI_STATE</type>
<position>283.5,-1850</position>
<input>
<ID>ENABLE_0</ID>557 </input>
<input>
<ID>IN_0</ID>558 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>855</ID>
<type>AA_AND2</type>
<position>434.5,-1851.5</position>
<input>
<ID>IN_0</ID>562 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>561 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>856</ID>
<type>AE_DFF_LOW</type>
<position>350.5,-1841.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>560 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>857</ID>
<type>BA_TRI_STATE</type>
<position>375,-1851.5</position>
<input>
<ID>ENABLE_0</ID>559 </input>
<input>
<ID>IN_0</ID>560 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>858</ID>
<type>AA_AND2</type>
<position>360.5,-1851.5</position>
<input>
<ID>IN_0</ID>560 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>559 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>859</ID>
<type>AE_DFF_LOW</type>
<position>424,-1841.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>562 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>860</ID>
<type>BA_TRI_STATE</type>
<position>448.5,-1851.5</position>
<input>
<ID>ENABLE_0</ID>561 </input>
<input>
<ID>IN_0</ID>562 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>861</ID>
<type>AA_AND2</type>
<position>592.5,-1853.5</position>
<input>
<ID>IN_0</ID>566 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>565 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>862</ID>
<type>AE_DFF_LOW</type>
<position>508.5,-1841.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>564 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>863</ID>
<type>BA_TRI_STATE</type>
<position>533,-1853.5</position>
<input>
<ID>ENABLE_0</ID>563 </input>
<input>
<ID>IN_0</ID>564 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>864</ID>
<type>AA_AND2</type>
<position>518.5,-1853.5</position>
<input>
<ID>IN_0</ID>564 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>563 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>865</ID>
<type>AE_DFF_LOW</type>
<position>582,-1841.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>566 </output>
<input>
<ID>clock</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>866</ID>
<type>BA_TRI_STATE</type>
<position>606.5,-1853.5</position>
<input>
<ID>ENABLE_0</ID>565 </input>
<input>
<ID>IN_0</ID>566 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>867</ID>
<type>AA_AND2</type>
<position>-4,-1842.5</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>567 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>868</ID>
<type>BA_TRI_STATE</type>
<position>-25.5,-1861.5</position>
<input>
<ID>ENABLE_0</ID>549 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>550 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>869</ID>
<type>AA_AND2</type>
<position>108.5,-1758</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>572 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>870</ID>
<type>AE_DFF_LOW</type>
<position>24.5,-1751.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>571 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>871</ID>
<type>BA_TRI_STATE</type>
<position>49,-1758</position>
<input>
<ID>ENABLE_0</ID>570 </input>
<input>
<ID>IN_0</ID>571 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>872</ID>
<type>AA_AND2</type>
<position>34.5,-1758</position>
<input>
<ID>IN_0</ID>571 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>570 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>873</ID>
<type>AE_DFF_LOW</type>
<position>98,-1751.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>573 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>874</ID>
<type>BA_TRI_STATE</type>
<position>122.5,-1758</position>
<input>
<ID>ENABLE_0</ID>572 </input>
<input>
<ID>IN_0</ID>573 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>875</ID>
<type>AA_AND2</type>
<position>266.5,-1760</position>
<input>
<ID>IN_0</ID>577 </input>
<input>
<ID>IN_1</ID>569 </input>
<output>
<ID>OUT</ID>576 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>876</ID>
<type>AE_DFF_LOW</type>
<position>182.5,-1751.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>575 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>877</ID>
<type>BA_TRI_STATE</type>
<position>207,-1760</position>
<input>
<ID>ENABLE_0</ID>574 </input>
<input>
<ID>IN_0</ID>575 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>878</ID>
<type>AA_AND2</type>
<position>192,-2631.5</position>
<input>
<ID>IN_0</ID>727 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>726 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>879</ID>
<type>AE_DFF_LOW</type>
<position>256.5,-2623</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>729 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>880</ID>
<type>BA_TRI_STATE</type>
<position>280,-2631.5</position>
<input>
<ID>ENABLE_0</ID>728 </input>
<input>
<ID>IN_0</ID>729 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>881</ID>
<type>AA_AND2</type>
<position>431,-2633</position>
<input>
<ID>IN_0</ID>733 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>732 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>882</ID>
<type>AE_DFF_LOW</type>
<position>347,-2623</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>731 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>883</ID>
<type>BA_TRI_STATE</type>
<position>371.5,-2633</position>
<input>
<ID>ENABLE_0</ID>730 </input>
<input>
<ID>IN_0</ID>731 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>884</ID>
<type>AA_AND2</type>
<position>357,-2633</position>
<input>
<ID>IN_0</ID>731 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>730 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>885</ID>
<type>AE_DFF_LOW</type>
<position>420.5,-2623</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>733 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>886</ID>
<type>BA_TRI_STATE</type>
<position>445,-2633</position>
<input>
<ID>ENABLE_0</ID>732 </input>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>887</ID>
<type>AA_AND2</type>
<position>589,-2635</position>
<input>
<ID>IN_0</ID>737 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>736 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>888</ID>
<type>AE_DFF_LOW</type>
<position>505,-2623</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>735 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>889</ID>
<type>BA_TRI_STATE</type>
<position>529.5,-2635</position>
<input>
<ID>ENABLE_0</ID>734 </input>
<input>
<ID>IN_0</ID>735 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>890</ID>
<type>AA_AND2</type>
<position>515,-2635</position>
<input>
<ID>IN_0</ID>735 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>734 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>891</ID>
<type>AE_DFF_LOW</type>
<position>578.5,-2623</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>737 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>892</ID>
<type>BA_TRI_STATE</type>
<position>603,-2635</position>
<input>
<ID>ENABLE_0</ID>736 </input>
<input>
<ID>IN_0</ID>737 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>893</ID>
<type>AA_AND2</type>
<position>-7.5,-2624</position>
<input>
<ID>IN_0</ID>720 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>894</ID>
<type>BA_TRI_STATE</type>
<position>-29,-2643</position>
<input>
<ID>ENABLE_0</ID>720 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>721 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>895</ID>
<type>AA_AND2</type>
<position>115,-2887.5</position>
<input>
<ID>IN_0</ID>744 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>743 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>896</ID>
<type>AE_DFF_LOW</type>
<position>31,-2881</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>742 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>897</ID>
<type>BA_TRI_STATE</type>
<position>55.5,-2887.5</position>
<input>
<ID>ENABLE_0</ID>741 </input>
<input>
<ID>IN_0</ID>742 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>898</ID>
<type>AA_AND2</type>
<position>41,-2887.5</position>
<input>
<ID>IN_0</ID>742 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>899</ID>
<type>AE_DFF_LOW</type>
<position>104.5,-2881</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>744 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>900</ID>
<type>BA_TRI_STATE</type>
<position>129,-2887.5</position>
<input>
<ID>ENABLE_0</ID>743 </input>
<input>
<ID>IN_0</ID>744 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>901</ID>
<type>AA_AND2</type>
<position>273,-2889.5</position>
<input>
<ID>IN_0</ID>748 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>747 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>902</ID>
<type>AE_DFF_LOW</type>
<position>189,-2881</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>746 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>903</ID>
<type>BA_TRI_STATE</type>
<position>213.5,-2889.5</position>
<input>
<ID>ENABLE_0</ID>745 </input>
<input>
<ID>IN_0</ID>746 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>904</ID>
<type>AA_AND2</type>
<position>199,-2889.5</position>
<input>
<ID>IN_0</ID>746 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>745 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>905</ID>
<type>AE_DFF_LOW</type>
<position>263.5,-2881</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>748 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>906</ID>
<type>BA_TRI_STATE</type>
<position>287,-2889.5</position>
<input>
<ID>ENABLE_0</ID>747 </input>
<input>
<ID>IN_0</ID>748 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>907</ID>
<type>AA_AND2</type>
<position>438,-2891</position>
<input>
<ID>IN_0</ID>752 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>751 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>908</ID>
<type>AE_DFF_LOW</type>
<position>354,-2881</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>750 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>909</ID>
<type>BA_TRI_STATE</type>
<position>378.5,-2891</position>
<input>
<ID>ENABLE_0</ID>749 </input>
<input>
<ID>IN_0</ID>750 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>910</ID>
<type>AA_AND2</type>
<position>364,-2891</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>749 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>911</ID>
<type>AE_DFF_LOW</type>
<position>427.5,-2881</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>752 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>912</ID>
<type>BA_TRI_STATE</type>
<position>452,-2891</position>
<input>
<ID>ENABLE_0</ID>751 </input>
<input>
<ID>IN_0</ID>752 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>913</ID>
<type>AA_AND2</type>
<position>596,-2893</position>
<input>
<ID>IN_0</ID>756 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>755 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>914</ID>
<type>AE_DFF_LOW</type>
<position>512,-2881</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>754 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>915</ID>
<type>BA_TRI_STATE</type>
<position>536.5,-2893</position>
<input>
<ID>ENABLE_0</ID>753 </input>
<input>
<ID>IN_0</ID>754 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>916</ID>
<type>AA_AND2</type>
<position>522,-2893</position>
<input>
<ID>IN_0</ID>754 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>753 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>917</ID>
<type>AE_DFF_LOW</type>
<position>585.5,-2881</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>756 </output>
<input>
<ID>clock</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>918</ID>
<type>BA_TRI_STATE</type>
<position>610,-2893</position>
<input>
<ID>ENABLE_0</ID>755 </input>
<input>
<ID>IN_0</ID>756 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>919</ID>
<type>AA_AND2</type>
<position>-0.5,-2882</position>
<input>
<ID>IN_0</ID>739 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>757 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>920</ID>
<type>BA_TRI_STATE</type>
<position>-22,-2901</position>
<input>
<ID>ENABLE_0</ID>739 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>740 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>921</ID>
<type>AA_AND2</type>
<position>112,-2797.5</position>
<input>
<ID>IN_0</ID>763 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>762 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>922</ID>
<type>AE_DFF_LOW</type>
<position>28,-2791</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>761 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>923</ID>
<type>BA_TRI_STATE</type>
<position>52.5,-2797.5</position>
<input>
<ID>ENABLE_0</ID>760 </input>
<input>
<ID>IN_0</ID>761 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>924</ID>
<type>AA_AND2</type>
<position>38,-2797.5</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>760 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>925</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-2791</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>763 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>926</ID>
<type>BA_TRI_STATE</type>
<position>126,-2797.5</position>
<input>
<ID>ENABLE_0</ID>762 </input>
<input>
<ID>IN_0</ID>763 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>927</ID>
<type>AA_AND2</type>
<position>270,-2799.5</position>
<input>
<ID>IN_0</ID>767 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>928</ID>
<type>AE_DFF_LOW</type>
<position>186,-2791</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>765 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>929</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-2799.5</position>
<input>
<ID>ENABLE_0</ID>764 </input>
<input>
<ID>IN_0</ID>765 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>930</ID>
<type>AA_AND2</type>
<position>196,-2799.5</position>
<input>
<ID>IN_0</ID>765 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>764 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>931</ID>
<type>AE_DFF_LOW</type>
<position>260.5,-2791</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>767 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>932</ID>
<type>BA_TRI_STATE</type>
<position>284,-2799.5</position>
<input>
<ID>ENABLE_0</ID>766 </input>
<input>
<ID>IN_0</ID>767 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>933</ID>
<type>AA_AND2</type>
<position>435,-2801</position>
<input>
<ID>IN_0</ID>771 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>770 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>934</ID>
<type>AE_DFF_LOW</type>
<position>351,-2791</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>769 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>935</ID>
<type>BA_TRI_STATE</type>
<position>375.5,-2801</position>
<input>
<ID>ENABLE_0</ID>768 </input>
<input>
<ID>IN_0</ID>769 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>936</ID>
<type>AA_AND2</type>
<position>361,-2801</position>
<input>
<ID>IN_0</ID>769 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>768 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>937</ID>
<type>AE_DFF_LOW</type>
<position>424.5,-2791</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>771 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>938</ID>
<type>BA_TRI_STATE</type>
<position>449,-2801</position>
<input>
<ID>ENABLE_0</ID>770 </input>
<input>
<ID>IN_0</ID>771 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>939</ID>
<type>AA_AND2</type>
<position>593,-2803</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>774 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>940</ID>
<type>AE_DFF_LOW</type>
<position>509,-2791</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>773 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>941</ID>
<type>BA_TRI_STATE</type>
<position>533.5,-2803</position>
<input>
<ID>ENABLE_0</ID>772 </input>
<input>
<ID>IN_0</ID>773 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>942</ID>
<type>AA_AND2</type>
<position>519,-2803</position>
<input>
<ID>IN_0</ID>773 </input>
<input>
<ID>IN_1</ID>759 </input>
<output>
<ID>OUT</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>943</ID>
<type>AE_DFF_LOW</type>
<position>582.5,-2791</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>775 </output>
<input>
<ID>clock</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>944</ID>
<type>BA_TRI_STATE</type>
<position>607,-2803</position>
<input>
<ID>ENABLE_0</ID>774 </input>
<input>
<ID>IN_0</ID>775 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>945</ID>
<type>AA_AND2</type>
<position>-3.5,-2792</position>
<input>
<ID>IN_0</ID>758 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>776 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>946</ID>
<type>BA_TRI_STATE</type>
<position>-25,-2811</position>
<input>
<ID>ENABLE_0</ID>758 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>759 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>947</ID>
<type>BE_DECODER_3x8</type>
<position>-122.5,-2582.5</position>
<input>
<ID>ENABLE</ID>1396 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>739 </output>
<output>
<ID>OUT_1</ID>758 </output>
<output>
<ID>OUT_2</ID>701 </output>
<output>
<ID>OUT_3</ID>720 </output>
<output>
<ID>OUT_4</ID>663 </output>
<output>
<ID>OUT_5</ID>682 </output>
<output>
<ID>OUT_6</ID>625 </output>
<output>
<ID>OUT_7</ID>644 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>948</ID>
<type>AA_AND2</type>
<position>109,-2343.5</position>
<input>
<ID>IN_0</ID>630 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>629 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>949</ID>
<type>AE_DFF_LOW</type>
<position>25,-2337</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>628 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>950</ID>
<type>BA_TRI_STATE</type>
<position>49.5,-2343.5</position>
<input>
<ID>ENABLE_0</ID>627 </input>
<input>
<ID>IN_0</ID>628 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>951</ID>
<type>AA_AND2</type>
<position>35,-2343.5</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>952</ID>
<type>AE_DFF_LOW</type>
<position>98.5,-2337</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>630 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>953</ID>
<type>BA_TRI_STATE</type>
<position>123,-2343.5</position>
<input>
<ID>ENABLE_0</ID>629 </input>
<input>
<ID>IN_0</ID>630 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>954</ID>
<type>AA_AND2</type>
<position>267,-2345.5</position>
<input>
<ID>IN_0</ID>634 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>633 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>955</ID>
<type>AE_DFF_LOW</type>
<position>183,-2337</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>632 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>956</ID>
<type>BA_TRI_STATE</type>
<position>207.5,-2345.5</position>
<input>
<ID>ENABLE_0</ID>631 </input>
<input>
<ID>IN_0</ID>632 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>957</ID>
<type>AA_AND2</type>
<position>193,-2345.5</position>
<input>
<ID>IN_0</ID>632 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>631 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>958</ID>
<type>AE_DFF_LOW</type>
<position>257.5,-2337</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>634 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>959</ID>
<type>BA_TRI_STATE</type>
<position>281,-2345.5</position>
<input>
<ID>ENABLE_0</ID>633 </input>
<input>
<ID>IN_0</ID>634 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>960</ID>
<type>AA_AND2</type>
<position>432,-2347</position>
<input>
<ID>IN_0</ID>638 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>637 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>961</ID>
<type>AE_DFF_LOW</type>
<position>348,-2337</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>636 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>962</ID>
<type>BA_TRI_STATE</type>
<position>372.5,-2347</position>
<input>
<ID>ENABLE_0</ID>635 </input>
<input>
<ID>IN_0</ID>636 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>963</ID>
<type>AA_AND2</type>
<position>358,-2347</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>635 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>964</ID>
<type>AE_DFF_LOW</type>
<position>421.5,-2337</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>638 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>965</ID>
<type>BA_TRI_STATE</type>
<position>446,-2347</position>
<input>
<ID>ENABLE_0</ID>637 </input>
<input>
<ID>IN_0</ID>638 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>966</ID>
<type>AA_AND2</type>
<position>590,-2349</position>
<input>
<ID>IN_0</ID>642 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>967</ID>
<type>AE_DFF_LOW</type>
<position>506,-2337</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>640 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>968</ID>
<type>BA_TRI_STATE</type>
<position>530.5,-2349</position>
<input>
<ID>ENABLE_0</ID>639 </input>
<input>
<ID>IN_0</ID>640 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>969</ID>
<type>AA_AND2</type>
<position>516,-2349</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>639 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>970</ID>
<type>AE_DFF_LOW</type>
<position>579.5,-2337</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>642 </output>
<input>
<ID>clock</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>971</ID>
<type>BA_TRI_STATE</type>
<position>604,-2349</position>
<input>
<ID>ENABLE_0</ID>641 </input>
<input>
<ID>IN_0</ID>642 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>972</ID>
<type>AA_AND2</type>
<position>-6.5,-2338</position>
<input>
<ID>IN_0</ID>625 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>643 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>973</ID>
<type>BA_TRI_STATE</type>
<position>-28,-2357</position>
<input>
<ID>ENABLE_0</ID>625 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>626 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>974</ID>
<type>AA_AND2</type>
<position>106,-2253.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>648 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>975</ID>
<type>AE_DFF_LOW</type>
<position>22,-2247</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>647 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>976</ID>
<type>BA_TRI_STATE</type>
<position>46.5,-2253.5</position>
<input>
<ID>ENABLE_0</ID>646 </input>
<input>
<ID>IN_0</ID>647 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>977</ID>
<type>AA_AND2</type>
<position>32,-2253.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>978</ID>
<type>AE_DFF_LOW</type>
<position>95.5,-2247</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>649 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>979</ID>
<type>BA_TRI_STATE</type>
<position>120,-2253.5</position>
<input>
<ID>ENABLE_0</ID>648 </input>
<input>
<ID>IN_0</ID>649 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>980</ID>
<type>AA_AND2</type>
<position>264,-2255.5</position>
<input>
<ID>IN_0</ID>653 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>981</ID>
<type>AE_DFF_LOW</type>
<position>180,-2247</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>651 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>982</ID>
<type>BA_TRI_STATE</type>
<position>204.5,-2255.5</position>
<input>
<ID>ENABLE_0</ID>650 </input>
<input>
<ID>IN_0</ID>651 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>983</ID>
<type>AA_AND2</type>
<position>190,-2255.5</position>
<input>
<ID>IN_0</ID>651 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>984</ID>
<type>AE_DFF_LOW</type>
<position>254.5,-2247</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>653 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>985</ID>
<type>BA_TRI_STATE</type>
<position>278,-2255.5</position>
<input>
<ID>ENABLE_0</ID>652 </input>
<input>
<ID>IN_0</ID>653 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>986</ID>
<type>AA_AND2</type>
<position>429,-2257</position>
<input>
<ID>IN_0</ID>657 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>656 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>987</ID>
<type>AE_DFF_LOW</type>
<position>345,-2247</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>655 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>988</ID>
<type>BA_TRI_STATE</type>
<position>369.5,-2257</position>
<input>
<ID>ENABLE_0</ID>654 </input>
<input>
<ID>IN_0</ID>655 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>989</ID>
<type>AA_AND2</type>
<position>355,-2257</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>990</ID>
<type>AE_DFF_LOW</type>
<position>418.5,-2247</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>657 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>991</ID>
<type>BA_TRI_STATE</type>
<position>443,-2257</position>
<input>
<ID>ENABLE_0</ID>656 </input>
<input>
<ID>IN_0</ID>657 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>992</ID>
<type>AA_AND2</type>
<position>587,-2259</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>660 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>993</ID>
<type>AE_DFF_LOW</type>
<position>503,-2247</position>
<output>
<ID>OUT_0</ID>659 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>994</ID>
<type>BA_TRI_STATE</type>
<position>527.5,-2259</position>
<input>
<ID>ENABLE_0</ID>658 </input>
<input>
<ID>IN_0</ID>659 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>995</ID>
<type>AA_AND2</type>
<position>513,-2259</position>
<input>
<ID>IN_0</ID>659 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>658 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>996</ID>
<type>AE_DFF_LOW</type>
<position>576.5,-2247</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>661 </output>
<input>
<ID>clock</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>997</ID>
<type>BA_TRI_STATE</type>
<position>601,-2259</position>
<input>
<ID>ENABLE_0</ID>660 </input>
<input>
<ID>IN_0</ID>661 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>998</ID>
<type>AA_AND2</type>
<position>-9.5,-2248</position>
<input>
<ID>IN_0</ID>644 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>662 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>999</ID>
<type>BA_TRI_STATE</type>
<position>-31,-2267</position>
<input>
<ID>ENABLE_0</ID>644 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>645 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1000</ID>
<type>AA_AND2</type>
<position>113,-2511.5</position>
<input>
<ID>IN_0</ID>668 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>667 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1001</ID>
<type>AE_DFF_LOW</type>
<position>29,-2505</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>666 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1002</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-2511.5</position>
<input>
<ID>ENABLE_0</ID>665 </input>
<input>
<ID>IN_0</ID>666 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1003</ID>
<type>AA_AND2</type>
<position>39,-2511.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>665 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1004</ID>
<type>AE_DFF_LOW</type>
<position>102.5,-2505</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>668 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1005</ID>
<type>BA_TRI_STATE</type>
<position>127,-2511.5</position>
<input>
<ID>ENABLE_0</ID>667 </input>
<input>
<ID>IN_0</ID>668 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1006</ID>
<type>AA_AND2</type>
<position>271,-2513.5</position>
<input>
<ID>IN_0</ID>672 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1007</ID>
<type>AE_DFF_LOW</type>
<position>187,-2505</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>670 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1008</ID>
<type>BA_TRI_STATE</type>
<position>211.5,-2513.5</position>
<input>
<ID>ENABLE_0</ID>669 </input>
<input>
<ID>IN_0</ID>670 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1009</ID>
<type>AA_AND2</type>
<position>197,-2513.5</position>
<input>
<ID>IN_0</ID>670 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>669 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1010</ID>
<type>AE_DFF_LOW</type>
<position>261.5,-2505</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>672 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1011</ID>
<type>BA_TRI_STATE</type>
<position>285,-2513.5</position>
<input>
<ID>ENABLE_0</ID>671 </input>
<input>
<ID>IN_0</ID>672 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1012</ID>
<type>AA_AND2</type>
<position>436,-2515</position>
<input>
<ID>IN_0</ID>676 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>675 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1013</ID>
<type>AE_DFF_LOW</type>
<position>352,-2505</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>674 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1014</ID>
<type>BA_TRI_STATE</type>
<position>376.5,-2515</position>
<input>
<ID>ENABLE_0</ID>673 </input>
<input>
<ID>IN_0</ID>674 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1015</ID>
<type>AA_AND2</type>
<position>362,-2515</position>
<input>
<ID>IN_0</ID>674 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>673 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1016</ID>
<type>AE_DFF_LOW</type>
<position>425.5,-2505</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>676 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1017</ID>
<type>BA_TRI_STATE</type>
<position>450,-2515</position>
<input>
<ID>ENABLE_0</ID>675 </input>
<input>
<ID>IN_0</ID>676 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1018</ID>
<type>AA_AND2</type>
<position>594,-2517</position>
<input>
<ID>IN_0</ID>680 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>679 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1019</ID>
<type>AE_DFF_LOW</type>
<position>510,-2505</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>678 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1020</ID>
<type>BA_TRI_STATE</type>
<position>534.5,-2517</position>
<input>
<ID>ENABLE_0</ID>677 </input>
<input>
<ID>IN_0</ID>678 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1021</ID>
<type>AA_AND2</type>
<position>520,-2517</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1022</ID>
<type>AE_DFF_LOW</type>
<position>583.5,-2505</position>
<input>
<ID>IN_0</ID>1463 </input>
<output>
<ID>OUT_0</ID>680 </output>
<input>
<ID>clock</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1023</ID>
<type>BA_TRI_STATE</type>
<position>608,-2517</position>
<input>
<ID>ENABLE_0</ID>679 </input>
<input>
<ID>IN_0</ID>680 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1024</ID>
<type>AA_AND2</type>
<position>-2.5,-2506</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>681 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1025</ID>
<type>BA_TRI_STATE</type>
<position>-24,-2525</position>
<input>
<ID>ENABLE_0</ID>663 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>664 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1026</ID>
<type>AA_AND2</type>
<position>110,-2421.5</position>
<input>
<ID>IN_0</ID>687 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>686 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1027</ID>
<type>AE_DFF_LOW</type>
<position>26,-2415</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>685 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1028</ID>
<type>BA_TRI_STATE</type>
<position>50.5,-2421.5</position>
<input>
<ID>ENABLE_0</ID>684 </input>
<input>
<ID>IN_0</ID>685 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1029</ID>
<type>AA_AND2</type>
<position>36,-2421.5</position>
<input>
<ID>IN_0</ID>685 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>684 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1030</ID>
<type>AE_DFF_LOW</type>
<position>99.5,-2415</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>687 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1031</ID>
<type>BA_TRI_STATE</type>
<position>124,-2421.5</position>
<input>
<ID>ENABLE_0</ID>686 </input>
<input>
<ID>IN_0</ID>687 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1032</ID>
<type>AA_AND2</type>
<position>268,-2423.5</position>
<input>
<ID>IN_0</ID>691 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>690 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1033</ID>
<type>AE_DFF_LOW</type>
<position>184,-2415</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>689 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1034</ID>
<type>BA_TRI_STATE</type>
<position>208.5,-2423.5</position>
<input>
<ID>ENABLE_0</ID>688 </input>
<input>
<ID>IN_0</ID>689 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1035</ID>
<type>AA_AND2</type>
<position>194,-2423.5</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>688 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1036</ID>
<type>AE_DFF_LOW</type>
<position>258.5,-2415</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>691 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1037</ID>
<type>BA_TRI_STATE</type>
<position>282,-2423.5</position>
<input>
<ID>ENABLE_0</ID>690 </input>
<input>
<ID>IN_0</ID>691 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1038</ID>
<type>AA_AND2</type>
<position>433,-2425</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>694 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1039</ID>
<type>AE_DFF_LOW</type>
<position>349,-2415</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>693 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1040</ID>
<type>BA_TRI_STATE</type>
<position>373.5,-2425</position>
<input>
<ID>ENABLE_0</ID>692 </input>
<input>
<ID>IN_0</ID>693 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1041</ID>
<type>AA_AND2</type>
<position>359,-2425</position>
<input>
<ID>IN_0</ID>693 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>692 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1042</ID>
<type>AE_DFF_LOW</type>
<position>422.5,-2415</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>695 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1043</ID>
<type>BA_TRI_STATE</type>
<position>447,-2425</position>
<input>
<ID>ENABLE_0</ID>694 </input>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1044</ID>
<type>AA_AND2</type>
<position>591,-2427</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1045</ID>
<type>AE_DFF_LOW</type>
<position>507,-2415</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>697 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1046</ID>
<type>BA_TRI_STATE</type>
<position>531.5,-2427</position>
<input>
<ID>ENABLE_0</ID>696 </input>
<input>
<ID>IN_0</ID>697 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1047</ID>
<type>AA_AND2</type>
<position>517,-2427</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>696 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1048</ID>
<type>AE_DFF_LOW</type>
<position>580.5,-2415</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>699 </output>
<input>
<ID>clock</ID>700 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1049</ID>
<type>BA_TRI_STATE</type>
<position>605,-2427</position>
<input>
<ID>ENABLE_0</ID>698 </input>
<input>
<ID>IN_0</ID>699 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1050</ID>
<type>AA_AND2</type>
<position>-5.5,-2416</position>
<input>
<ID>IN_0</ID>682 </input>
<output>
<ID>OUT</ID>700 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1051</ID>
<type>BA_TRI_STATE</type>
<position>-27,-2435</position>
<input>
<ID>ENABLE_0</ID>682 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>683 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1052</ID>
<type>AA_AND2</type>
<position>111,-2719.5</position>
<input>
<ID>IN_0</ID>706 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>705 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1053</ID>
<type>AE_DFF_LOW</type>
<position>27,-2713</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>704 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1054</ID>
<type>BA_TRI_STATE</type>
<position>51.5,-2719.5</position>
<input>
<ID>ENABLE_0</ID>703 </input>
<input>
<ID>IN_0</ID>704 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1055</ID>
<type>AA_AND2</type>
<position>37,-2719.5</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>703 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1056</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-2713</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>706 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1057</ID>
<type>BA_TRI_STATE</type>
<position>125,-2719.5</position>
<input>
<ID>ENABLE_0</ID>705 </input>
<input>
<ID>IN_0</ID>706 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1058</ID>
<type>AA_AND2</type>
<position>269,-2721.5</position>
<input>
<ID>IN_0</ID>710 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1059</ID>
<type>AE_DFF_LOW</type>
<position>185,-2713</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>708 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1060</ID>
<type>BA_TRI_STATE</type>
<position>209.5,-2721.5</position>
<input>
<ID>ENABLE_0</ID>707 </input>
<input>
<ID>IN_0</ID>708 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1061</ID>
<type>AA_AND2</type>
<position>195,-2721.5</position>
<input>
<ID>IN_0</ID>708 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>707 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1062</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-2713</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>710 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1063</ID>
<type>BA_TRI_STATE</type>
<position>283,-2721.5</position>
<input>
<ID>ENABLE_0</ID>709 </input>
<input>
<ID>IN_0</ID>710 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1064</ID>
<type>AA_AND2</type>
<position>434,-2723</position>
<input>
<ID>IN_0</ID>714 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>713 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1065</ID>
<type>AE_DFF_LOW</type>
<position>350,-2713</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>712 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1066</ID>
<type>BA_TRI_STATE</type>
<position>374.5,-2723</position>
<input>
<ID>ENABLE_0</ID>711 </input>
<input>
<ID>IN_0</ID>712 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1067</ID>
<type>AA_AND2</type>
<position>360,-2723</position>
<input>
<ID>IN_0</ID>712 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>711 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1068</ID>
<type>AE_DFF_LOW</type>
<position>423.5,-2713</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>714 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1069</ID>
<type>BA_TRI_STATE</type>
<position>448,-2723</position>
<input>
<ID>ENABLE_0</ID>713 </input>
<input>
<ID>IN_0</ID>714 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1070</ID>
<type>AA_AND2</type>
<position>592,-2725</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>717 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1071</ID>
<type>AE_DFF_LOW</type>
<position>508,-2713</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>716 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1072</ID>
<type>BA_TRI_STATE</type>
<position>532.5,-2725</position>
<input>
<ID>ENABLE_0</ID>715 </input>
<input>
<ID>IN_0</ID>716 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1073</ID>
<type>AA_AND2</type>
<position>518,-2725</position>
<input>
<ID>IN_0</ID>716 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>715 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1074</ID>
<type>AE_DFF_LOW</type>
<position>581.5,-2713</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>718 </output>
<input>
<ID>clock</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1075</ID>
<type>BA_TRI_STATE</type>
<position>606,-2725</position>
<input>
<ID>ENABLE_0</ID>717 </input>
<input>
<ID>IN_0</ID>718 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1076</ID>
<type>AA_AND2</type>
<position>-4.5,-2714</position>
<input>
<ID>IN_0</ID>701 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>719 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1077</ID>
<type>BA_TRI_STATE</type>
<position>-26,-2733</position>
<input>
<ID>ENABLE_0</ID>701 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>702 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1078</ID>
<type>AA_AND2</type>
<position>108,-2629.5</position>
<input>
<ID>IN_0</ID>725 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>724 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1079</ID>
<type>AE_DFF_LOW</type>
<position>24,-2623</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>723 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1080</ID>
<type>BA_TRI_STATE</type>
<position>48.5,-2629.5</position>
<input>
<ID>ENABLE_0</ID>1457 </input>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1081</ID>
<type>AA_AND2</type>
<position>34,-2629.5</position>
<input>
<ID>IN_0</ID>723 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>1457 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1082</ID>
<type>AE_DFF_LOW</type>
<position>97.5,-2623</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>725 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1083</ID>
<type>BA_TRI_STATE</type>
<position>122,-2629.5</position>
<input>
<ID>ENABLE_0</ID>724 </input>
<input>
<ID>IN_0</ID>725 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1084</ID>
<type>AA_AND2</type>
<position>266,-2631.5</position>
<input>
<ID>IN_0</ID>729 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>728 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1085</ID>
<type>AE_DFF_LOW</type>
<position>182,-2623</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>727 </output>
<input>
<ID>clock</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1086</ID>
<type>BA_TRI_STATE</type>
<position>206.5,-2631.5</position>
<input>
<ID>ENABLE_0</ID>726 </input>
<input>
<ID>IN_0</ID>727 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1087</ID>
<type>AA_AND2</type>
<position>110,-3237.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1088</ID>
<type>AE_DFF_LOW</type>
<position>26,-3231</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>780 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1089</ID>
<type>BA_TRI_STATE</type>
<position>50.5,-3237.5</position>
<input>
<ID>ENABLE_0</ID>779 </input>
<input>
<ID>IN_0</ID>780 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1090</ID>
<type>AA_AND2</type>
<position>36,-3237.5</position>
<input>
<ID>IN_0</ID>780 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>779 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1091</ID>
<type>AE_DFF_LOW</type>
<position>99.5,-3231</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>782 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1092</ID>
<type>BA_TRI_STATE</type>
<position>124,-3237.5</position>
<input>
<ID>ENABLE_0</ID>781 </input>
<input>
<ID>IN_0</ID>782 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1093</ID>
<type>AA_AND2</type>
<position>268,-3239.5</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>785 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1094</ID>
<type>AE_DFF_LOW</type>
<position>184,-3231</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>784 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1095</ID>
<type>BA_TRI_STATE</type>
<position>208.5,-3239.5</position>
<input>
<ID>ENABLE_0</ID>783 </input>
<input>
<ID>IN_0</ID>784 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1096</ID>
<type>AA_AND2</type>
<position>194,-3239.5</position>
<input>
<ID>IN_0</ID>784 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1097</ID>
<type>AE_DFF_LOW</type>
<position>258.5,-3231</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>786 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1098</ID>
<type>BA_TRI_STATE</type>
<position>282,-3239.5</position>
<input>
<ID>ENABLE_0</ID>785 </input>
<input>
<ID>IN_0</ID>786 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1099</ID>
<type>AA_AND2</type>
<position>433,-3241</position>
<input>
<ID>IN_0</ID>790 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>789 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1100</ID>
<type>AE_DFF_LOW</type>
<position>349,-3231</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>788 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1101</ID>
<type>BA_TRI_STATE</type>
<position>373.5,-3241</position>
<input>
<ID>ENABLE_0</ID>787 </input>
<input>
<ID>IN_0</ID>788 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1102</ID>
<type>AA_AND2</type>
<position>359,-3241</position>
<input>
<ID>IN_0</ID>788 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>787 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1103</ID>
<type>AE_DFF_LOW</type>
<position>422.5,-3231</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>790 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1104</ID>
<type>BA_TRI_STATE</type>
<position>447,-3241</position>
<input>
<ID>ENABLE_0</ID>789 </input>
<input>
<ID>IN_0</ID>790 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1105</ID>
<type>AA_AND2</type>
<position>591,-3243</position>
<input>
<ID>IN_0</ID>794 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1106</ID>
<type>AE_DFF_LOW</type>
<position>507,-3231</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>792 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1107</ID>
<type>BA_TRI_STATE</type>
<position>531.5,-3243</position>
<input>
<ID>ENABLE_0</ID>791 </input>
<input>
<ID>IN_0</ID>792 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1108</ID>
<type>AA_AND2</type>
<position>517,-3243</position>
<input>
<ID>IN_0</ID>792 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>791 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1109</ID>
<type>AE_DFF_LOW</type>
<position>580.5,-3231</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>794 </output>
<input>
<ID>clock</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1110</ID>
<type>BA_TRI_STATE</type>
<position>605,-3243</position>
<input>
<ID>ENABLE_0</ID>793 </input>
<input>
<ID>IN_0</ID>794 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1111</ID>
<type>AA_AND2</type>
<position>-5.5,-3232</position>
<input>
<ID>IN_0</ID>777 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>795 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1112</ID>
<type>BA_TRI_STATE</type>
<position>-27,-3251</position>
<input>
<ID>ENABLE_0</ID>777 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>778 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1113</ID>
<type>AA_AND2</type>
<position>107,-3147.5</position>
<input>
<ID>IN_0</ID>801 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>800 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1114</ID>
<type>AE_DFF_LOW</type>
<position>23,-3141</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>799 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1115</ID>
<type>BA_TRI_STATE</type>
<position>47.5,-3147.5</position>
<input>
<ID>ENABLE_0</ID>798 </input>
<input>
<ID>IN_0</ID>799 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1116</ID>
<type>AA_AND2</type>
<position>33,-3147.5</position>
<input>
<ID>IN_0</ID>799 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>798 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1117</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-3141</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>801 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1118</ID>
<type>BA_TRI_STATE</type>
<position>121,-3147.5</position>
<input>
<ID>ENABLE_0</ID>800 </input>
<input>
<ID>IN_0</ID>801 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1119</ID>
<type>AA_AND2</type>
<position>265,-3149.5</position>
<input>
<ID>IN_0</ID>805 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>804 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1120</ID>
<type>AE_DFF_LOW</type>
<position>181,-3141</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>803 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1121</ID>
<type>BA_TRI_STATE</type>
<position>205.5,-3149.5</position>
<input>
<ID>ENABLE_0</ID>802 </input>
<input>
<ID>IN_0</ID>803 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1122</ID>
<type>AA_AND2</type>
<position>191,-3149.5</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>802 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1123</ID>
<type>AE_DFF_LOW</type>
<position>255.5,-3141</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>805 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1124</ID>
<type>BA_TRI_STATE</type>
<position>279,-3149.5</position>
<input>
<ID>ENABLE_0</ID>804 </input>
<input>
<ID>IN_0</ID>805 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1125</ID>
<type>AA_AND2</type>
<position>430,-3151</position>
<input>
<ID>IN_0</ID>809 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>808 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1126</ID>
<type>AE_DFF_LOW</type>
<position>346,-3141</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>807 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1127</ID>
<type>BA_TRI_STATE</type>
<position>370.5,-3151</position>
<input>
<ID>ENABLE_0</ID>806 </input>
<input>
<ID>IN_0</ID>807 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1128</ID>
<type>AA_AND2</type>
<position>356,-3151</position>
<input>
<ID>IN_0</ID>807 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>806 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1129</ID>
<type>AE_DFF_LOW</type>
<position>419.5,-3141</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>809 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1130</ID>
<type>BA_TRI_STATE</type>
<position>444,-3151</position>
<input>
<ID>ENABLE_0</ID>808 </input>
<input>
<ID>IN_0</ID>809 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1131</ID>
<type>AA_AND2</type>
<position>588,-3153</position>
<input>
<ID>IN_0</ID>813 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>812 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1132</ID>
<type>AE_DFF_LOW</type>
<position>504,-3141</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>811 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1133</ID>
<type>BA_TRI_STATE</type>
<position>528.5,-3153</position>
<input>
<ID>ENABLE_0</ID>810 </input>
<input>
<ID>IN_0</ID>811 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1134</ID>
<type>AA_AND2</type>
<position>514,-3153</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>810 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1135</ID>
<type>AE_DFF_LOW</type>
<position>577.5,-3141</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>813 </output>
<input>
<ID>clock</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1136</ID>
<type>BA_TRI_STATE</type>
<position>602,-3153</position>
<input>
<ID>ENABLE_0</ID>812 </input>
<input>
<ID>IN_0</ID>813 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1137</ID>
<type>AA_AND2</type>
<position>-8.5,-3142</position>
<input>
<ID>IN_0</ID>796 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>814 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1138</ID>
<type>BA_TRI_STATE</type>
<position>-30,-3161</position>
<input>
<ID>ENABLE_0</ID>796 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>797 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1139</ID>
<type>AA_AND2</type>
<position>114,-3405.5</position>
<input>
<ID>IN_0</ID>820 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1140</ID>
<type>AE_DFF_LOW</type>
<position>30,-3399</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>818 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1141</ID>
<type>BA_TRI_STATE</type>
<position>54.5,-3405.5</position>
<input>
<ID>ENABLE_0</ID>817 </input>
<input>
<ID>IN_0</ID>818 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1142</ID>
<type>AA_AND2</type>
<position>40,-3405.5</position>
<input>
<ID>IN_0</ID>818 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1143</ID>
<type>AE_DFF_LOW</type>
<position>103.5,-3399</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>820 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1144</ID>
<type>BA_TRI_STATE</type>
<position>128,-3405.5</position>
<input>
<ID>ENABLE_0</ID>819 </input>
<input>
<ID>IN_0</ID>820 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1145</ID>
<type>AA_AND2</type>
<position>272,-3407.5</position>
<input>
<ID>IN_0</ID>824 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>823 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1146</ID>
<type>AE_DFF_LOW</type>
<position>188,-3399</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>822 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1147</ID>
<type>BA_TRI_STATE</type>
<position>212.5,-3407.5</position>
<input>
<ID>ENABLE_0</ID>821 </input>
<input>
<ID>IN_0</ID>822 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1148</ID>
<type>AA_AND2</type>
<position>198,-3407.5</position>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>821 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1149</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-3399</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>824 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1150</ID>
<type>BA_TRI_STATE</type>
<position>286,-3407.5</position>
<input>
<ID>ENABLE_0</ID>823 </input>
<input>
<ID>IN_0</ID>824 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1151</ID>
<type>AA_AND2</type>
<position>437,-3409</position>
<input>
<ID>IN_0</ID>828 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>827 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1152</ID>
<type>AE_DFF_LOW</type>
<position>353,-3399</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>826 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1153</ID>
<type>BA_TRI_STATE</type>
<position>377.5,-3409</position>
<input>
<ID>ENABLE_0</ID>825 </input>
<input>
<ID>IN_0</ID>826 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1154</ID>
<type>AA_AND2</type>
<position>363,-3409</position>
<input>
<ID>IN_0</ID>826 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>825 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1155</ID>
<type>AE_DFF_LOW</type>
<position>426.5,-3399</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>828 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1156</ID>
<type>BA_TRI_STATE</type>
<position>451,-3409</position>
<input>
<ID>ENABLE_0</ID>827 </input>
<input>
<ID>IN_0</ID>828 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1157</ID>
<type>AA_AND2</type>
<position>595,-3411</position>
<input>
<ID>IN_0</ID>832 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>831 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1158</ID>
<type>AE_DFF_LOW</type>
<position>511,-3399</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>830 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1159</ID>
<type>BA_TRI_STATE</type>
<position>535.5,-3411</position>
<input>
<ID>ENABLE_0</ID>829 </input>
<input>
<ID>IN_0</ID>830 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1160</ID>
<type>AA_AND2</type>
<position>521,-3411</position>
<input>
<ID>IN_0</ID>830 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>829 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1161</ID>
<type>AE_DFF_LOW</type>
<position>584.5,-3399</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>832 </output>
<input>
<ID>clock</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1162</ID>
<type>BA_TRI_STATE</type>
<position>609,-3411</position>
<input>
<ID>ENABLE_0</ID>831 </input>
<input>
<ID>IN_0</ID>832 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1163</ID>
<type>AA_AND2</type>
<position>-1.5,-3400</position>
<input>
<ID>IN_0</ID>815 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>833 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1164</ID>
<type>BA_TRI_STATE</type>
<position>-23,-3419</position>
<input>
<ID>ENABLE_0</ID>815 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>816 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1165</ID>
<type>AA_AND2</type>
<position>111,-3315.5</position>
<input>
<ID>IN_0</ID>839 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>838 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1166</ID>
<type>AE_DFF_LOW</type>
<position>27,-3309</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>837 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1167</ID>
<type>BA_TRI_STATE</type>
<position>51.5,-3315.5</position>
<input>
<ID>ENABLE_0</ID>836 </input>
<input>
<ID>IN_0</ID>837 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1168</ID>
<type>AA_AND2</type>
<position>37,-3315.5</position>
<input>
<ID>IN_0</ID>837 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>836 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1169</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-3309</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>839 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1170</ID>
<type>BA_TRI_STATE</type>
<position>125,-3315.5</position>
<input>
<ID>ENABLE_0</ID>838 </input>
<input>
<ID>IN_0</ID>839 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1171</ID>
<type>AA_AND2</type>
<position>269,-3317.5</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>842 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1172</ID>
<type>AE_DFF_LOW</type>
<position>185,-3309</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>841 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1173</ID>
<type>BA_TRI_STATE</type>
<position>209.5,-3317.5</position>
<input>
<ID>ENABLE_0</ID>840 </input>
<input>
<ID>IN_0</ID>841 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1174</ID>
<type>AA_AND2</type>
<position>195,-3317.5</position>
<input>
<ID>IN_0</ID>841 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>840 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1175</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-3309</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>843 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1176</ID>
<type>BA_TRI_STATE</type>
<position>283,-3317.5</position>
<input>
<ID>ENABLE_0</ID>842 </input>
<input>
<ID>IN_0</ID>843 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1177</ID>
<type>AA_AND2</type>
<position>434,-3319</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>846 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1178</ID>
<type>AE_DFF_LOW</type>
<position>350,-3309</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>845 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1179</ID>
<type>BA_TRI_STATE</type>
<position>374.5,-3319</position>
<input>
<ID>ENABLE_0</ID>844 </input>
<input>
<ID>IN_0</ID>845 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1180</ID>
<type>AA_AND2</type>
<position>360,-3319</position>
<input>
<ID>IN_0</ID>845 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>844 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1181</ID>
<type>AE_DFF_LOW</type>
<position>423.5,-3309</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>847 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1182</ID>
<type>BA_TRI_STATE</type>
<position>448,-3319</position>
<input>
<ID>ENABLE_0</ID>846 </input>
<input>
<ID>IN_0</ID>847 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1183</ID>
<type>AA_AND2</type>
<position>592,-3321</position>
<input>
<ID>IN_0</ID>851 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>850 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1184</ID>
<type>AE_DFF_LOW</type>
<position>508,-3309</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>849 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1185</ID>
<type>BA_TRI_STATE</type>
<position>532.5,-3321</position>
<input>
<ID>ENABLE_0</ID>848 </input>
<input>
<ID>IN_0</ID>849 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1186</ID>
<type>AA_AND2</type>
<position>518,-3321</position>
<input>
<ID>IN_0</ID>849 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>848 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1187</ID>
<type>AE_DFF_LOW</type>
<position>581.5,-3309</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>851 </output>
<input>
<ID>clock</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1188</ID>
<type>BA_TRI_STATE</type>
<position>606,-3321</position>
<input>
<ID>ENABLE_0</ID>850 </input>
<input>
<ID>IN_0</ID>851 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1189</ID>
<type>AA_AND2</type>
<position>-4.5,-3310</position>
<input>
<ID>IN_0</ID>834 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>852 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1190</ID>
<type>BA_TRI_STATE</type>
<position>-26,-3329</position>
<input>
<ID>ENABLE_0</ID>834 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>835 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1191</ID>
<type>AA_AND2</type>
<position>112,-3613.5</position>
<input>
<ID>IN_0</ID>858 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>857 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1192</ID>
<type>AE_DFF_LOW</type>
<position>28,-3607</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>856 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1193</ID>
<type>BA_TRI_STATE</type>
<position>52.5,-3613.5</position>
<input>
<ID>ENABLE_0</ID>855 </input>
<input>
<ID>IN_0</ID>856 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1194</ID>
<type>AA_AND2</type>
<position>38,-3613.5</position>
<input>
<ID>IN_0</ID>856 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>855 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1195</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-3607</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>858 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1196</ID>
<type>BA_TRI_STATE</type>
<position>126,-3613.5</position>
<input>
<ID>ENABLE_0</ID>857 </input>
<input>
<ID>IN_0</ID>858 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1197</ID>
<type>AA_AND2</type>
<position>270,-3615.5</position>
<input>
<ID>IN_0</ID>862 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>861 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1198</ID>
<type>AE_DFF_LOW</type>
<position>186,-3607</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>860 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1199</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-3615.5</position>
<input>
<ID>ENABLE_0</ID>859 </input>
<input>
<ID>IN_0</ID>860 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1200</ID>
<type>AA_AND2</type>
<position>196,-3615.5</position>
<input>
<ID>IN_0</ID>860 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>859 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1201</ID>
<type>AE_DFF_LOW</type>
<position>260.5,-3607</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>862 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1202</ID>
<type>BA_TRI_STATE</type>
<position>284,-3615.5</position>
<input>
<ID>ENABLE_0</ID>861 </input>
<input>
<ID>IN_0</ID>862 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1203</ID>
<type>AA_AND2</type>
<position>435,-3617</position>
<input>
<ID>IN_0</ID>866 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>865 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1204</ID>
<type>AE_DFF_LOW</type>
<position>351,-3607</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>864 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1205</ID>
<type>BA_TRI_STATE</type>
<position>375.5,-3617</position>
<input>
<ID>ENABLE_0</ID>863 </input>
<input>
<ID>IN_0</ID>864 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1206</ID>
<type>AA_AND2</type>
<position>361,-3617</position>
<input>
<ID>IN_0</ID>864 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>863 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1207</ID>
<type>AE_DFF_LOW</type>
<position>424.5,-3607</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>866 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1208</ID>
<type>BA_TRI_STATE</type>
<position>449,-3617</position>
<input>
<ID>ENABLE_0</ID>865 </input>
<input>
<ID>IN_0</ID>866 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1209</ID>
<type>AA_AND2</type>
<position>593,-3619</position>
<input>
<ID>IN_0</ID>870 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>869 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1210</ID>
<type>AE_DFF_LOW</type>
<position>509,-3607</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>868 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1211</ID>
<type>BA_TRI_STATE</type>
<position>533.5,-3619</position>
<input>
<ID>ENABLE_0</ID>867 </input>
<input>
<ID>IN_0</ID>868 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1212</ID>
<type>AA_AND2</type>
<position>519,-3619</position>
<input>
<ID>IN_0</ID>868 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>867 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1213</ID>
<type>AE_DFF_LOW</type>
<position>582.5,-3607</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>870 </output>
<input>
<ID>clock</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1214</ID>
<type>BA_TRI_STATE</type>
<position>607,-3619</position>
<input>
<ID>ENABLE_0</ID>869 </input>
<input>
<ID>IN_0</ID>870 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1215</ID>
<type>AA_AND2</type>
<position>-3.5,-3608</position>
<input>
<ID>IN_0</ID>853 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>871 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1216</ID>
<type>BA_TRI_STATE</type>
<position>-25,-3627</position>
<input>
<ID>ENABLE_0</ID>853 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>854 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1217</ID>
<type>AA_AND2</type>
<position>109,-3523.5</position>
<input>
<ID>IN_0</ID>877 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>876 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1218</ID>
<type>AE_DFF_LOW</type>
<position>25,-3517</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>875 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1219</ID>
<type>BA_TRI_STATE</type>
<position>49.5,-3523.5</position>
<input>
<ID>ENABLE_0</ID>874 </input>
<input>
<ID>IN_0</ID>875 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1220</ID>
<type>AA_AND2</type>
<position>35,-3523.5</position>
<input>
<ID>IN_0</ID>875 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>874 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1221</ID>
<type>AE_DFF_LOW</type>
<position>98.5,-3517</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>877 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1222</ID>
<type>BA_TRI_STATE</type>
<position>123,-3523.5</position>
<input>
<ID>ENABLE_0</ID>876 </input>
<input>
<ID>IN_0</ID>877 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1223</ID>
<type>AA_AND2</type>
<position>267,-3525.5</position>
<input>
<ID>IN_0</ID>881 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>880 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1224</ID>
<type>AE_DFF_LOW</type>
<position>183,-3517</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>879 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1225</ID>
<type>BA_TRI_STATE</type>
<position>207.5,-3525.5</position>
<input>
<ID>ENABLE_0</ID>878 </input>
<input>
<ID>IN_0</ID>879 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1226</ID>
<type>AA_AND2</type>
<position>193,-3525.5</position>
<input>
<ID>IN_0</ID>879 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>878 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1227</ID>
<type>AE_DFF_LOW</type>
<position>257.5,-3517</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>881 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1228</ID>
<type>BA_TRI_STATE</type>
<position>281,-3525.5</position>
<input>
<ID>ENABLE_0</ID>880 </input>
<input>
<ID>IN_0</ID>881 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1229</ID>
<type>AA_AND2</type>
<position>432,-3527</position>
<input>
<ID>IN_0</ID>885 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1230</ID>
<type>AE_DFF_LOW</type>
<position>348,-3517</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>883 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1231</ID>
<type>BA_TRI_STATE</type>
<position>372.5,-3527</position>
<input>
<ID>ENABLE_0</ID>882 </input>
<input>
<ID>IN_0</ID>883 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1232</ID>
<type>AA_AND2</type>
<position>358,-3527</position>
<input>
<ID>IN_0</ID>883 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>882 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1233</ID>
<type>AE_DFF_LOW</type>
<position>421.5,-3517</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>885 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1234</ID>
<type>BA_TRI_STATE</type>
<position>446,-3527</position>
<input>
<ID>ENABLE_0</ID>884 </input>
<input>
<ID>IN_0</ID>885 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1235</ID>
<type>AA_AND2</type>
<position>590,-3529</position>
<input>
<ID>IN_0</ID>889 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>888 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1236</ID>
<type>AE_DFF_LOW</type>
<position>506,-3517</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>887 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1237</ID>
<type>BA_TRI_STATE</type>
<position>530.5,-3529</position>
<input>
<ID>ENABLE_0</ID>886 </input>
<input>
<ID>IN_0</ID>887 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1238</ID>
<type>AA_AND2</type>
<position>516,-3529</position>
<input>
<ID>IN_0</ID>887 </input>
<input>
<ID>IN_1</ID>873 </input>
<output>
<ID>OUT</ID>886 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1239</ID>
<type>AE_DFF_LOW</type>
<position>579.5,-3517</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>889 </output>
<input>
<ID>clock</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1240</ID>
<type>BA_TRI_STATE</type>
<position>604,-3529</position>
<input>
<ID>ENABLE_0</ID>888 </input>
<input>
<ID>IN_0</ID>889 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1241</ID>
<type>AA_AND2</type>
<position>-6.5,-3518</position>
<input>
<ID>IN_0</ID>872 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>890 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1242</ID>
<type>BA_TRI_STATE</type>
<position>-28,-3537</position>
<input>
<ID>ENABLE_0</ID>872 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>873 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1243</ID>
<type>AA_AND2</type>
<position>116,-3781.5</position>
<input>
<ID>IN_0</ID>896 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>895 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1244</ID>
<type>AE_DFF_LOW</type>
<position>32,-3775</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>894 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1245</ID>
<type>BA_TRI_STATE</type>
<position>56.5,-3781.5</position>
<input>
<ID>ENABLE_0</ID>893 </input>
<input>
<ID>IN_0</ID>894 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1246</ID>
<type>AA_AND2</type>
<position>42,-3781.5</position>
<input>
<ID>IN_0</ID>894 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>893 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1247</ID>
<type>AE_DFF_LOW</type>
<position>105.5,-3775</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>896 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1248</ID>
<type>BA_TRI_STATE</type>
<position>130,-3781.5</position>
<input>
<ID>ENABLE_0</ID>895 </input>
<input>
<ID>IN_0</ID>896 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1249</ID>
<type>AA_AND2</type>
<position>274,-3783.5</position>
<input>
<ID>IN_0</ID>900 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>899 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1250</ID>
<type>AE_DFF_LOW</type>
<position>190,-3775</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>898 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1251</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-3783.5</position>
<input>
<ID>ENABLE_0</ID>897 </input>
<input>
<ID>IN_0</ID>898 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1252</ID>
<type>AA_AND2</type>
<position>200,-3783.5</position>
<input>
<ID>IN_0</ID>898 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>897 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1253</ID>
<type>AE_DFF_LOW</type>
<position>264.5,-3775</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>900 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1254</ID>
<type>BA_TRI_STATE</type>
<position>288,-3783.5</position>
<input>
<ID>ENABLE_0</ID>899 </input>
<input>
<ID>IN_0</ID>900 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1255</ID>
<type>AA_AND2</type>
<position>439,-3785</position>
<input>
<ID>IN_0</ID>904 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>903 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1256</ID>
<type>AE_DFF_LOW</type>
<position>355,-3775</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>902 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1257</ID>
<type>BA_TRI_STATE</type>
<position>379.5,-3785</position>
<input>
<ID>ENABLE_0</ID>901 </input>
<input>
<ID>IN_0</ID>902 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1258</ID>
<type>AA_AND2</type>
<position>365,-3785</position>
<input>
<ID>IN_0</ID>902 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>901 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1259</ID>
<type>AE_DFF_LOW</type>
<position>428.5,-3775</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>904 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1260</ID>
<type>BA_TRI_STATE</type>
<position>453,-3785</position>
<input>
<ID>ENABLE_0</ID>903 </input>
<input>
<ID>IN_0</ID>904 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1261</ID>
<type>AA_AND2</type>
<position>597,-3787</position>
<input>
<ID>IN_0</ID>908 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>907 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1262</ID>
<type>AE_DFF_LOW</type>
<position>513,-3775</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>906 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1263</ID>
<type>BA_TRI_STATE</type>
<position>537.5,-3787</position>
<input>
<ID>ENABLE_0</ID>905 </input>
<input>
<ID>IN_0</ID>906 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1264</ID>
<type>AA_AND2</type>
<position>523,-3787</position>
<input>
<ID>IN_0</ID>906 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>905 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1265</ID>
<type>AE_DFF_LOW</type>
<position>586.5,-3775</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>908 </output>
<input>
<ID>clock</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1266</ID>
<type>BA_TRI_STATE</type>
<position>611,-3787</position>
<input>
<ID>ENABLE_0</ID>907 </input>
<input>
<ID>IN_0</ID>908 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1267</ID>
<type>AA_AND2</type>
<position>0.5,-3776</position>
<input>
<ID>IN_0</ID>891 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>909 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1268</ID>
<type>BA_TRI_STATE</type>
<position>-21,-3795</position>
<input>
<ID>ENABLE_0</ID>891 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>892 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1269</ID>
<type>AA_AND2</type>
<position>113,-3691.5</position>
<input>
<ID>IN_0</ID>915 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>914 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1270</ID>
<type>AE_DFF_LOW</type>
<position>29,-3685</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>913 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1271</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-3691.5</position>
<input>
<ID>ENABLE_0</ID>912 </input>
<input>
<ID>IN_0</ID>913 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1272</ID>
<type>AA_AND2</type>
<position>39,-3691.5</position>
<input>
<ID>IN_0</ID>913 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>912 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1273</ID>
<type>AE_DFF_LOW</type>
<position>102.5,-3685</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>915 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1274</ID>
<type>BA_TRI_STATE</type>
<position>127,-3691.5</position>
<input>
<ID>ENABLE_0</ID>914 </input>
<input>
<ID>IN_0</ID>915 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1275</ID>
<type>AA_AND2</type>
<position>271,-3693.5</position>
<input>
<ID>IN_0</ID>919 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>918 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1276</ID>
<type>AE_DFF_LOW</type>
<position>187,-3685</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>917 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1277</ID>
<type>BA_TRI_STATE</type>
<position>211.5,-3693.5</position>
<input>
<ID>ENABLE_0</ID>916 </input>
<input>
<ID>IN_0</ID>917 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1278</ID>
<type>AA_AND2</type>
<position>197,-3693.5</position>
<input>
<ID>IN_0</ID>917 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>916 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1279</ID>
<type>AE_DFF_LOW</type>
<position>261.5,-3685</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>919 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1280</ID>
<type>BA_TRI_STATE</type>
<position>285,-3693.5</position>
<input>
<ID>ENABLE_0</ID>918 </input>
<input>
<ID>IN_0</ID>919 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1281</ID>
<type>AA_AND2</type>
<position>436,-3695</position>
<input>
<ID>IN_0</ID>923 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>922 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1282</ID>
<type>AE_DFF_LOW</type>
<position>352,-3685</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>921 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1283</ID>
<type>BA_TRI_STATE</type>
<position>376.5,-3695</position>
<input>
<ID>ENABLE_0</ID>920 </input>
<input>
<ID>IN_0</ID>921 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1284</ID>
<type>AA_AND2</type>
<position>362,-3695</position>
<input>
<ID>IN_0</ID>921 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>920 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1285</ID>
<type>AE_DFF_LOW</type>
<position>425.5,-3685</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>923 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1286</ID>
<type>BA_TRI_STATE</type>
<position>450,-3695</position>
<input>
<ID>ENABLE_0</ID>922 </input>
<input>
<ID>IN_0</ID>923 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1287</ID>
<type>AA_AND2</type>
<position>594,-3697</position>
<input>
<ID>IN_0</ID>927 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>926 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1288</ID>
<type>AE_DFF_LOW</type>
<position>510,-3685</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>925 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1289</ID>
<type>BA_TRI_STATE</type>
<position>534.5,-3697</position>
<input>
<ID>ENABLE_0</ID>924 </input>
<input>
<ID>IN_0</ID>925 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1290</ID>
<type>AA_AND2</type>
<position>520,-3697</position>
<input>
<ID>IN_0</ID>925 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>924 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1291</ID>
<type>AE_DFF_LOW</type>
<position>583.5,-3685</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>927 </output>
<input>
<ID>clock</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1292</ID>
<type>BA_TRI_STATE</type>
<position>608,-3697</position>
<input>
<ID>ENABLE_0</ID>926 </input>
<input>
<ID>IN_0</ID>927 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1293</ID>
<type>AA_AND2</type>
<position>-2.5,-3686</position>
<input>
<ID>IN_0</ID>910 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>928 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1294</ID>
<type>BA_TRI_STATE</type>
<position>-24,-3705</position>
<input>
<ID>ENABLE_0</ID>910 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>911 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1295</ID>
<type>BE_DECODER_3x8</type>
<position>-121.5,-3476.5</position>
<input>
<ID>ENABLE</ID>1397 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>891 </output>
<output>
<ID>OUT_1</ID>910 </output>
<output>
<ID>OUT_2</ID>853 </output>
<output>
<ID>OUT_3</ID>872 </output>
<output>
<ID>OUT_4</ID>815 </output>
<output>
<ID>OUT_5</ID>834 </output>
<output>
<ID>OUT_6</ID>777 </output>
<output>
<ID>OUT_7</ID>796 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1296</ID>
<type>AA_AND2</type>
<position>193,-4351</position>
<input>
<ID>IN_0</ID>1031 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1297</ID>
<type>AE_DFF_LOW</type>
<position>257.5,-4342.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1033 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1298</ID>
<type>BA_TRI_STATE</type>
<position>281,-4351</position>
<input>
<ID>ENABLE_0</ID>1032 </input>
<input>
<ID>IN_0</ID>1033 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1299</ID>
<type>AA_AND2</type>
<position>432,-4352.5</position>
<input>
<ID>IN_0</ID>1037 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1036 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1300</ID>
<type>AE_DFF_LOW</type>
<position>348,-4342.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1035 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1301</ID>
<type>BA_TRI_STATE</type>
<position>372.5,-4352.5</position>
<input>
<ID>ENABLE_0</ID>1034 </input>
<input>
<ID>IN_0</ID>1035 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1302</ID>
<type>AA_AND2</type>
<position>358,-4352.5</position>
<input>
<ID>IN_0</ID>1035 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1034 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1303</ID>
<type>AE_DFF_LOW</type>
<position>421.5,-4342.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1037 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1304</ID>
<type>BA_TRI_STATE</type>
<position>446,-4352.5</position>
<input>
<ID>ENABLE_0</ID>1036 </input>
<input>
<ID>IN_0</ID>1037 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1305</ID>
<type>AA_AND2</type>
<position>590,-4354.5</position>
<input>
<ID>IN_0</ID>1041 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1040 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1306</ID>
<type>AE_DFF_LOW</type>
<position>506,-4342.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1039 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1307</ID>
<type>BA_TRI_STATE</type>
<position>530.5,-4354.5</position>
<input>
<ID>ENABLE_0</ID>1038 </input>
<input>
<ID>IN_0</ID>1039 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1308</ID>
<type>AA_AND2</type>
<position>516,-4354.5</position>
<input>
<ID>IN_0</ID>1039 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1038 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1309</ID>
<type>AE_DFF_LOW</type>
<position>579.5,-4342.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1041 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1310</ID>
<type>BA_TRI_STATE</type>
<position>604,-4354.5</position>
<input>
<ID>ENABLE_0</ID>1040 </input>
<input>
<ID>IN_0</ID>1041 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1311</ID>
<type>AA_AND2</type>
<position>-6.5,-4343.5</position>
<input>
<ID>IN_0</ID>1024 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1042 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1312</ID>
<type>BA_TRI_STATE</type>
<position>-28,-4362.5</position>
<input>
<ID>ENABLE_0</ID>1024 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1025 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1313</ID>
<type>AA_AND2</type>
<position>116,-4607</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1047 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1314</ID>
<type>AE_DFF_LOW</type>
<position>32,-4600.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1046 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1315</ID>
<type>BA_TRI_STATE</type>
<position>56.5,-4607</position>
<input>
<ID>ENABLE_0</ID>1045 </input>
<input>
<ID>IN_0</ID>1046 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1316</ID>
<type>AA_AND2</type>
<position>42,-4607</position>
<input>
<ID>IN_0</ID>1046 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1045 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1317</ID>
<type>AE_DFF_LOW</type>
<position>105.5,-4600.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1048 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1318</ID>
<type>BA_TRI_STATE</type>
<position>130,-4607</position>
<input>
<ID>ENABLE_0</ID>1047 </input>
<input>
<ID>IN_0</ID>1048 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1319</ID>
<type>AA_AND2</type>
<position>274,-4609</position>
<input>
<ID>IN_0</ID>1052 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1051 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1320</ID>
<type>AE_DFF_LOW</type>
<position>190,-4600.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1050 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1321</ID>
<type>BA_TRI_STATE</type>
<position>214.5,-4609</position>
<input>
<ID>ENABLE_0</ID>1049 </input>
<input>
<ID>IN_0</ID>1050 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1322</ID>
<type>AA_AND2</type>
<position>200,-4609</position>
<input>
<ID>IN_0</ID>1050 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1049 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1323</ID>
<type>AE_DFF_LOW</type>
<position>264.5,-4600.5</position>
<output>
<ID>OUT_0</ID>1052 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1324</ID>
<type>BA_TRI_STATE</type>
<position>288,-4609</position>
<input>
<ID>ENABLE_0</ID>1051 </input>
<input>
<ID>IN_0</ID>1052 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1325</ID>
<type>AA_AND2</type>
<position>439,-4610.5</position>
<input>
<ID>IN_0</ID>1056 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1055 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1326</ID>
<type>AE_DFF_LOW</type>
<position>355,-4600.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1054 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1327</ID>
<type>BA_TRI_STATE</type>
<position>379.5,-4610.5</position>
<input>
<ID>ENABLE_0</ID>1053 </input>
<input>
<ID>IN_0</ID>1054 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1328</ID>
<type>AA_AND2</type>
<position>365,-4610.5</position>
<input>
<ID>IN_0</ID>1054 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1053 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1329</ID>
<type>AE_DFF_LOW</type>
<position>428.5,-4600.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1056 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1330</ID>
<type>BA_TRI_STATE</type>
<position>453,-4610.5</position>
<input>
<ID>ENABLE_0</ID>1055 </input>
<input>
<ID>IN_0</ID>1056 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1331</ID>
<type>AA_AND2</type>
<position>597,-4612.5</position>
<input>
<ID>IN_0</ID>1060 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1059 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1332</ID>
<type>AE_DFF_LOW</type>
<position>513,-4600.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1058 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1333</ID>
<type>BA_TRI_STATE</type>
<position>537.5,-4612.5</position>
<input>
<ID>ENABLE_0</ID>1057 </input>
<input>
<ID>IN_0</ID>1058 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1334</ID>
<type>AA_AND2</type>
<position>523,-4612.5</position>
<input>
<ID>IN_0</ID>1058 </input>
<input>
<ID>IN_1</ID>1044 </input>
<output>
<ID>OUT</ID>1057 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1335</ID>
<type>AE_DFF_LOW</type>
<position>586.5,-4600.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1060 </output>
<input>
<ID>clock</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1336</ID>
<type>BA_TRI_STATE</type>
<position>611,-4612.5</position>
<input>
<ID>ENABLE_0</ID>1059 </input>
<input>
<ID>IN_0</ID>1060 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1337</ID>
<type>AA_AND2</type>
<position>0.5,-4601.5</position>
<input>
<ID>IN_0</ID>1043 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1338</ID>
<type>BA_TRI_STATE</type>
<position>-21,-4620.5</position>
<input>
<ID>ENABLE_0</ID>1043 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1044 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1339</ID>
<type>AA_AND2</type>
<position>113,-4517</position>
<input>
<ID>IN_0</ID>1067 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1066 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1340</ID>
<type>AE_DFF_LOW</type>
<position>29,-4510.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1065 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1341</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-4517</position>
<input>
<ID>ENABLE_0</ID>1064 </input>
<input>
<ID>IN_0</ID>1065 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1342</ID>
<type>AA_AND2</type>
<position>39,-4517</position>
<input>
<ID>IN_0</ID>1065 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1343</ID>
<type>AE_DFF_LOW</type>
<position>102.5,-4510.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1067 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1344</ID>
<type>BA_TRI_STATE</type>
<position>127,-4517</position>
<input>
<ID>ENABLE_0</ID>1066 </input>
<input>
<ID>IN_0</ID>1067 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1345</ID>
<type>AA_AND2</type>
<position>271,-4519</position>
<input>
<ID>IN_0</ID>1071 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1346</ID>
<type>AE_DFF_LOW</type>
<position>187,-4510.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1069 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1347</ID>
<type>BA_TRI_STATE</type>
<position>211.5,-4519</position>
<input>
<ID>ENABLE_0</ID>1068 </input>
<input>
<ID>IN_0</ID>1069 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1348</ID>
<type>AA_AND2</type>
<position>197,-4519</position>
<input>
<ID>IN_0</ID>1069 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1349</ID>
<type>AE_DFF_LOW</type>
<position>261.5,-4510.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1071 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1350</ID>
<type>BA_TRI_STATE</type>
<position>285,-4519</position>
<input>
<ID>ENABLE_0</ID>1070 </input>
<input>
<ID>IN_0</ID>1071 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1351</ID>
<type>AA_AND2</type>
<position>436,-4520.5</position>
<input>
<ID>IN_0</ID>1075 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1352</ID>
<type>AE_DFF_LOW</type>
<position>352,-4510.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1073 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1353</ID>
<type>BA_TRI_STATE</type>
<position>376.5,-4520.5</position>
<input>
<ID>ENABLE_0</ID>1072 </input>
<input>
<ID>IN_0</ID>1073 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1354</ID>
<type>AA_AND2</type>
<position>362,-4520.5</position>
<input>
<ID>IN_0</ID>1073 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1072 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1355</ID>
<type>AE_DFF_LOW</type>
<position>425.5,-4510.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1075 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1356</ID>
<type>BA_TRI_STATE</type>
<position>450,-4520.5</position>
<input>
<ID>ENABLE_0</ID>1074 </input>
<input>
<ID>IN_0</ID>1075 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1357</ID>
<type>AA_AND2</type>
<position>594,-4522.5</position>
<input>
<ID>IN_0</ID>1079 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1078 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1358</ID>
<type>AE_DFF_LOW</type>
<position>510,-4510.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1077 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1359</ID>
<type>BA_TRI_STATE</type>
<position>534.5,-4522.5</position>
<input>
<ID>ENABLE_0</ID>1076 </input>
<input>
<ID>IN_0</ID>1077 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1360</ID>
<type>AA_AND2</type>
<position>520,-4522.5</position>
<input>
<ID>IN_0</ID>1077 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1076 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1361</ID>
<type>AE_DFF_LOW</type>
<position>583.5,-4510.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1079 </output>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1362</ID>
<type>BA_TRI_STATE</type>
<position>608,-4522.5</position>
<input>
<ID>ENABLE_0</ID>1078 </input>
<input>
<ID>IN_0</ID>1079 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1363</ID>
<type>AA_AND2</type>
<position>-2.5,-4511.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1364</ID>
<type>BA_TRI_STATE</type>
<position>-24,-4530.5</position>
<input>
<ID>ENABLE_0</ID>1062 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1063 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1365</ID>
<type>BE_DECODER_3x8</type>
<position>-121.5,-4302</position>
<input>
<ID>ENABLE</ID>1398 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>1043 </output>
<output>
<ID>OUT_1</ID>1062 </output>
<output>
<ID>OUT_2</ID>1005 </output>
<output>
<ID>OUT_3</ID>1024 </output>
<output>
<ID>OUT_4</ID>967 </output>
<output>
<ID>OUT_5</ID>986 </output>
<output>
<ID>OUT_6</ID>929 </output>
<output>
<ID>OUT_7</ID>948 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1366</ID>
<type>AA_AND2</type>
<position>110,-4063</position>
<input>
<ID>IN_0</ID>934 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>933 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1367</ID>
<type>AE_DFF_LOW</type>
<position>26,-4056.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>932 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1368</ID>
<type>BA_TRI_STATE</type>
<position>50.5,-4063</position>
<input>
<ID>ENABLE_0</ID>931 </input>
<input>
<ID>IN_0</ID>932 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1369</ID>
<type>AA_AND2</type>
<position>36,-4063</position>
<input>
<ID>IN_0</ID>932 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>931 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1370</ID>
<type>AE_DFF_LOW</type>
<position>99.5,-4056.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>934 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1371</ID>
<type>BA_TRI_STATE</type>
<position>124,-4063</position>
<input>
<ID>ENABLE_0</ID>933 </input>
<input>
<ID>IN_0</ID>934 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1372</ID>
<type>AA_AND2</type>
<position>268,-4065</position>
<input>
<ID>IN_0</ID>938 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>937 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1373</ID>
<type>AE_DFF_LOW</type>
<position>184,-4056.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>936 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1374</ID>
<type>BA_TRI_STATE</type>
<position>208.5,-4065</position>
<input>
<ID>ENABLE_0</ID>935 </input>
<input>
<ID>IN_0</ID>936 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1375</ID>
<type>AA_AND2</type>
<position>194,-4065</position>
<input>
<ID>IN_0</ID>936 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>935 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1376</ID>
<type>AE_DFF_LOW</type>
<position>258.5,-4056.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>938 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1377</ID>
<type>BA_TRI_STATE</type>
<position>282,-4065</position>
<input>
<ID>ENABLE_0</ID>937 </input>
<input>
<ID>IN_0</ID>938 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1378</ID>
<type>AA_AND2</type>
<position>433,-4066.5</position>
<input>
<ID>IN_0</ID>942 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>941 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1379</ID>
<type>AE_DFF_LOW</type>
<position>349,-4056.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>940 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1380</ID>
<type>BA_TRI_STATE</type>
<position>373.5,-4066.5</position>
<input>
<ID>ENABLE_0</ID>939 </input>
<input>
<ID>IN_0</ID>940 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1381</ID>
<type>AA_AND2</type>
<position>359,-4066.5</position>
<input>
<ID>IN_0</ID>940 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>939 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1382</ID>
<type>AE_DFF_LOW</type>
<position>422.5,-4056.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>942 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1383</ID>
<type>BA_TRI_STATE</type>
<position>447,-4066.5</position>
<input>
<ID>ENABLE_0</ID>941 </input>
<input>
<ID>IN_0</ID>942 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1384</ID>
<type>AA_AND2</type>
<position>591,-4068.5</position>
<input>
<ID>IN_0</ID>946 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1385</ID>
<type>AE_DFF_LOW</type>
<position>507,-4056.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>944 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1386</ID>
<type>BA_TRI_STATE</type>
<position>531.5,-4068.5</position>
<input>
<ID>ENABLE_0</ID>943 </input>
<input>
<ID>IN_0</ID>944 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1387</ID>
<type>AA_AND2</type>
<position>517,-4068.5</position>
<input>
<ID>IN_0</ID>944 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>943 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1388</ID>
<type>AE_DFF_LOW</type>
<position>580.5,-4056.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>946 </output>
<input>
<ID>clock</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1389</ID>
<type>BA_TRI_STATE</type>
<position>605,-4068.5</position>
<input>
<ID>ENABLE_0</ID>945 </input>
<input>
<ID>IN_0</ID>946 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1390</ID>
<type>AA_AND2</type>
<position>-5.5,-4057.5</position>
<input>
<ID>IN_0</ID>929 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>947 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1391</ID>
<type>BA_TRI_STATE</type>
<position>-27,-4076.5</position>
<input>
<ID>ENABLE_0</ID>929 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>930 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1392</ID>
<type>AA_AND2</type>
<position>107,-3973</position>
<input>
<ID>IN_0</ID>953 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>952 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1393</ID>
<type>AE_DFF_LOW</type>
<position>23,-3966.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>951 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1394</ID>
<type>BA_TRI_STATE</type>
<position>47.5,-3973</position>
<input>
<ID>ENABLE_0</ID>950 </input>
<input>
<ID>IN_0</ID>951 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1395</ID>
<type>AA_AND2</type>
<position>33,-3973</position>
<input>
<ID>IN_0</ID>951 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>950 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1396</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-3966.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>953 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1397</ID>
<type>BA_TRI_STATE</type>
<position>121,-3973</position>
<input>
<ID>ENABLE_0</ID>952 </input>
<input>
<ID>IN_0</ID>953 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1398</ID>
<type>AA_AND2</type>
<position>265,-3975</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>956 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1399</ID>
<type>AE_DFF_LOW</type>
<position>181,-3966.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>955 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1400</ID>
<type>BA_TRI_STATE</type>
<position>205.5,-3975</position>
<input>
<ID>ENABLE_0</ID>954 </input>
<input>
<ID>IN_0</ID>955 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1401</ID>
<type>AA_AND2</type>
<position>191,-3975</position>
<input>
<ID>IN_0</ID>955 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>954 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1402</ID>
<type>AE_DFF_LOW</type>
<position>255.5,-3966.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>957 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1403</ID>
<type>BA_TRI_STATE</type>
<position>279,-3975</position>
<input>
<ID>ENABLE_0</ID>956 </input>
<input>
<ID>IN_0</ID>957 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1404</ID>
<type>AA_AND2</type>
<position>430,-3976.5</position>
<input>
<ID>IN_0</ID>961 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>960 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1405</ID>
<type>AE_DFF_LOW</type>
<position>346,-3966.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>959 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1406</ID>
<type>BA_TRI_STATE</type>
<position>370.5,-3976.5</position>
<input>
<ID>ENABLE_0</ID>958 </input>
<input>
<ID>IN_0</ID>959 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1407</ID>
<type>AA_AND2</type>
<position>356,-3976.5</position>
<input>
<ID>IN_0</ID>959 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>958 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1408</ID>
<type>AE_DFF_LOW</type>
<position>419.5,-3966.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>961 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1409</ID>
<type>BA_TRI_STATE</type>
<position>444,-3976.5</position>
<input>
<ID>ENABLE_0</ID>960 </input>
<input>
<ID>IN_0</ID>961 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1410</ID>
<type>AA_AND2</type>
<position>588,-3978.5</position>
<input>
<ID>IN_0</ID>965 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>964 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1411</ID>
<type>AE_DFF_LOW</type>
<position>504,-3966.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>963 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1412</ID>
<type>BA_TRI_STATE</type>
<position>528.5,-3978.5</position>
<input>
<ID>ENABLE_0</ID>962 </input>
<input>
<ID>IN_0</ID>963 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1413</ID>
<type>AA_AND2</type>
<position>514,-3978.5</position>
<input>
<ID>IN_0</ID>963 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>962 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1414</ID>
<type>AE_DFF_LOW</type>
<position>577.5,-3966.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>965 </output>
<input>
<ID>clock</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1415</ID>
<type>BA_TRI_STATE</type>
<position>602,-3978.5</position>
<input>
<ID>ENABLE_0</ID>964 </input>
<input>
<ID>IN_0</ID>965 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1416</ID>
<type>AA_AND2</type>
<position>-8.5,-3967.5</position>
<input>
<ID>IN_0</ID>948 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>966 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1417</ID>
<type>BA_TRI_STATE</type>
<position>-30,-3986.5</position>
<input>
<ID>ENABLE_0</ID>948 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>949 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1418</ID>
<type>AA_AND2</type>
<position>114,-4231</position>
<input>
<ID>IN_0</ID>972 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>971 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1419</ID>
<type>AE_DFF_LOW</type>
<position>30,-4224.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>970 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1420</ID>
<type>BA_TRI_STATE</type>
<position>54.5,-4231</position>
<input>
<ID>ENABLE_0</ID>969 </input>
<input>
<ID>IN_0</ID>970 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1421</ID>
<type>AA_AND2</type>
<position>40,-4231</position>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>969 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1422</ID>
<type>AE_DFF_LOW</type>
<position>103.5,-4224.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>972 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1423</ID>
<type>BA_TRI_STATE</type>
<position>128,-4231</position>
<input>
<ID>ENABLE_0</ID>971 </input>
<input>
<ID>IN_0</ID>972 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1424</ID>
<type>AA_AND2</type>
<position>272,-4233</position>
<input>
<ID>IN_0</ID>976 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>975 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1425</ID>
<type>AE_DFF_LOW</type>
<position>188,-4224.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>974 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1426</ID>
<type>BA_TRI_STATE</type>
<position>212.5,-4233</position>
<input>
<ID>ENABLE_0</ID>973 </input>
<input>
<ID>IN_0</ID>974 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1427</ID>
<type>AA_AND2</type>
<position>198,-4233</position>
<input>
<ID>IN_0</ID>974 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>973 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1428</ID>
<type>AE_DFF_LOW</type>
<position>262.5,-4224.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>976 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1429</ID>
<type>BA_TRI_STATE</type>
<position>286,-4233</position>
<input>
<ID>ENABLE_0</ID>975 </input>
<input>
<ID>IN_0</ID>976 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1430</ID>
<type>AA_AND2</type>
<position>437,-4234.5</position>
<input>
<ID>IN_0</ID>980 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>979 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1431</ID>
<type>AE_DFF_LOW</type>
<position>353,-4224.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>978 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1432</ID>
<type>BA_TRI_STATE</type>
<position>377.5,-4234.5</position>
<input>
<ID>ENABLE_0</ID>977 </input>
<input>
<ID>IN_0</ID>978 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1433</ID>
<type>AA_AND2</type>
<position>363,-4234.5</position>
<input>
<ID>IN_0</ID>978 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>977 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1434</ID>
<type>AE_DFF_LOW</type>
<position>426.5,-4224.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>980 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1435</ID>
<type>BA_TRI_STATE</type>
<position>451,-4234.5</position>
<input>
<ID>ENABLE_0</ID>979 </input>
<input>
<ID>IN_0</ID>980 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1436</ID>
<type>AA_AND2</type>
<position>595,-4236.5</position>
<input>
<ID>IN_0</ID>984 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>983 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1437</ID>
<type>AE_DFF_LOW</type>
<position>511,-4224.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>982 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1438</ID>
<type>BA_TRI_STATE</type>
<position>535.5,-4236.5</position>
<input>
<ID>ENABLE_0</ID>981 </input>
<input>
<ID>IN_0</ID>982 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1439</ID>
<type>AA_AND2</type>
<position>521,-4236.5</position>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>968 </input>
<output>
<ID>OUT</ID>981 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1440</ID>
<type>AE_DFF_LOW</type>
<position>584.5,-4224.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>984 </output>
<input>
<ID>clock</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1441</ID>
<type>BA_TRI_STATE</type>
<position>609,-4236.5</position>
<input>
<ID>ENABLE_0</ID>983 </input>
<input>
<ID>IN_0</ID>984 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1442</ID>
<type>AA_AND2</type>
<position>-1.5,-4225.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>985 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1443</ID>
<type>BA_TRI_STATE</type>
<position>-23,-4244.5</position>
<input>
<ID>ENABLE_0</ID>967 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>968 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1444</ID>
<type>AA_AND2</type>
<position>111,-4141</position>
<input>
<ID>IN_0</ID>991 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>990 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1445</ID>
<type>AE_DFF_LOW</type>
<position>27,-4134.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>989 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1446</ID>
<type>BA_TRI_STATE</type>
<position>51.5,-4141</position>
<input>
<ID>ENABLE_0</ID>988 </input>
<input>
<ID>IN_0</ID>989 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1447</ID>
<type>AA_AND2</type>
<position>37,-4141</position>
<input>
<ID>IN_0</ID>989 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>988 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1448</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-4134.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>991 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1449</ID>
<type>BA_TRI_STATE</type>
<position>125,-4141</position>
<input>
<ID>ENABLE_0</ID>990 </input>
<input>
<ID>IN_0</ID>991 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1450</ID>
<type>AA_AND2</type>
<position>269,-4143</position>
<input>
<ID>IN_0</ID>995 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>994 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1451</ID>
<type>AE_DFF_LOW</type>
<position>185,-4134.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>993 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1452</ID>
<type>BA_TRI_STATE</type>
<position>209.5,-4143</position>
<input>
<ID>ENABLE_0</ID>992 </input>
<input>
<ID>IN_0</ID>993 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1453</ID>
<type>AA_AND2</type>
<position>195,-4143</position>
<input>
<ID>IN_0</ID>993 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>992 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1454</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-4134.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>995 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1455</ID>
<type>BA_TRI_STATE</type>
<position>283,-4143</position>
<input>
<ID>ENABLE_0</ID>994 </input>
<input>
<ID>IN_0</ID>995 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1456</ID>
<type>AA_AND2</type>
<position>434,-4144.5</position>
<input>
<ID>IN_0</ID>999 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>998 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1457</ID>
<type>AE_DFF_LOW</type>
<position>350,-4134.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>997 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1458</ID>
<type>BA_TRI_STATE</type>
<position>374.5,-4144.5</position>
<input>
<ID>ENABLE_0</ID>996 </input>
<input>
<ID>IN_0</ID>997 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1459</ID>
<type>AA_AND2</type>
<position>360,-4144.5</position>
<input>
<ID>IN_0</ID>997 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>996 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1460</ID>
<type>AE_DFF_LOW</type>
<position>423.5,-4134.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>999 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1461</ID>
<type>BA_TRI_STATE</type>
<position>448,-4144.5</position>
<input>
<ID>ENABLE_0</ID>998 </input>
<input>
<ID>IN_0</ID>999 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1462</ID>
<type>AA_AND2</type>
<position>592,-4146.5</position>
<input>
<ID>IN_0</ID>1003 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>1002 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1463</ID>
<type>AE_DFF_LOW</type>
<position>508,-4134.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1001 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1464</ID>
<type>BA_TRI_STATE</type>
<position>532.5,-4146.5</position>
<input>
<ID>ENABLE_0</ID>1000 </input>
<input>
<ID>IN_0</ID>1001 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1465</ID>
<type>AA_AND2</type>
<position>518,-4146.5</position>
<input>
<ID>IN_0</ID>1001 </input>
<input>
<ID>IN_1</ID>987 </input>
<output>
<ID>OUT</ID>1000 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1466</ID>
<type>AE_DFF_LOW</type>
<position>581.5,-4134.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1003 </output>
<input>
<ID>clock</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1467</ID>
<type>BA_TRI_STATE</type>
<position>606,-4146.5</position>
<input>
<ID>ENABLE_0</ID>1002 </input>
<input>
<ID>IN_0</ID>1003 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1468</ID>
<type>AA_AND2</type>
<position>-4.5,-4135.5</position>
<input>
<ID>IN_0</ID>986 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1004 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1469</ID>
<type>BA_TRI_STATE</type>
<position>-26,-4154.5</position>
<input>
<ID>ENABLE_0</ID>986 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>987 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1470</ID>
<type>AA_AND2</type>
<position>112,-4439</position>
<input>
<ID>IN_0</ID>1010 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1009 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1471</ID>
<type>AE_DFF_LOW</type>
<position>28,-4432.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1008 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1472</ID>
<type>BA_TRI_STATE</type>
<position>52.5,-4439</position>
<input>
<ID>ENABLE_0</ID>1007 </input>
<input>
<ID>IN_0</ID>1008 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1473</ID>
<type>AA_AND2</type>
<position>38,-4439</position>
<input>
<ID>IN_0</ID>1008 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1007 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1474</ID>
<type>AE_DFF_LOW</type>
<position>101.5,-4432.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1010 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1475</ID>
<type>BA_TRI_STATE</type>
<position>126,-4439</position>
<input>
<ID>ENABLE_0</ID>1009 </input>
<input>
<ID>IN_0</ID>1010 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1476</ID>
<type>AA_AND2</type>
<position>270,-4441</position>
<input>
<ID>IN_0</ID>1014 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1013 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1477</ID>
<type>AE_DFF_LOW</type>
<position>186,-4432.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1012 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1478</ID>
<type>BA_TRI_STATE</type>
<position>210.5,-4441</position>
<input>
<ID>ENABLE_0</ID>1011 </input>
<input>
<ID>IN_0</ID>1012 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1479</ID>
<type>AA_AND2</type>
<position>196,-4441</position>
<input>
<ID>IN_0</ID>1012 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1011 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1480</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-4432.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1014 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1481</ID>
<type>BA_TRI_STATE</type>
<position>284,-4441</position>
<input>
<ID>ENABLE_0</ID>1013 </input>
<input>
<ID>IN_0</ID>1014 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1482</ID>
<type>AA_AND2</type>
<position>435,-4442.5</position>
<input>
<ID>IN_0</ID>1018 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1017 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1483</ID>
<type>AE_DFF_LOW</type>
<position>351,-4432.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1016 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1484</ID>
<type>BA_TRI_STATE</type>
<position>375.5,-4442.5</position>
<input>
<ID>ENABLE_0</ID>1015 </input>
<input>
<ID>IN_0</ID>1016 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1485</ID>
<type>AA_AND2</type>
<position>361,-4442.5</position>
<input>
<ID>IN_0</ID>1016 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1015 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1486</ID>
<type>AE_DFF_LOW</type>
<position>424.5,-4432.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1018 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1487</ID>
<type>BA_TRI_STATE</type>
<position>449,-4442.5</position>
<input>
<ID>ENABLE_0</ID>1017 </input>
<input>
<ID>IN_0</ID>1018 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1488</ID>
<type>AA_AND2</type>
<position>593,-4444.5</position>
<input>
<ID>IN_0</ID>1022 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1021 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1489</ID>
<type>AE_DFF_LOW</type>
<position>509,-4432.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1020 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1490</ID>
<type>BA_TRI_STATE</type>
<position>533.5,-4444.5</position>
<input>
<ID>ENABLE_0</ID>1019 </input>
<input>
<ID>IN_0</ID>1020 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1491</ID>
<type>AA_AND2</type>
<position>519,-4444.5</position>
<input>
<ID>IN_0</ID>1020 </input>
<input>
<ID>IN_1</ID>1006 </input>
<output>
<ID>OUT</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1492</ID>
<type>AE_DFF_LOW</type>
<position>582.5,-4432.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1022 </output>
<input>
<ID>clock</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1493</ID>
<type>BA_TRI_STATE</type>
<position>607,-4444.5</position>
<input>
<ID>ENABLE_0</ID>1021 </input>
<input>
<ID>IN_0</ID>1022 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1494</ID>
<type>AA_AND2</type>
<position>-3.5,-4433.5</position>
<input>
<ID>IN_0</ID>1005 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1023 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1495</ID>
<type>BA_TRI_STATE</type>
<position>-25,-4452.5</position>
<input>
<ID>ENABLE_0</ID>1005 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1006 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1496</ID>
<type>AA_AND2</type>
<position>109,-4349</position>
<input>
<ID>IN_0</ID>1029 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1028 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1497</ID>
<type>AE_DFF_LOW</type>
<position>25,-4342.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1027 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1498</ID>
<type>BA_TRI_STATE</type>
<position>49.5,-4349</position>
<input>
<ID>ENABLE_0</ID>1026 </input>
<input>
<ID>IN_0</ID>1027 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1499</ID>
<type>AA_AND2</type>
<position>35,-4349</position>
<input>
<ID>IN_0</ID>1027 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1026 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1500</ID>
<type>AE_DFF_LOW</type>
<position>98.5,-4342.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1029 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1501</ID>
<type>BA_TRI_STATE</type>
<position>123,-4349</position>
<input>
<ID>ENABLE_0</ID>1028 </input>
<input>
<ID>IN_0</ID>1029 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1502</ID>
<type>AA_AND2</type>
<position>267,-4351</position>
<input>
<ID>IN_0</ID>1033 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1032 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1503</ID>
<type>AE_DFF_LOW</type>
<position>183,-4342.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1031 </output>
<input>
<ID>clock</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1504</ID>
<type>BA_TRI_STATE</type>
<position>207.5,-4351</position>
<input>
<ID>ENABLE_0</ID>1030 </input>
<input>
<ID>IN_0</ID>1031 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1505</ID>
<type>AA_AND2</type>
<position>190.5,-5275.5</position>
<input>
<ID>IN_0</ID>1183 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1182 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1506</ID>
<type>AE_DFF_LOW</type>
<position>255,-5267</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1185 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1507</ID>
<type>BA_TRI_STATE</type>
<position>278.5,-5275.5</position>
<input>
<ID>ENABLE_0</ID>1184 </input>
<input>
<ID>IN_0</ID>1185 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1508</ID>
<type>AA_AND2</type>
<position>429.5,-5277</position>
<input>
<ID>IN_0</ID>1189 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1509</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-5267</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1187 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1510</ID>
<type>BA_TRI_STATE</type>
<position>370,-5277</position>
<input>
<ID>ENABLE_0</ID>1186 </input>
<input>
<ID>IN_0</ID>1187 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1511</ID>
<type>AA_AND2</type>
<position>355.5,-5277</position>
<input>
<ID>IN_0</ID>1187 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1512</ID>
<type>AE_DFF_LOW</type>
<position>419,-5267</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1189 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1513</ID>
<type>BA_TRI_STATE</type>
<position>443.5,-5277</position>
<input>
<ID>ENABLE_0</ID>1188 </input>
<input>
<ID>IN_0</ID>1189 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1514</ID>
<type>AA_AND2</type>
<position>587.5,-5279</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1515</ID>
<type>AE_DFF_LOW</type>
<position>503.5,-5267</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1191 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1516</ID>
<type>BA_TRI_STATE</type>
<position>528,-5279</position>
<input>
<ID>ENABLE_0</ID>1190 </input>
<input>
<ID>IN_0</ID>1191 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1517</ID>
<type>AA_AND2</type>
<position>513.5,-5279</position>
<input>
<ID>IN_0</ID>1191 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1518</ID>
<type>AE_DFF_LOW</type>
<position>577,-5267</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1193 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1519</ID>
<type>BA_TRI_STATE</type>
<position>601.5,-5279</position>
<input>
<ID>ENABLE_0</ID>1192 </input>
<input>
<ID>IN_0</ID>1193 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1520</ID>
<type>AA_AND2</type>
<position>-9,-5268</position>
<input>
<ID>IN_0</ID>1176 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1521</ID>
<type>BA_TRI_STATE</type>
<position>-30.5,-5287</position>
<input>
<ID>ENABLE_0</ID>1176 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1177 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1522</ID>
<type>AA_AND2</type>
<position>113.5,-5531.5</position>
<input>
<ID>IN_0</ID>1200 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1523</ID>
<type>AE_DFF_LOW</type>
<position>29.5,-5525</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1198 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1524</ID>
<type>BA_TRI_STATE</type>
<position>54,-5531.5</position>
<input>
<ID>ENABLE_0</ID>1197 </input>
<input>
<ID>IN_0</ID>1198 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1525</ID>
<type>AA_AND2</type>
<position>39.5,-5531.5</position>
<input>
<ID>IN_0</ID>1198 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1526</ID>
<type>AE_DFF_LOW</type>
<position>103,-5525</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1200 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1527</ID>
<type>BA_TRI_STATE</type>
<position>127.5,-5531.5</position>
<input>
<ID>ENABLE_0</ID>1199 </input>
<input>
<ID>IN_0</ID>1200 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1528</ID>
<type>AA_AND2</type>
<position>271.5,-5533.5</position>
<input>
<ID>IN_0</ID>1204 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1529</ID>
<type>AE_DFF_LOW</type>
<position>187.5,-5525</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1202 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1530</ID>
<type>BA_TRI_STATE</type>
<position>212,-5533.5</position>
<input>
<ID>ENABLE_0</ID>1201 </input>
<input>
<ID>IN_0</ID>1202 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1531</ID>
<type>AA_AND2</type>
<position>197.5,-5533.5</position>
<input>
<ID>IN_0</ID>1202 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1532</ID>
<type>AE_DFF_LOW</type>
<position>262,-5525</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1204 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1533</ID>
<type>BA_TRI_STATE</type>
<position>285.5,-5533.5</position>
<input>
<ID>ENABLE_0</ID>1203 </input>
<input>
<ID>IN_0</ID>1204 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1534</ID>
<type>AA_AND2</type>
<position>436.5,-5535</position>
<input>
<ID>IN_0</ID>1208 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1535</ID>
<type>AE_DFF_LOW</type>
<position>352.5,-5525</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1206 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1536</ID>
<type>BA_TRI_STATE</type>
<position>377,-5535</position>
<input>
<ID>ENABLE_0</ID>1205 </input>
<input>
<ID>IN_0</ID>1206 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1537</ID>
<type>AA_AND2</type>
<position>362.5,-5535</position>
<input>
<ID>IN_0</ID>1206 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1538</ID>
<type>AE_DFF_LOW</type>
<position>426,-5525</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1208 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1539</ID>
<type>BA_TRI_STATE</type>
<position>450.5,-5535</position>
<input>
<ID>ENABLE_0</ID>1207 </input>
<input>
<ID>IN_0</ID>1208 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1540</ID>
<type>AA_AND2</type>
<position>594.5,-5537</position>
<input>
<ID>IN_0</ID>1212 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1541</ID>
<type>AE_DFF_LOW</type>
<position>510.5,-5525</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1210 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1542</ID>
<type>BA_TRI_STATE</type>
<position>535,-5537</position>
<input>
<ID>ENABLE_0</ID>1209 </input>
<input>
<ID>IN_0</ID>1210 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1543</ID>
<type>AA_AND2</type>
<position>520.5,-5537</position>
<input>
<ID>IN_0</ID>1210 </input>
<input>
<ID>IN_1</ID>1196 </input>
<output>
<ID>OUT</ID>1209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1544</ID>
<type>AE_DFF_LOW</type>
<position>584,-5525</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1212 </output>
<input>
<ID>clock</ID>1213 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1545</ID>
<type>BA_TRI_STATE</type>
<position>608.5,-5537</position>
<input>
<ID>ENABLE_0</ID>1211 </input>
<input>
<ID>IN_0</ID>1212 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1546</ID>
<type>AA_AND2</type>
<position>-2,-5526</position>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1547</ID>
<type>BA_TRI_STATE</type>
<position>-23.5,-5545</position>
<input>
<ID>ENABLE_0</ID>1195 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1196 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1548</ID>
<type>AA_AND2</type>
<position>110.5,-5441.5</position>
<input>
<ID>IN_0</ID>1219 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1549</ID>
<type>AE_DFF_LOW</type>
<position>26.5,-5435</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1217 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1550</ID>
<type>BA_TRI_STATE</type>
<position>51,-5441.5</position>
<input>
<ID>ENABLE_0</ID>1216 </input>
<input>
<ID>IN_0</ID>1217 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1551</ID>
<type>AA_AND2</type>
<position>36.5,-5441.5</position>
<input>
<ID>IN_0</ID>1217 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1552</ID>
<type>AE_DFF_LOW</type>
<position>100,-5435</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1219 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1553</ID>
<type>BA_TRI_STATE</type>
<position>124.5,-5441.5</position>
<input>
<ID>ENABLE_0</ID>1218 </input>
<input>
<ID>IN_0</ID>1219 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1554</ID>
<type>AA_AND2</type>
<position>268.5,-5443.5</position>
<input>
<ID>IN_0</ID>1223 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1555</ID>
<type>AE_DFF_LOW</type>
<position>184.5,-5435</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1221 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1556</ID>
<type>BA_TRI_STATE</type>
<position>209,-5443.5</position>
<input>
<ID>ENABLE_0</ID>1220 </input>
<input>
<ID>IN_0</ID>1221 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1557</ID>
<type>AA_AND2</type>
<position>194.5,-5443.5</position>
<input>
<ID>IN_0</ID>1221 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1558</ID>
<type>AE_DFF_LOW</type>
<position>259,-5435</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1223 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1559</ID>
<type>BA_TRI_STATE</type>
<position>282.5,-5443.5</position>
<input>
<ID>ENABLE_0</ID>1222 </input>
<input>
<ID>IN_0</ID>1223 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1560</ID>
<type>AA_AND2</type>
<position>433.5,-5445</position>
<input>
<ID>IN_0</ID>1227 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1561</ID>
<type>AE_DFF_LOW</type>
<position>349.5,-5435</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1225 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1562</ID>
<type>BA_TRI_STATE</type>
<position>374,-5445</position>
<input>
<ID>ENABLE_0</ID>1224 </input>
<input>
<ID>IN_0</ID>1225 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1563</ID>
<type>AA_AND2</type>
<position>359.5,-5445</position>
<input>
<ID>IN_0</ID>1225 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1564</ID>
<type>AE_DFF_LOW</type>
<position>423,-5435</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1227 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1565</ID>
<type>BA_TRI_STATE</type>
<position>447.5,-5445</position>
<input>
<ID>ENABLE_0</ID>1226 </input>
<input>
<ID>IN_0</ID>1227 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1566</ID>
<type>AA_AND2</type>
<position>591.5,-5447</position>
<input>
<ID>IN_0</ID>1231 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1567</ID>
<type>AE_DFF_LOW</type>
<position>507.5,-5435</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1229 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1568</ID>
<type>BA_TRI_STATE</type>
<position>532,-5447</position>
<input>
<ID>ENABLE_0</ID>1228 </input>
<input>
<ID>IN_0</ID>1229 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1569</ID>
<type>AA_AND2</type>
<position>517.5,-5447</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1215 </input>
<output>
<ID>OUT</ID>1228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1570</ID>
<type>AE_DFF_LOW</type>
<position>581,-5435</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1231 </output>
<input>
<ID>clock</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1571</ID>
<type>BA_TRI_STATE</type>
<position>605.5,-5447</position>
<input>
<ID>ENABLE_0</ID>1230 </input>
<input>
<ID>IN_0</ID>1231 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1572</ID>
<type>AA_AND2</type>
<position>-5,-5436</position>
<input>
<ID>IN_0</ID>1214 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1573</ID>
<type>BA_TRI_STATE</type>
<position>-26.5,-5455</position>
<input>
<ID>ENABLE_0</ID>1214 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1215 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1574</ID>
<type>BE_DECODER_3x8</type>
<position>-124,-5226.5</position>
<input>
<ID>ENABLE</ID>1399 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>1195 </output>
<output>
<ID>OUT_1</ID>1214 </output>
<output>
<ID>OUT_2</ID>1157 </output>
<output>
<ID>OUT_3</ID>1176 </output>
<output>
<ID>OUT_4</ID>1119 </output>
<output>
<ID>OUT_5</ID>1138 </output>
<output>
<ID>OUT_6</ID>1081 </output>
<output>
<ID>OUT_7</ID>1100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1575</ID>
<type>AA_AND2</type>
<position>107.5,-4987.5</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1085 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1576</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-4981</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1084 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1577</ID>
<type>BA_TRI_STATE</type>
<position>48,-4987.5</position>
<input>
<ID>ENABLE_0</ID>1083 </input>
<input>
<ID>IN_0</ID>1084 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1578</ID>
<type>AA_AND2</type>
<position>33.5,-4987.5</position>
<input>
<ID>IN_0</ID>1084 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1083 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1579</ID>
<type>AE_DFF_LOW</type>
<position>97,-4981</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1086 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1580</ID>
<type>BA_TRI_STATE</type>
<position>121.5,-4987.5</position>
<input>
<ID>ENABLE_0</ID>1085 </input>
<input>
<ID>IN_0</ID>1086 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1581</ID>
<type>AA_AND2</type>
<position>265.5,-4989.5</position>
<input>
<ID>IN_0</ID>1090 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1089 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1582</ID>
<type>AE_DFF_LOW</type>
<position>181.5,-4981</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1088 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1583</ID>
<type>BA_TRI_STATE</type>
<position>206,-4989.5</position>
<input>
<ID>ENABLE_0</ID>1087 </input>
<input>
<ID>IN_0</ID>1088 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1584</ID>
<type>AA_AND2</type>
<position>191.5,-4989.5</position>
<input>
<ID>IN_0</ID>1088 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1087 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1585</ID>
<type>AE_DFF_LOW</type>
<position>256,-4981</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1090 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1586</ID>
<type>BA_TRI_STATE</type>
<position>279.5,-4989.5</position>
<input>
<ID>ENABLE_0</ID>1089 </input>
<input>
<ID>IN_0</ID>1090 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1587</ID>
<type>AA_AND2</type>
<position>430.5,-4991</position>
<input>
<ID>IN_0</ID>1094 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1093 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1588</ID>
<type>AE_DFF_LOW</type>
<position>346.5,-4981</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1092 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1589</ID>
<type>BA_TRI_STATE</type>
<position>371,-4991</position>
<input>
<ID>ENABLE_0</ID>1091 </input>
<input>
<ID>IN_0</ID>1092 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1590</ID>
<type>AA_AND2</type>
<position>356.5,-4991</position>
<input>
<ID>IN_0</ID>1092 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1091 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1591</ID>
<type>AE_DFF_LOW</type>
<position>420,-4981</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1094 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1592</ID>
<type>BA_TRI_STATE</type>
<position>444.5,-4991</position>
<input>
<ID>ENABLE_0</ID>1093 </input>
<input>
<ID>IN_0</ID>1094 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1593</ID>
<type>AA_AND2</type>
<position>588.5,-4993</position>
<input>
<ID>IN_0</ID>1098 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1097 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1594</ID>
<type>AE_DFF_LOW</type>
<position>504.5,-4981</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1096 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1595</ID>
<type>BA_TRI_STATE</type>
<position>529,-4993</position>
<input>
<ID>ENABLE_0</ID>1095 </input>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1596</ID>
<type>AA_AND2</type>
<position>514.5,-4993</position>
<input>
<ID>IN_0</ID>1096 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1095 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1597</ID>
<type>AE_DFF_LOW</type>
<position>578,-4981</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1098 </output>
<input>
<ID>clock</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1598</ID>
<type>BA_TRI_STATE</type>
<position>602.5,-4993</position>
<input>
<ID>ENABLE_0</ID>1097 </input>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1599</ID>
<type>AA_AND2</type>
<position>-8,-4982</position>
<input>
<ID>IN_0</ID>1081 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1099 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1600</ID>
<type>BA_TRI_STATE</type>
<position>-29.5,-5001</position>
<input>
<ID>ENABLE_0</ID>1081 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1082 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1601</ID>
<type>AA_AND2</type>
<position>104.5,-4897.5</position>
<input>
<ID>IN_0</ID>1105 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1602</ID>
<type>AE_DFF_LOW</type>
<position>20.5,-4891</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1603</ID>
<type>BA_TRI_STATE</type>
<position>45,-4897.5</position>
<input>
<ID>ENABLE_0</ID>1102 </input>
<input>
<ID>IN_0</ID>1103 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1604</ID>
<type>AA_AND2</type>
<position>30.5,-4897.5</position>
<input>
<ID>IN_0</ID>1103 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1605</ID>
<type>AE_DFF_LOW</type>
<position>94,-4891</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1606</ID>
<type>BA_TRI_STATE</type>
<position>118.5,-4897.5</position>
<input>
<ID>ENABLE_0</ID>1104 </input>
<input>
<ID>IN_0</ID>1105 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1607</ID>
<type>AA_AND2</type>
<position>262.5,-4899.5</position>
<input>
<ID>IN_0</ID>1109 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1608</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-4891</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1107 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1609</ID>
<type>BA_TRI_STATE</type>
<position>203,-4899.5</position>
<input>
<ID>ENABLE_0</ID>1106 </input>
<input>
<ID>IN_0</ID>1107 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1610</ID>
<type>AA_AND2</type>
<position>188.5,-4899.5</position>
<input>
<ID>IN_0</ID>1107 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1611</ID>
<type>AE_DFF_LOW</type>
<position>253,-4891</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1109 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1612</ID>
<type>BA_TRI_STATE</type>
<position>276.5,-4899.5</position>
<input>
<ID>ENABLE_0</ID>1108 </input>
<input>
<ID>IN_0</ID>1109 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1613</ID>
<type>AA_AND2</type>
<position>427.5,-4901</position>
<input>
<ID>IN_0</ID>1113 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1614</ID>
<type>AE_DFF_LOW</type>
<position>343.5,-4891</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1111 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1615</ID>
<type>BA_TRI_STATE</type>
<position>368,-4901</position>
<input>
<ID>ENABLE_0</ID>1110 </input>
<input>
<ID>IN_0</ID>1111 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1616</ID>
<type>AA_AND2</type>
<position>353.5,-4901</position>
<input>
<ID>IN_0</ID>1111 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1617</ID>
<type>AE_DFF_LOW</type>
<position>417,-4891</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1113 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1618</ID>
<type>BA_TRI_STATE</type>
<position>441.5,-4901</position>
<input>
<ID>ENABLE_0</ID>1112 </input>
<input>
<ID>IN_0</ID>1113 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1619</ID>
<type>AA_AND2</type>
<position>585.5,-4903</position>
<input>
<ID>IN_0</ID>1117 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1620</ID>
<type>AE_DFF_LOW</type>
<position>501.5,-4891</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1115 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1621</ID>
<type>BA_TRI_STATE</type>
<position>526,-4903</position>
<input>
<ID>ENABLE_0</ID>1114 </input>
<input>
<ID>IN_0</ID>1115 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1622</ID>
<type>AA_AND2</type>
<position>511.5,-4903</position>
<input>
<ID>IN_0</ID>1115 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1623</ID>
<type>AE_DFF_LOW</type>
<position>575,-4891</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1117 </output>
<input>
<ID>clock</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1624</ID>
<type>BA_TRI_STATE</type>
<position>599.5,-4903</position>
<input>
<ID>ENABLE_0</ID>1116 </input>
<input>
<ID>IN_0</ID>1117 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1625</ID>
<type>AA_AND2</type>
<position>-11,-4892</position>
<input>
<ID>IN_0</ID>1100 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1626</ID>
<type>BA_TRI_STATE</type>
<position>-32.5,-4911</position>
<input>
<ID>ENABLE_0</ID>1100 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1101 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1627</ID>
<type>AA_AND2</type>
<position>111.5,-5155.5</position>
<input>
<ID>IN_0</ID>1124 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1628</ID>
<type>AE_DFF_LOW</type>
<position>27.5,-5149</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1122 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1629</ID>
<type>BA_TRI_STATE</type>
<position>52,-5155.5</position>
<input>
<ID>ENABLE_0</ID>1121 </input>
<input>
<ID>IN_0</ID>1122 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1630</ID>
<type>AA_AND2</type>
<position>37.5,-5155.5</position>
<input>
<ID>IN_0</ID>1122 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1631</ID>
<type>AE_DFF_LOW</type>
<position>101,-5149</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1124 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1632</ID>
<type>BA_TRI_STATE</type>
<position>125.5,-5155.5</position>
<input>
<ID>ENABLE_0</ID>1123 </input>
<input>
<ID>IN_0</ID>1124 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1633</ID>
<type>AA_AND2</type>
<position>269.5,-5157.5</position>
<input>
<ID>IN_0</ID>1128 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1634</ID>
<type>AE_DFF_LOW</type>
<position>185.5,-5149</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1126 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1635</ID>
<type>BA_TRI_STATE</type>
<position>210,-5157.5</position>
<input>
<ID>ENABLE_0</ID>1125 </input>
<input>
<ID>IN_0</ID>1126 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1636</ID>
<type>AA_AND2</type>
<position>195.5,-5157.5</position>
<input>
<ID>IN_0</ID>1126 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1637</ID>
<type>AE_DFF_LOW</type>
<position>260,-5149</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1128 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1638</ID>
<type>BA_TRI_STATE</type>
<position>283.5,-5157.5</position>
<input>
<ID>ENABLE_0</ID>1127 </input>
<input>
<ID>IN_0</ID>1128 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1639</ID>
<type>AA_AND2</type>
<position>434.5,-5159</position>
<input>
<ID>IN_0</ID>1132 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1640</ID>
<type>AE_DFF_LOW</type>
<position>350.5,-5149</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1130 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1641</ID>
<type>BA_TRI_STATE</type>
<position>375,-5159</position>
<input>
<ID>ENABLE_0</ID>1129 </input>
<input>
<ID>IN_0</ID>1130 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1642</ID>
<type>AA_AND2</type>
<position>360.5,-5159</position>
<input>
<ID>IN_0</ID>1130 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1643</ID>
<type>AE_DFF_LOW</type>
<position>424,-5149</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1132 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1644</ID>
<type>BA_TRI_STATE</type>
<position>448.5,-5159</position>
<input>
<ID>ENABLE_0</ID>1131 </input>
<input>
<ID>IN_0</ID>1132 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1645</ID>
<type>AA_AND2</type>
<position>592.5,-5161</position>
<input>
<ID>IN_0</ID>1136 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1646</ID>
<type>AE_DFF_LOW</type>
<position>508.5,-5149</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1134 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1647</ID>
<type>BA_TRI_STATE</type>
<position>533,-5161</position>
<input>
<ID>ENABLE_0</ID>1133 </input>
<input>
<ID>IN_0</ID>1134 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1648</ID>
<type>AA_AND2</type>
<position>518.5,-5161</position>
<input>
<ID>IN_0</ID>1134 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1649</ID>
<type>AE_DFF_LOW</type>
<position>582,-5149</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1136 </output>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1650</ID>
<type>BA_TRI_STATE</type>
<position>606.5,-5161</position>
<input>
<ID>ENABLE_0</ID>1135 </input>
<input>
<ID>IN_0</ID>1136 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1651</ID>
<type>AA_AND2</type>
<position>-4,-5150</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1652</ID>
<type>BA_TRI_STATE</type>
<position>-25.5,-5169</position>
<input>
<ID>ENABLE_0</ID>1119 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1120 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1653</ID>
<type>AA_AND2</type>
<position>108.5,-5065.5</position>
<input>
<ID>IN_0</ID>1143 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1654</ID>
<type>AE_DFF_LOW</type>
<position>24.5,-5059</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1657</ID>
<type>AE_DFF_LOW</type>
<position>98,-5059</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1143 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1658</ID>
<type>BA_TRI_STATE</type>
<position>122.5,-5065.5</position>
<input>
<ID>ENABLE_0</ID>1142 </input>
<input>
<ID>IN_0</ID>1143 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1659</ID>
<type>AA_AND2</type>
<position>266.5,-5067.5</position>
<input>
<ID>IN_0</ID>1147 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1660</ID>
<type>AE_DFF_LOW</type>
<position>182.5,-5059</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1145 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1661</ID>
<type>BA_TRI_STATE</type>
<position>207,-5067.5</position>
<input>
<ID>ENABLE_0</ID>1144 </input>
<input>
<ID>IN_0</ID>1145 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1662</ID>
<type>AA_AND2</type>
<position>192.5,-5067.5</position>
<input>
<ID>IN_0</ID>1145 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1663</ID>
<type>AE_DFF_LOW</type>
<position>257,-5059</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1147 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1664</ID>
<type>BA_TRI_STATE</type>
<position>280.5,-5067.5</position>
<input>
<ID>ENABLE_0</ID>1146 </input>
<input>
<ID>IN_0</ID>1147 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1665</ID>
<type>AA_AND2</type>
<position>431.5,-5069</position>
<input>
<ID>IN_0</ID>1151 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1666</ID>
<type>AE_DFF_LOW</type>
<position>347.5,-5059</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1149 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1667</ID>
<type>BA_TRI_STATE</type>
<position>372,-5069</position>
<input>
<ID>ENABLE_0</ID>1148 </input>
<input>
<ID>IN_0</ID>1149 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1668</ID>
<type>AA_AND2</type>
<position>357.5,-5069</position>
<input>
<ID>IN_0</ID>1149 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1669</ID>
<type>AE_DFF_LOW</type>
<position>421,-5059</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1151 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1670</ID>
<type>BA_TRI_STATE</type>
<position>445.5,-5069</position>
<input>
<ID>ENABLE_0</ID>1150 </input>
<input>
<ID>IN_0</ID>1151 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1671</ID>
<type>AA_AND2</type>
<position>589.5,-5071</position>
<input>
<ID>IN_0</ID>1155 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1672</ID>
<type>AE_DFF_LOW</type>
<position>505.5,-5059</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1153 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1673</ID>
<type>BA_TRI_STATE</type>
<position>530,-5071</position>
<input>
<ID>ENABLE_0</ID>1463 </input>
<input>
<ID>IN_0</ID>1153 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1674</ID>
<type>AA_AND2</type>
<position>515.5,-5071</position>
<input>
<ID>IN_0</ID>1153 </input>
<input>
<ID>IN_1</ID>1139 </input>
<output>
<ID>OUT</ID>1463 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1675</ID>
<type>AE_DFF_LOW</type>
<position>579,-5059</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1155 </output>
<input>
<ID>clock</ID>1156 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1676</ID>
<type>BA_TRI_STATE</type>
<position>603.5,-5071</position>
<input>
<ID>ENABLE_0</ID>1154 </input>
<input>
<ID>IN_0</ID>1155 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1677</ID>
<type>AA_AND2</type>
<position>-7,-5060</position>
<input>
<ID>IN_0</ID>1138 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1678</ID>
<type>BA_TRI_STATE</type>
<position>-28.5,-5079</position>
<input>
<ID>ENABLE_0</ID>1138 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1139 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1679</ID>
<type>AA_AND2</type>
<position>109.5,-5363.5</position>
<input>
<ID>IN_0</ID>1162 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1680</ID>
<type>AE_DFF_LOW</type>
<position>25.5,-5357</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1160 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1681</ID>
<type>BA_TRI_STATE</type>
<position>50,-5363.5</position>
<input>
<ID>ENABLE_0</ID>1159 </input>
<input>
<ID>IN_0</ID>1160 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1682</ID>
<type>AA_AND2</type>
<position>35.5,-5363.5</position>
<input>
<ID>IN_0</ID>1160 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1683</ID>
<type>AE_DFF_LOW</type>
<position>99,-5357</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1162 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1684</ID>
<type>BA_TRI_STATE</type>
<position>123.5,-5363.5</position>
<input>
<ID>ENABLE_0</ID>1161 </input>
<input>
<ID>IN_0</ID>1162 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1685</ID>
<type>AA_AND2</type>
<position>267.5,-5365.5</position>
<input>
<ID>IN_0</ID>1166 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1686</ID>
<type>AE_DFF_LOW</type>
<position>183.5,-5357</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1164 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1687</ID>
<type>BA_TRI_STATE</type>
<position>208,-5365.5</position>
<input>
<ID>ENABLE_0</ID>1163 </input>
<input>
<ID>IN_0</ID>1164 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1688</ID>
<type>AA_AND2</type>
<position>193.5,-5365.5</position>
<input>
<ID>IN_0</ID>1164 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1689</ID>
<type>AE_DFF_LOW</type>
<position>258,-5357</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1166 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1690</ID>
<type>BA_TRI_STATE</type>
<position>281.5,-5365.5</position>
<input>
<ID>ENABLE_0</ID>1165 </input>
<input>
<ID>IN_0</ID>1166 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1691</ID>
<type>AA_AND2</type>
<position>432.5,-5367</position>
<input>
<ID>IN_0</ID>1170 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1692</ID>
<type>AE_DFF_LOW</type>
<position>348.5,-5357</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1168 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1693</ID>
<type>BA_TRI_STATE</type>
<position>373,-5367</position>
<input>
<ID>ENABLE_0</ID>1167 </input>
<input>
<ID>IN_0</ID>1168 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1694</ID>
<type>AA_AND2</type>
<position>358.5,-5367</position>
<input>
<ID>IN_0</ID>1168 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1695</ID>
<type>AE_DFF_LOW</type>
<position>422,-5357</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1170 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1696</ID>
<type>BA_TRI_STATE</type>
<position>446.5,-5367</position>
<input>
<ID>ENABLE_0</ID>1169 </input>
<input>
<ID>IN_0</ID>1170 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1697</ID>
<type>AA_AND2</type>
<position>590.5,-5369</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1698</ID>
<type>AE_DFF_LOW</type>
<position>506.5,-5357</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1172 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1699</ID>
<type>BA_TRI_STATE</type>
<position>531,-5369</position>
<input>
<ID>ENABLE_0</ID>1171 </input>
<input>
<ID>IN_0</ID>1172 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1700</ID>
<type>AA_AND2</type>
<position>516.5,-5369</position>
<input>
<ID>IN_0</ID>1172 </input>
<input>
<ID>IN_1</ID>1158 </input>
<output>
<ID>OUT</ID>1171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1701</ID>
<type>AE_DFF_LOW</type>
<position>580,-5357</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1174 </output>
<input>
<ID>clock</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1702</ID>
<type>BA_TRI_STATE</type>
<position>604.5,-5369</position>
<input>
<ID>ENABLE_0</ID>1173 </input>
<input>
<ID>IN_0</ID>1174 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1703</ID>
<type>AA_AND2</type>
<position>-6,-5358</position>
<input>
<ID>IN_0</ID>1157 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1704</ID>
<type>BA_TRI_STATE</type>
<position>-27.5,-5377</position>
<input>
<ID>ENABLE_0</ID>1157 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1158 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1705</ID>
<type>AA_AND2</type>
<position>106.5,-5273.5</position>
<input>
<ID>IN_0</ID>1181 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1706</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-5267</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1179 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1707</ID>
<type>BA_TRI_STATE</type>
<position>47,-5273.5</position>
<input>
<ID>ENABLE_0</ID>1178 </input>
<input>
<ID>IN_0</ID>1179 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1708</ID>
<type>AA_AND2</type>
<position>32.5,-5273.5</position>
<input>
<ID>IN_0</ID>1179 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1709</ID>
<type>AE_DFF_LOW</type>
<position>96,-5267</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1181 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1710</ID>
<type>BA_TRI_STATE</type>
<position>120.5,-5273.5</position>
<input>
<ID>ENABLE_0</ID>1180 </input>
<input>
<ID>IN_0</ID>1181 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1711</ID>
<type>AA_AND2</type>
<position>264.5,-5275.5</position>
<input>
<ID>IN_0</ID>1185 </input>
<input>
<ID>IN_1</ID>1177 </input>
<output>
<ID>OUT</ID>1184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1712</ID>
<type>AE_DFF_LOW</type>
<position>180.5,-5267</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1183 </output>
<input>
<ID>clock</ID>1194 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1713</ID>
<type>BA_TRI_STATE</type>
<position>205,-5275.5</position>
<input>
<ID>ENABLE_0</ID>1182 </input>
<input>
<ID>IN_0</ID>1183 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1714</ID>
<type>AA_AND2</type>
<position>190,-6147</position>
<input>
<ID>IN_0</ID>1335 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1334 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1715</ID>
<type>AE_DFF_LOW</type>
<position>254.5,-6138.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1337 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1716</ID>
<type>BA_TRI_STATE</type>
<position>278,-6147</position>
<input>
<ID>ENABLE_0</ID>1336 </input>
<input>
<ID>IN_0</ID>1337 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1717</ID>
<type>AA_AND2</type>
<position>429,-6148.5</position>
<input>
<ID>IN_0</ID>1341 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1718</ID>
<type>AE_DFF_LOW</type>
<position>345,-6138.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1339 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1719</ID>
<type>BA_TRI_STATE</type>
<position>369.5,-6148.5</position>
<input>
<ID>ENABLE_0</ID>1338 </input>
<input>
<ID>IN_0</ID>1339 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1720</ID>
<type>AA_AND2</type>
<position>355,-6148.5</position>
<input>
<ID>IN_0</ID>1339 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1721</ID>
<type>AE_DFF_LOW</type>
<position>418.5,-6138.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1341 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1722</ID>
<type>BA_TRI_STATE</type>
<position>443,-6148.5</position>
<input>
<ID>ENABLE_0</ID>1340 </input>
<input>
<ID>IN_0</ID>1341 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1723</ID>
<type>AA_AND2</type>
<position>587,-6150.5</position>
<input>
<ID>IN_0</ID>1345 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1344 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1724</ID>
<type>AE_DFF_LOW</type>
<position>503,-6138.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1343 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1725</ID>
<type>BA_TRI_STATE</type>
<position>527.5,-6150.5</position>
<input>
<ID>ENABLE_0</ID>1342 </input>
<input>
<ID>IN_0</ID>1343 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1726</ID>
<type>AA_AND2</type>
<position>513,-6150.5</position>
<input>
<ID>IN_0</ID>1343 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1727</ID>
<type>AE_DFF_LOW</type>
<position>576.5,-6138.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1345 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1728</ID>
<type>BA_TRI_STATE</type>
<position>601,-6150.5</position>
<input>
<ID>ENABLE_0</ID>1344 </input>
<input>
<ID>IN_0</ID>1345 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1729</ID>
<type>AA_AND2</type>
<position>-9.5,-6139.5</position>
<input>
<ID>IN_0</ID>1328 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1346 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1730</ID>
<type>BA_TRI_STATE</type>
<position>-31,-6158.5</position>
<input>
<ID>ENABLE_0</ID>1328 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1329 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1731</ID>
<type>AA_AND2</type>
<position>113,-6403</position>
<input>
<ID>IN_0</ID>1352 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1351 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1732</ID>
<type>AE_DFF_LOW</type>
<position>29,-6396.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1350 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1733</ID>
<type>BA_TRI_STATE</type>
<position>53.5,-6403</position>
<input>
<ID>ENABLE_0</ID>1349 </input>
<input>
<ID>IN_0</ID>1350 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1734</ID>
<type>AA_AND2</type>
<position>39,-6403</position>
<input>
<ID>IN_0</ID>1350 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1349 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1735</ID>
<type>AE_DFF_LOW</type>
<position>102.5,-6396.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1352 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1736</ID>
<type>BA_TRI_STATE</type>
<position>127,-6403</position>
<input>
<ID>ENABLE_0</ID>1351 </input>
<input>
<ID>IN_0</ID>1352 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1737</ID>
<type>AA_AND2</type>
<position>271,-6405</position>
<input>
<ID>IN_0</ID>1356 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1738</ID>
<type>AE_DFF_LOW</type>
<position>187,-6396.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1354 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1739</ID>
<type>BA_TRI_STATE</type>
<position>211.5,-6405</position>
<input>
<ID>ENABLE_0</ID>1353 </input>
<input>
<ID>IN_0</ID>1354 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1740</ID>
<type>AA_AND2</type>
<position>197,-6405</position>
<input>
<ID>IN_0</ID>1354 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1353 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1741</ID>
<type>AE_DFF_LOW</type>
<position>261.5,-6396.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1356 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1742</ID>
<type>BA_TRI_STATE</type>
<position>285,-6405</position>
<input>
<ID>ENABLE_0</ID>1355 </input>
<input>
<ID>IN_0</ID>1356 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1743</ID>
<type>AA_AND2</type>
<position>436,-6406.5</position>
<input>
<ID>IN_0</ID>1360 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1359 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1744</ID>
<type>AE_DFF_LOW</type>
<position>352,-6396.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1358 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1745</ID>
<type>BA_TRI_STATE</type>
<position>376.5,-6406.5</position>
<input>
<ID>ENABLE_0</ID>1357 </input>
<input>
<ID>IN_0</ID>1358 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1746</ID>
<type>AA_AND2</type>
<position>362,-6406.5</position>
<input>
<ID>IN_0</ID>1358 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1357 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1747</ID>
<type>AE_DFF_LOW</type>
<position>425.5,-6396.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1360 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1748</ID>
<type>BA_TRI_STATE</type>
<position>450,-6406.5</position>
<input>
<ID>ENABLE_0</ID>1359 </input>
<input>
<ID>IN_0</ID>1360 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1749</ID>
<type>AA_AND2</type>
<position>594,-6408.5</position>
<input>
<ID>IN_0</ID>1364 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1363 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1750</ID>
<type>AE_DFF_LOW</type>
<position>510,-6396.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1362 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1751</ID>
<type>BA_TRI_STATE</type>
<position>534.5,-6408.5</position>
<input>
<ID>ENABLE_0</ID>1361 </input>
<input>
<ID>IN_0</ID>1362 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1752</ID>
<type>AA_AND2</type>
<position>520,-6408.5</position>
<input>
<ID>IN_0</ID>1362 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1361 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1753</ID>
<type>AE_DFF_LOW</type>
<position>583.5,-6396.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1364 </output>
<input>
<ID>clock</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1754</ID>
<type>BA_TRI_STATE</type>
<position>608,-6408.5</position>
<input>
<ID>ENABLE_0</ID>1363 </input>
<input>
<ID>IN_0</ID>1364 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1755</ID>
<type>AA_AND2</type>
<position>-2.5,-6397.5</position>
<input>
<ID>IN_0</ID>1347 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1365 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1756</ID>
<type>BA_TRI_STATE</type>
<position>-24,-6416.5</position>
<input>
<ID>ENABLE_0</ID>1347 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1348 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1757</ID>
<type>AA_AND2</type>
<position>110,-6313</position>
<input>
<ID>IN_0</ID>1371 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1758</ID>
<type>AE_DFF_LOW</type>
<position>26,-6306.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1369 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1759</ID>
<type>BA_TRI_STATE</type>
<position>50.5,-6313</position>
<input>
<ID>ENABLE_0</ID>1368 </input>
<input>
<ID>IN_0</ID>1369 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1760</ID>
<type>AA_AND2</type>
<position>36,-6313</position>
<input>
<ID>IN_0</ID>1369 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1368 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1761</ID>
<type>AE_DFF_LOW</type>
<position>99.5,-6306.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1371 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1762</ID>
<type>BA_TRI_STATE</type>
<position>124,-6313</position>
<input>
<ID>ENABLE_0</ID>1370 </input>
<input>
<ID>IN_0</ID>1371 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1763</ID>
<type>AA_AND2</type>
<position>268,-6315</position>
<input>
<ID>IN_0</ID>1375 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1764</ID>
<type>AE_DFF_LOW</type>
<position>184,-6306.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1373 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1765</ID>
<type>BA_TRI_STATE</type>
<position>208.5,-6315</position>
<input>
<ID>ENABLE_0</ID>1372 </input>
<input>
<ID>IN_0</ID>1373 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1766</ID>
<type>AA_AND2</type>
<position>194,-6315</position>
<input>
<ID>IN_0</ID>1373 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1372 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1767</ID>
<type>AE_DFF_LOW</type>
<position>258.5,-6306.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1375 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1768</ID>
<type>BA_TRI_STATE</type>
<position>282,-6315</position>
<input>
<ID>ENABLE_0</ID>1374 </input>
<input>
<ID>IN_0</ID>1375 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1769</ID>
<type>AA_AND2</type>
<position>433,-6316.5</position>
<input>
<ID>IN_0</ID>1379 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1378 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1770</ID>
<type>AE_DFF_LOW</type>
<position>349,-6306.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1377 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1771</ID>
<type>BA_TRI_STATE</type>
<position>373.5,-6316.5</position>
<input>
<ID>ENABLE_0</ID>1376 </input>
<input>
<ID>IN_0</ID>1377 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1772</ID>
<type>AA_AND2</type>
<position>359,-6316.5</position>
<input>
<ID>IN_0</ID>1377 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1376 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1773</ID>
<type>AE_DFF_LOW</type>
<position>422.5,-6306.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1379 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1774</ID>
<type>BA_TRI_STATE</type>
<position>447,-6316.5</position>
<input>
<ID>ENABLE_0</ID>1378 </input>
<input>
<ID>IN_0</ID>1379 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1775</ID>
<type>AA_AND2</type>
<position>591,-6318.5</position>
<input>
<ID>IN_0</ID>1383 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1776</ID>
<type>AE_DFF_LOW</type>
<position>507,-6306.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1381 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1777</ID>
<type>BA_TRI_STATE</type>
<position>531.5,-6318.5</position>
<input>
<ID>ENABLE_0</ID>1380 </input>
<input>
<ID>IN_0</ID>1381 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1778</ID>
<type>AA_AND2</type>
<position>517,-6318.5</position>
<input>
<ID>IN_0</ID>1381 </input>
<input>
<ID>IN_1</ID>1367 </input>
<output>
<ID>OUT</ID>1380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1779</ID>
<type>AE_DFF_LOW</type>
<position>580.5,-6306.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1383 </output>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1780</ID>
<type>BA_TRI_STATE</type>
<position>605,-6318.5</position>
<input>
<ID>ENABLE_0</ID>1382 </input>
<input>
<ID>IN_0</ID>1383 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1781</ID>
<type>AA_AND2</type>
<position>-5.5,-6307.5</position>
<input>
<ID>IN_0</ID>1366 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1384 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1782</ID>
<type>BA_TRI_STATE</type>
<position>-27,-6326.5</position>
<input>
<ID>ENABLE_0</ID>1366 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1367 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1783</ID>
<type>BE_DECODER_3x8</type>
<position>-124.5,-6098</position>
<input>
<ID>ENABLE</ID>1400 </input>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1386 </input>
<input>
<ID>IN_2</ID>1385 </input>
<output>
<ID>OUT_0</ID>1347 </output>
<output>
<ID>OUT_1</ID>1366 </output>
<output>
<ID>OUT_2</ID>1309 </output>
<output>
<ID>OUT_3</ID>1328 </output>
<output>
<ID>OUT_4</ID>1271 </output>
<output>
<ID>OUT_5</ID>1290 </output>
<output>
<ID>OUT_6</ID>1233 </output>
<output>
<ID>OUT_7</ID>1252 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1784</ID>
<type>AA_AND2</type>
<position>107,-5859</position>
<input>
<ID>IN_0</ID>1238 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1785</ID>
<type>AE_DFF_LOW</type>
<position>23,-5852.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1236 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1786</ID>
<type>BA_TRI_STATE</type>
<position>47.5,-5859</position>
<input>
<ID>ENABLE_0</ID>1235 </input>
<input>
<ID>IN_0</ID>1236 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1787</ID>
<type>AA_AND2</type>
<position>33,-5859</position>
<input>
<ID>IN_0</ID>1236 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1788</ID>
<type>AE_DFF_LOW</type>
<position>96.5,-5852.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1238 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1789</ID>
<type>BA_TRI_STATE</type>
<position>121,-5859</position>
<input>
<ID>ENABLE_0</ID>1237 </input>
<input>
<ID>IN_0</ID>1238 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1790</ID>
<type>AA_AND2</type>
<position>265,-5861</position>
<input>
<ID>IN_0</ID>1242 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1791</ID>
<type>AE_DFF_LOW</type>
<position>181,-5852.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1240 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1792</ID>
<type>BA_TRI_STATE</type>
<position>205.5,-5861</position>
<input>
<ID>ENABLE_0</ID>1239 </input>
<input>
<ID>IN_0</ID>1240 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1793</ID>
<type>AA_AND2</type>
<position>191,-5861</position>
<input>
<ID>IN_0</ID>1240 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1794</ID>
<type>AE_DFF_LOW</type>
<position>255.5,-5852.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1242 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1795</ID>
<type>BA_TRI_STATE</type>
<position>279,-5861</position>
<input>
<ID>ENABLE_0</ID>1241 </input>
<input>
<ID>IN_0</ID>1242 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1796</ID>
<type>AA_AND2</type>
<position>430,-5862.5</position>
<input>
<ID>IN_0</ID>1246 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1797</ID>
<type>AE_DFF_LOW</type>
<position>346,-5852.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1244 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1798</ID>
<type>BA_TRI_STATE</type>
<position>370.5,-5862.5</position>
<input>
<ID>ENABLE_0</ID>1243 </input>
<input>
<ID>IN_0</ID>1244 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1799</ID>
<type>AA_AND2</type>
<position>356,-5862.5</position>
<input>
<ID>IN_0</ID>1244 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1800</ID>
<type>AE_DFF_LOW</type>
<position>419.5,-5852.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1246 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1801</ID>
<type>BA_TRI_STATE</type>
<position>444,-5862.5</position>
<input>
<ID>ENABLE_0</ID>1245 </input>
<input>
<ID>IN_0</ID>1246 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1802</ID>
<type>AA_AND2</type>
<position>588,-5864.5</position>
<input>
<ID>IN_0</ID>1250 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1803</ID>
<type>AE_DFF_LOW</type>
<position>504,-5852.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1248 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1804</ID>
<type>BA_TRI_STATE</type>
<position>528.5,-5864.5</position>
<input>
<ID>ENABLE_0</ID>1247 </input>
<input>
<ID>IN_0</ID>1248 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1805</ID>
<type>AA_AND2</type>
<position>514,-5864.5</position>
<input>
<ID>IN_0</ID>1248 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1806</ID>
<type>AE_DFF_LOW</type>
<position>577.5,-5852.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1250 </output>
<input>
<ID>clock</ID>1251 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1807</ID>
<type>BA_TRI_STATE</type>
<position>602,-5864.5</position>
<input>
<ID>ENABLE_0</ID>1249 </input>
<input>
<ID>IN_0</ID>1250 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1808</ID>
<type>AA_AND2</type>
<position>-8.5,-5853.5</position>
<input>
<ID>IN_0</ID>1233 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1809</ID>
<type>BA_TRI_STATE</type>
<position>-30,-5872.5</position>
<input>
<ID>ENABLE_0</ID>1233 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1234 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1810</ID>
<type>AA_AND2</type>
<position>104,-5769</position>
<input>
<ID>IN_0</ID>1257 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1256 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1811</ID>
<type>AE_DFF_LOW</type>
<position>20,-5762.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1255 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1812</ID>
<type>BA_TRI_STATE</type>
<position>44.5,-5769</position>
<input>
<ID>ENABLE_0</ID>1254 </input>
<input>
<ID>IN_0</ID>1255 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1813</ID>
<type>AA_AND2</type>
<position>30,-5769</position>
<input>
<ID>IN_0</ID>1255 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1814</ID>
<type>AE_DFF_LOW</type>
<position>93.5,-5762.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1257 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1815</ID>
<type>BA_TRI_STATE</type>
<position>118,-5769</position>
<input>
<ID>ENABLE_0</ID>1256 </input>
<input>
<ID>IN_0</ID>1257 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1816</ID>
<type>AA_AND2</type>
<position>262,-5771</position>
<input>
<ID>IN_0</ID>1261 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1817</ID>
<type>AE_DFF_LOW</type>
<position>178,-5762.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1259 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1818</ID>
<type>BA_TRI_STATE</type>
<position>202.5,-5771</position>
<input>
<ID>ENABLE_0</ID>1258 </input>
<input>
<ID>IN_0</ID>1259 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1819</ID>
<type>AA_AND2</type>
<position>188,-5771</position>
<input>
<ID>IN_0</ID>1259 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1258 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1820</ID>
<type>AE_DFF_LOW</type>
<position>252.5,-5762.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1261 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1821</ID>
<type>BA_TRI_STATE</type>
<position>276,-5771</position>
<input>
<ID>ENABLE_0</ID>1260 </input>
<input>
<ID>IN_0</ID>1261 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1822</ID>
<type>AA_AND2</type>
<position>427,-5772.5</position>
<input>
<ID>IN_0</ID>1265 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1264 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1823</ID>
<type>AE_DFF_LOW</type>
<position>343,-5762.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1263 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1824</ID>
<type>BA_TRI_STATE</type>
<position>367.5,-5772.5</position>
<input>
<ID>ENABLE_0</ID>1262 </input>
<input>
<ID>IN_0</ID>1263 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1825</ID>
<type>AA_AND2</type>
<position>353,-5772.5</position>
<input>
<ID>IN_0</ID>1263 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1826</ID>
<type>AE_DFF_LOW</type>
<position>416.5,-5762.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1265 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1827</ID>
<type>BA_TRI_STATE</type>
<position>441,-5772.5</position>
<input>
<ID>ENABLE_0</ID>1264 </input>
<input>
<ID>IN_0</ID>1265 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1828</ID>
<type>AA_AND2</type>
<position>585,-5774.5</position>
<input>
<ID>IN_0</ID>1269 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1829</ID>
<type>AE_DFF_LOW</type>
<position>501,-5762.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1267 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1830</ID>
<type>BA_TRI_STATE</type>
<position>525.5,-5774.5</position>
<input>
<ID>ENABLE_0</ID>1266 </input>
<input>
<ID>IN_0</ID>1267 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1831</ID>
<type>AA_AND2</type>
<position>511,-5774.5</position>
<input>
<ID>IN_0</ID>1267 </input>
<input>
<ID>IN_1</ID>1253 </input>
<output>
<ID>OUT</ID>1266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1832</ID>
<type>AE_DFF_LOW</type>
<position>574.5,-5762.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1269 </output>
<input>
<ID>clock</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1833</ID>
<type>BA_TRI_STATE</type>
<position>599,-5774.5</position>
<input>
<ID>ENABLE_0</ID>1268 </input>
<input>
<ID>IN_0</ID>1269 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1834</ID>
<type>AA_AND2</type>
<position>-11.5,-5763.5</position>
<input>
<ID>IN_0</ID>1252 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1835</ID>
<type>BA_TRI_STATE</type>
<position>-33,-5782.5</position>
<input>
<ID>ENABLE_0</ID>1252 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1253 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1836</ID>
<type>AA_AND2</type>
<position>111,-6027</position>
<input>
<ID>IN_0</ID>1276 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1837</ID>
<type>AE_DFF_LOW</type>
<position>27,-6020.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1274 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1838</ID>
<type>BA_TRI_STATE</type>
<position>51.5,-6027</position>
<input>
<ID>ENABLE_0</ID>1273 </input>
<input>
<ID>IN_0</ID>1274 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1839</ID>
<type>AA_AND2</type>
<position>37,-6027</position>
<input>
<ID>IN_0</ID>1274 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1840</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-6020.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1276 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1841</ID>
<type>BA_TRI_STATE</type>
<position>125,-6027</position>
<input>
<ID>ENABLE_0</ID>1275 </input>
<input>
<ID>IN_0</ID>1276 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1842</ID>
<type>AA_AND2</type>
<position>269,-6029</position>
<input>
<ID>IN_0</ID>1280 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1279 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1843</ID>
<type>AE_DFF_LOW</type>
<position>185,-6020.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1278 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1844</ID>
<type>BA_TRI_STATE</type>
<position>209.5,-6029</position>
<input>
<ID>ENABLE_0</ID>1277 </input>
<input>
<ID>IN_0</ID>1278 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1845</ID>
<type>AA_AND2</type>
<position>195,-6029</position>
<input>
<ID>IN_0</ID>1278 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1846</ID>
<type>AE_DFF_LOW</type>
<position>259.5,-6020.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1280 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1847</ID>
<type>BA_TRI_STATE</type>
<position>283,-6029</position>
<input>
<ID>ENABLE_0</ID>1279 </input>
<input>
<ID>IN_0</ID>1280 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1848</ID>
<type>AA_AND2</type>
<position>434,-6030.5</position>
<input>
<ID>IN_0</ID>1284 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1849</ID>
<type>AE_DFF_LOW</type>
<position>350,-6020.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1282 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1850</ID>
<type>BA_TRI_STATE</type>
<position>374.5,-6030.5</position>
<input>
<ID>ENABLE_0</ID>1281 </input>
<input>
<ID>IN_0</ID>1282 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1851</ID>
<type>AA_AND2</type>
<position>360,-6030.5</position>
<input>
<ID>IN_0</ID>1282 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1852</ID>
<type>AE_DFF_LOW</type>
<position>423.5,-6020.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1284 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1853</ID>
<type>BA_TRI_STATE</type>
<position>448,-6030.5</position>
<input>
<ID>ENABLE_0</ID>1283 </input>
<input>
<ID>IN_0</ID>1284 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1854</ID>
<type>AA_AND2</type>
<position>592,-6032.5</position>
<input>
<ID>IN_0</ID>1288 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1855</ID>
<type>AE_DFF_LOW</type>
<position>508,-6020.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1286 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1856</ID>
<type>BA_TRI_STATE</type>
<position>532.5,-6032.5</position>
<input>
<ID>ENABLE_0</ID>1285 </input>
<input>
<ID>IN_0</ID>1286 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1857</ID>
<type>AA_AND2</type>
<position>518,-6032.5</position>
<input>
<ID>IN_0</ID>1286 </input>
<input>
<ID>IN_1</ID>1272 </input>
<output>
<ID>OUT</ID>1285 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1858</ID>
<type>AE_DFF_LOW</type>
<position>581.5,-6020.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1288 </output>
<input>
<ID>clock</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1859</ID>
<type>BA_TRI_STATE</type>
<position>606,-6032.5</position>
<input>
<ID>ENABLE_0</ID>1287 </input>
<input>
<ID>IN_0</ID>1288 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1860</ID>
<type>AA_AND2</type>
<position>-4.5,-6021.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1289 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1861</ID>
<type>BA_TRI_STATE</type>
<position>-26,-6040.5</position>
<input>
<ID>ENABLE_0</ID>1271 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1272 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1862</ID>
<type>AA_AND2</type>
<position>108,-5937</position>
<input>
<ID>IN_0</ID>1295 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1294 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1863</ID>
<type>AE_DFF_LOW</type>
<position>24,-5930.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1293 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1864</ID>
<type>BA_TRI_STATE</type>
<position>48.5,-5937</position>
<input>
<ID>ENABLE_0</ID>1292 </input>
<input>
<ID>IN_0</ID>1293 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1865</ID>
<type>AA_AND2</type>
<position>34,-5937</position>
<input>
<ID>IN_0</ID>1293 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1292 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1866</ID>
<type>AE_DFF_LOW</type>
<position>97.5,-5930.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1295 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1867</ID>
<type>BA_TRI_STATE</type>
<position>122,-5937</position>
<input>
<ID>ENABLE_0</ID>1294 </input>
<input>
<ID>IN_0</ID>1295 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1868</ID>
<type>AA_AND2</type>
<position>266,-5939</position>
<input>
<ID>IN_0</ID>1299 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1298 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1869</ID>
<type>AE_DFF_LOW</type>
<position>182,-5930.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1297 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1870</ID>
<type>BA_TRI_STATE</type>
<position>206.5,-5939</position>
<input>
<ID>ENABLE_0</ID>1296 </input>
<input>
<ID>IN_0</ID>1297 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1871</ID>
<type>AA_AND2</type>
<position>192,-5939</position>
<input>
<ID>IN_0</ID>1297 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1296 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1872</ID>
<type>AE_DFF_LOW</type>
<position>256.5,-5930.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1299 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1873</ID>
<type>BA_TRI_STATE</type>
<position>280,-5939</position>
<input>
<ID>ENABLE_0</ID>1298 </input>
<input>
<ID>IN_0</ID>1299 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1874</ID>
<type>AA_AND2</type>
<position>431,-5940.5</position>
<input>
<ID>IN_0</ID>1303 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1302 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1875</ID>
<type>AE_DFF_LOW</type>
<position>347,-5930.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1301 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1876</ID>
<type>BA_TRI_STATE</type>
<position>371.5,-5940.5</position>
<input>
<ID>ENABLE_0</ID>1300 </input>
<input>
<ID>IN_0</ID>1301 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1877</ID>
<type>AA_AND2</type>
<position>357,-5940.5</position>
<input>
<ID>IN_0</ID>1301 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1300 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1878</ID>
<type>AE_DFF_LOW</type>
<position>420.5,-5930.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1303 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1879</ID>
<type>BA_TRI_STATE</type>
<position>445,-5940.5</position>
<input>
<ID>ENABLE_0</ID>1302 </input>
<input>
<ID>IN_0</ID>1303 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1880</ID>
<type>AA_AND2</type>
<position>589,-5942.5</position>
<input>
<ID>IN_0</ID>1307 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1306 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1881</ID>
<type>AE_DFF_LOW</type>
<position>505,-5930.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1305 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1882</ID>
<type>BA_TRI_STATE</type>
<position>529.5,-5942.5</position>
<input>
<ID>ENABLE_0</ID>1304 </input>
<input>
<ID>IN_0</ID>1305 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1883</ID>
<type>AA_AND2</type>
<position>515,-5942.5</position>
<input>
<ID>IN_0</ID>1305 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1304 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1884</ID>
<type>AE_DFF_LOW</type>
<position>578.5,-5930.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1307 </output>
<input>
<ID>clock</ID>1308 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1885</ID>
<type>BA_TRI_STATE</type>
<position>603,-5942.5</position>
<input>
<ID>ENABLE_0</ID>1306 </input>
<input>
<ID>IN_0</ID>1307 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1886</ID>
<type>AA_AND2</type>
<position>-7.5,-5931.5</position>
<input>
<ID>IN_0</ID>1290 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1887</ID>
<type>BA_TRI_STATE</type>
<position>-29,-5950.5</position>
<input>
<ID>ENABLE_0</ID>1290 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1291 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1888</ID>
<type>AA_AND2</type>
<position>109,-6235</position>
<input>
<ID>IN_0</ID>1314 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1313 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1889</ID>
<type>AE_DFF_LOW</type>
<position>25,-6228.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1312 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1890</ID>
<type>BA_TRI_STATE</type>
<position>49.5,-6235</position>
<input>
<ID>ENABLE_0</ID>1311 </input>
<input>
<ID>IN_0</ID>1312 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1891</ID>
<type>AA_AND2</type>
<position>35,-6235</position>
<input>
<ID>IN_0</ID>1312 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1311 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1892</ID>
<type>AE_DFF_LOW</type>
<position>98.5,-6228.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1314 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1893</ID>
<type>BA_TRI_STATE</type>
<position>123,-6235</position>
<input>
<ID>ENABLE_0</ID>1313 </input>
<input>
<ID>IN_0</ID>1314 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1894</ID>
<type>AA_AND2</type>
<position>267,-6237</position>
<input>
<ID>IN_0</ID>1318 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1317 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1895</ID>
<type>AE_DFF_LOW</type>
<position>183,-6228.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1316 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1896</ID>
<type>BA_TRI_STATE</type>
<position>207.5,-6237</position>
<input>
<ID>ENABLE_0</ID>1315 </input>
<input>
<ID>IN_0</ID>1316 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1897</ID>
<type>AA_AND2</type>
<position>193,-6237</position>
<input>
<ID>IN_0</ID>1316 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1315 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1898</ID>
<type>AE_DFF_LOW</type>
<position>257.5,-6228.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<output>
<ID>OUT_0</ID>1318 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1899</ID>
<type>BA_TRI_STATE</type>
<position>281,-6237</position>
<input>
<ID>ENABLE_0</ID>1317 </input>
<input>
<ID>IN_0</ID>1318 </input>
<output>
<ID>OUT_0</ID>1460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1900</ID>
<type>AA_AND2</type>
<position>432,-6238.5</position>
<input>
<ID>IN_0</ID>1322 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1321 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1901</ID>
<type>AE_DFF_LOW</type>
<position>348,-6228.5</position>
<input>
<ID>IN_0</ID>1469 </input>
<output>
<ID>OUT_0</ID>1320 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1902</ID>
<type>BA_TRI_STATE</type>
<position>372.5,-6238.5</position>
<input>
<ID>ENABLE_0</ID>1319 </input>
<input>
<ID>IN_0</ID>1320 </input>
<output>
<ID>OUT_0</ID>1461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1903</ID>
<type>AA_AND2</type>
<position>358,-6238.5</position>
<input>
<ID>IN_0</ID>1320 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1319 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1904</ID>
<type>AE_DFF_LOW</type>
<position>421.5,-6228.5</position>
<input>
<ID>IN_0</ID>1470 </input>
<output>
<ID>OUT_0</ID>1322 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1905</ID>
<type>BA_TRI_STATE</type>
<position>446,-6238.5</position>
<input>
<ID>ENABLE_0</ID>1321 </input>
<input>
<ID>IN_0</ID>1322 </input>
<output>
<ID>OUT_0</ID>1462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1906</ID>
<type>AA_AND2</type>
<position>590,-6240.5</position>
<input>
<ID>IN_0</ID>1326 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1907</ID>
<type>AE_DFF_LOW</type>
<position>506,-6228.5</position>
<input>
<ID>IN_0</ID>1471 </input>
<output>
<ID>OUT_0</ID>1324 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1908</ID>
<type>BA_TRI_STATE</type>
<position>530.5,-6240.5</position>
<input>
<ID>ENABLE_0</ID>1323 </input>
<input>
<ID>IN_0</ID>1324 </input>
<output>
<ID>OUT_0</ID>1463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1909</ID>
<type>AA_AND2</type>
<position>516,-6240.5</position>
<input>
<ID>IN_0</ID>1324 </input>
<input>
<ID>IN_1</ID>1310 </input>
<output>
<ID>OUT</ID>1323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1910</ID>
<type>AE_DFF_LOW</type>
<position>579.5,-6228.5</position>
<input>
<ID>IN_0</ID>1472 </input>
<output>
<ID>OUT_0</ID>1326 </output>
<input>
<ID>clock</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1911</ID>
<type>BA_TRI_STATE</type>
<position>604,-6240.5</position>
<input>
<ID>ENABLE_0</ID>1325 </input>
<input>
<ID>IN_0</ID>1326 </input>
<output>
<ID>OUT_0</ID>1464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1912</ID>
<type>AA_AND2</type>
<position>-6.5,-6229.5</position>
<input>
<ID>IN_0</ID>1309 </input>
<input>
<ID>IN_1</ID>1423 </input>
<output>
<ID>OUT</ID>1327 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1913</ID>
<type>BA_TRI_STATE</type>
<position>-28,-6248.5</position>
<input>
<ID>ENABLE_0</ID>1309 </input>
<input>
<ID>IN_0</ID>1456 </input>
<output>
<ID>OUT_0</ID>1310 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1914</ID>
<type>AA_AND2</type>
<position>106,-6145</position>
<input>
<ID>IN_0</ID>1333 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1332 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1915</ID>
<type>AE_DFF_LOW</type>
<position>22,-6138.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<output>
<ID>OUT_0</ID>1331 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1916</ID>
<type>BA_TRI_STATE</type>
<position>46.5,-6145</position>
<input>
<ID>ENABLE_0</ID>1330 </input>
<input>
<ID>IN_0</ID>1331 </input>
<output>
<ID>OUT_0</ID>1457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1917</ID>
<type>AA_AND2</type>
<position>32,-6145</position>
<input>
<ID>IN_0</ID>1331 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1330 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1918</ID>
<type>AE_DFF_LOW</type>
<position>95.5,-6138.5</position>
<input>
<ID>IN_0</ID>1466 </input>
<output>
<ID>OUT_0</ID>1333 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1919</ID>
<type>BA_TRI_STATE</type>
<position>120,-6145</position>
<input>
<ID>ENABLE_0</ID>1332 </input>
<input>
<ID>IN_0</ID>1333 </input>
<output>
<ID>OUT_0</ID>1458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1920</ID>
<type>AA_AND2</type>
<position>264,-6147</position>
<input>
<ID>IN_0</ID>1337 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1336 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1921</ID>
<type>AE_DFF_LOW</type>
<position>180,-6138.5</position>
<input>
<ID>IN_0</ID>1467 </input>
<output>
<ID>OUT_0</ID>1335 </output>
<input>
<ID>clock</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1922</ID>
<type>BA_TRI_STATE</type>
<position>204.5,-6147</position>
<input>
<ID>ENABLE_0</ID>1334 </input>
<input>
<ID>IN_0</ID>1335 </input>
<output>
<ID>OUT_0</ID>1459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1926</ID>
<type>AA_TOGGLE</type>
<position>-172,42</position>
<output>
<ID>OUT_0</ID>1385 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1928</ID>
<type>AA_TOGGLE</type>
<position>-172,36.5</position>
<output>
<ID>OUT_0</ID>1386 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1930</ID>
<type>AA_TOGGLE</type>
<position>-172,30</position>
<output>
<ID>OUT_0</ID>1387 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1935</ID>
<type>BE_DECODER_3x8</type>
<position>-144,22.5</position>
<input>
<ID>ENABLE</ID>1392 </input>
<input>
<ID>IN_0</ID>1391 </input>
<input>
<ID>IN_1</ID>1390 </input>
<input>
<ID>IN_2</ID>1389 </input>
<output>
<ID>OUT_0</ID>1400 </output>
<output>
<ID>OUT_1</ID>1399 </output>
<output>
<ID>OUT_2</ID>1398 </output>
<output>
<ID>OUT_3</ID>1397 </output>
<output>
<ID>OUT_4</ID>1396 </output>
<output>
<ID>OUT_5</ID>1395 </output>
<output>
<ID>OUT_6</ID>1394 </output>
<output>
<ID>OUT_7</ID>1393 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1937</ID>
<type>AA_TOGGLE</type>
<position>-172,21</position>
<output>
<ID>OUT_0</ID>1389 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1939</ID>
<type>AA_TOGGLE</type>
<position>-172.5,16.5</position>
<output>
<ID>OUT_0</ID>1390 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1941</ID>
<type>AA_TOGGLE</type>
<position>-172,12</position>
<output>
<ID>OUT_0</ID>1391 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1943</ID>
<type>AA_TOGGLE</type>
<position>-152.5,26</position>
<output>
<ID>OUT_0</ID>1392 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1945</ID>
<type>AA_LABEL</type>
<position>-156,27</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1947</ID>
<type>AA_LABEL</type>
<position>-178,42.5</position>
<gparam>LABEL_TEXT i/p 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1948</ID>
<type>AA_LABEL</type>
<position>-178,37</position>
<gparam>LABEL_TEXT i/p 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1949</ID>
<type>AA_LABEL</type>
<position>-178,30.5</position>
<gparam>LABEL_TEXT i/p 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1950</ID>
<type>AA_LABEL</type>
<position>-178,21.5</position>
<gparam>LABEL_TEXT i/p 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1951</ID>
<type>AA_LABEL</type>
<position>-178,16.5</position>
<gparam>LABEL_TEXT i/p 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1952</ID>
<type>AA_LABEL</type>
<position>-178,12.5</position>
<gparam>LABEL_TEXT i/p 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1961</ID>
<type>AA_TOGGLE</type>
<position>-244,-15.5</position>
<output>
<ID>OUT_0</ID>1430 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1963</ID>
<type>AA_TOGGLE</type>
<position>-233,-15</position>
<output>
<ID>OUT_0</ID>1431 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1964</ID>
<type>AA_TOGGLE</type>
<position>-223,-15</position>
<output>
<ID>OUT_0</ID>1432 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1965</ID>
<type>AA_TOGGLE</type>
<position>-215,-15</position>
<output>
<ID>OUT_0</ID>1433 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1972</ID>
<type>AA_TOGGLE</type>
<position>-283,-15</position>
<output>
<ID>OUT_0</ID>1427 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1973</ID>
<type>AA_TOGGLE</type>
<position>-272.5,-15</position>
<output>
<ID>OUT_0</ID>1434 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1974</ID>
<type>AA_TOGGLE</type>
<position>-262.5,-15</position>
<output>
<ID>OUT_0</ID>1428 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1975</ID>
<type>AA_TOGGLE</type>
<position>-255,-15</position>
<output>
<ID>OUT_0</ID>1429 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2003</ID>
<type>GA_LED</type>
<position>-281.5,61</position>
<input>
<ID>N_in3</ID>1403 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2004</ID>
<type>GA_LED</type>
<position>-271,61</position>
<input>
<ID>N_in3</ID>1404 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2005</ID>
<type>GA_LED</type>
<position>-261,61</position>
<input>
<ID>N_in3</ID>1405 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2006</ID>
<type>GA_LED</type>
<position>-253.5,61</position>
<input>
<ID>N_in3</ID>1406 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2007</ID>
<type>GA_LED</type>
<position>-242,61</position>
<input>
<ID>N_in3</ID>1407 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2022</ID>
<type>GA_LED</type>
<position>-223,61</position>
<input>
<ID>N_in3</ID>1409 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2024</ID>
<type>GA_LED</type>
<position>-233,61</position>
<input>
<ID>N_in3</ID>1408 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2026</ID>
<type>GA_LED</type>
<position>-215,61</position>
<input>
<ID>N_in3</ID>1410 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2028</ID>
<type>AA_TOGGLE</type>
<position>-303,29</position>
<output>
<ID>OUT_0</ID>1424 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2030</ID>
<type>AA_TOGGLE</type>
<position>-303,13</position>
<output>
<ID>OUT_0</ID>1426 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2032</ID>
<type>AA_TOGGLE</type>
<position>-303,20.5</position>
<output>
<ID>OUT_0</ID>1425 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2034</ID>
<type>AA_LABEL</type>
<position>-309.5,31.5</position>
<gparam>LABEL_TEXT Read</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2036</ID>
<type>AA_LABEL</type>
<position>-309,23.5</position>
<gparam>LABEL_TEXT Write</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2038</ID>
<type>AA_LABEL</type>
<position>-311,16</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2040</ID>
<type>AA_LABEL</type>
<position>-297,-14</position>
<gparam>LABEL_TEXT Data in</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2042</ID>
<type>AA_LABEL</type>
<position>-297.5,61.5</position>
<gparam>LABEL_TEXT Data out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2066</ID>
<type>DA_FROM</type>
<position>-281.5,68</position>
<input>
<ID>IN_0</ID>1403 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O1</lparam></gate>
<gate>
<ID>2068</ID>
<type>DA_FROM</type>
<position>-271,68</position>
<input>
<ID>IN_0</ID>1404 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O2</lparam></gate>
<gate>
<ID>2070</ID>
<type>DA_FROM</type>
<position>-261,68</position>
<input>
<ID>IN_0</ID>1405 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O3</lparam></gate>
<gate>
<ID>2072</ID>
<type>DA_FROM</type>
<position>-253.5,68</position>
<input>
<ID>IN_0</ID>1406 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O4</lparam></gate>
<gate>
<ID>2074</ID>
<type>DA_FROM</type>
<position>-242,68</position>
<input>
<ID>IN_0</ID>1407 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O5</lparam></gate>
<gate>
<ID>2076</ID>
<type>DA_FROM</type>
<position>-233,68</position>
<input>
<ID>IN_0</ID>1408 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O6</lparam></gate>
<gate>
<ID>2078</ID>
<type>DA_FROM</type>
<position>-223,68</position>
<input>
<ID>IN_0</ID>1409 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O7</lparam></gate>
<gate>
<ID>2080</ID>
<type>DA_FROM</type>
<position>-215,68</position>
<input>
<ID>IN_0</ID>1410 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O8</lparam></gate>
<gate>
<ID>2084</ID>
<type>DA_FROM</type>
<position>-8,-6450.5</position>
<input>
<ID>IN_0</ID>1423 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>2086</ID>
<type>DE_TO</type>
<position>-295.5,29</position>
<input>
<ID>IN_0</ID>1424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>2087</ID>
<type>DE_TO</type>
<position>-296,20.5</position>
<input>
<ID>IN_0</ID>1425 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>2088</ID>
<type>DE_TO</type>
<position>-296.5,13</position>
<input>
<ID>IN_0</ID>1426 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>2089</ID>
<type>DE_TO</type>
<position>-283,-8</position>
<input>
<ID>IN_0</ID>1427 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>2090</ID>
<type>DE_TO</type>
<position>-272.5,-8</position>
<input>
<ID>IN_0</ID>1434 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>2091</ID>
<type>DE_TO</type>
<position>-262.5,-8</position>
<input>
<ID>IN_0</ID>1428 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>2092</ID>
<type>DE_TO</type>
<position>-255,-8</position>
<input>
<ID>IN_0</ID>1429 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>2093</ID>
<type>DE_TO</type>
<position>-244,-8.5</position>
<input>
<ID>IN_0</ID>1430 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>2094</ID>
<type>DE_TO</type>
<position>-233,-8</position>
<input>
<ID>IN_0</ID>1431 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>2095</ID>
<type>DE_TO</type>
<position>-223,-8</position>
<input>
<ID>IN_0</ID>1432 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>2096</ID>
<type>DE_TO</type>
<position>-215,-8</position>
<input>
<ID>IN_0</ID>1433 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>2098</ID>
<type>BA_TRI_STATE</type>
<position>13,-6441</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1435 </input>
<output>
<ID>OUT_0</ID>1465 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2100</ID>
<type>DA_FROM</type>
<position>13,-6454</position>
<input>
<ID>IN_0</ID>1435 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>2101</ID>
<type>BA_TRI_STATE</type>
<position>75.5,-6441.5</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1436 </input>
<output>
<ID>OUT_0</ID>1466 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2102</ID>
<type>DA_FROM</type>
<position>75.5,-6455</position>
<input>
<ID>IN_0</ID>1436 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>2103</ID>
<type>BA_TRI_STATE</type>
<position>152,-6441.5</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1437 </input>
<output>
<ID>OUT_0</ID>1467 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2104</ID>
<type>DA_FROM</type>
<position>152,-6458</position>
<input>
<ID>IN_0</ID>1437 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>2105</ID>
<type>BA_TRI_STATE</type>
<position>234.5,-6441.5</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1438 </input>
<output>
<ID>OUT_0</ID>1468 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2106</ID>
<type>DA_FROM</type>
<position>234.5,-6457.5</position>
<input>
<ID>IN_0</ID>1438 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>2107</ID>
<type>BA_TRI_STATE</type>
<position>308,-6442</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1439 </input>
<output>
<ID>OUT_0</ID>1469 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2108</ID>
<type>DA_FROM</type>
<position>308,-6458</position>
<input>
<ID>IN_0</ID>1439 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>2109</ID>
<type>BA_TRI_STATE</type>
<position>396.5,-6442.5</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1440 </input>
<output>
<ID>OUT_0</ID>1470 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2110</ID>
<type>DA_FROM</type>
<position>397,-6458</position>
<input>
<ID>IN_0</ID>1440 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>2111</ID>
<type>BA_TRI_STATE</type>
<position>478,-6442.5</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1441 </input>
<output>
<ID>OUT_0</ID>1471 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2112</ID>
<type>DA_FROM</type>
<position>478,-6458.5</position>
<input>
<ID>IN_0</ID>1441 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>2113</ID>
<type>BA_TRI_STATE</type>
<position>562,-6442.5</position>
<input>
<ID>ENABLE_0</ID>1444 </input>
<input>
<ID>IN_0</ID>1442 </input>
<output>
<ID>OUT_0</ID>1472 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2114</ID>
<type>DA_FROM</type>
<position>562,-6458.5</position>
<input>
<ID>IN_0</ID>1442 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>2116</ID>
<type>DA_FROM</type>
<position>3.5,-6441</position>
<input>
<ID>IN_0</ID>1444 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>2118</ID>
<type>BA_TRI_STATE</type>
<position>63,426.5</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1457 </input>
<output>
<ID>OUT_0</ID>1445 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2119</ID>
<type>BA_TRI_STATE</type>
<position>143.5,426</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1458 </input>
<output>
<ID>OUT_0</ID>1447 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2127</ID>
<type>DE_TO</type>
<position>63,448.5</position>
<input>
<ID>IN_0</ID>1445 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O1</lparam></gate>
<gate>
<ID>2129</ID>
<type>DA_FROM</type>
<position>12,426.5</position>
<input>
<ID>IN_0</ID>1455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>2131</ID>
<type>DE_TO</type>
<position>143.5,447.5</position>
<input>
<ID>IN_0</ID>1447 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O2</lparam></gate>
<gate>
<ID>2132</ID>
<type>BA_TRI_STATE</type>
<position>220,428</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1459 </input>
<output>
<ID>OUT_0</ID>1448 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2133</ID>
<type>DE_TO</type>
<position>220,446.5</position>
<input>
<ID>IN_0</ID>1448 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O3</lparam></gate>
<gate>
<ID>2134</ID>
<type>BA_TRI_STATE</type>
<position>288,426.5</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1460 </input>
<output>
<ID>OUT_0</ID>1449 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2135</ID>
<type>DE_TO</type>
<position>288,448</position>
<input>
<ID>IN_0</ID>1449 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O4</lparam></gate>
<gate>
<ID>2136</ID>
<type>BA_TRI_STATE</type>
<position>379.5,428.5</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1461 </input>
<output>
<ID>OUT_0</ID>1450 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2137</ID>
<type>DE_TO</type>
<position>379.5,450</position>
<input>
<ID>IN_0</ID>1450 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O5</lparam></gate>
<gate>
<ID>2138</ID>
<type>BA_TRI_STATE</type>
<position>458.5,427.5</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1462 </input>
<output>
<ID>OUT_0</ID>1451 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2139</ID>
<type>DE_TO</type>
<position>458.5,449</position>
<input>
<ID>IN_0</ID>1451 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O6</lparam></gate>
<gate>
<ID>2140</ID>
<type>BA_TRI_STATE</type>
<position>543.5,424.5</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1463 </input>
<output>
<ID>OUT_0</ID>1452 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2141</ID>
<type>DE_TO</type>
<position>543.5,446</position>
<input>
<ID>IN_0</ID>1452 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O7</lparam></gate>
<gate>
<ID>2144</ID>
<type>BA_TRI_STATE</type>
<position>619.5,425</position>
<input>
<ID>ENABLE_0</ID>1455 </input>
<input>
<ID>IN_0</ID>1464 </input>
<output>
<ID>OUT_0</ID>1454 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2145</ID>
<type>DE_TO</type>
<position>619.5,446.5</position>
<input>
<ID>IN_0</ID>1454 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O8</lparam></gate>
<gate>
<ID>2147</ID>
<type>DA_FROM</type>
<position>-35,402</position>
<input>
<ID>IN_0</ID>1456 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-5066,40.5,-5066</points>
<connection>
<GID>58</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-5070.5,42.5,-5069</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-5070.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-5070.5,42.5,-5070.5</points>
<intersection>27.5 3</intersection>
<intersection>28.5 2</intersection>
<intersection>42.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>28.5,-5070.5,28.5,-5065</points>
<intersection>-5070.5 1</intersection>
<intersection>-5065 4</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-5070.5,27.5,-5057</points>
<connection>
<GID>1654</GID>
<name>OUT_0</name></connection>
<intersection>-5070.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28.5,-5065,29,-5065</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>28.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,41.5,-108,284.5</points>
<intersection>41.5 2</intersection>
<intersection>266.5 3</intersection>
<intersection>284.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,284.5,-6.5,284.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,41.5,-108,41.5</points>
<connection>
<GID>459</GID>
<name>OUT_6</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,266.5,-25,266.5</points>
<connection>
<GID>275</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-22.5,264.5,590,264.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>35 38</intersection>
<intersection>109 43</intersection>
<intersection>193 42</intersection>
<intersection>267 45</intersection>
<intersection>358 47</intersection>
<intersection>432 49</intersection>
<intersection>516 51</intersection>
<intersection>590 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>35,264.5,35,277</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>193,264.5,193,275</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>109,264.5,109,277</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>267,264.5,267,275</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>358,264.5,358,273.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>432,264.5,432,273.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>516,264.5,516,271.5</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>590,264.5,590,271.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>264.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,278,50.5,278</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<connection>
<GID>252</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,269.5,32,286.5</points>
<intersection>269.5 3</intersection>
<intersection>279 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,279,35,279</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,286.5,32,286.5</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,269.5,52.5,269.5</points>
<intersection>32 0</intersection>
<intersection>52.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52.5,269.5,52.5,275</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>269.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115,278,124,278</points>
<connection>
<GID>255</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>250</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,268,105.5,286.5</points>
<intersection>268 3</intersection>
<intersection>279 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,279,109,279</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,286.5,105.5,286.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105.5,268,126,268</points>
<intersection>105.5 0</intersection>
<intersection>126 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,268,126,275</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>268 3</intersection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,276,208.5,276</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<connection>
<GID>258</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,267.5,190,286.5</points>
<intersection>267.5 3</intersection>
<intersection>277 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,277,193,277</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,286.5,190,286.5</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>190,267.5,210.5,267.5</points>
<intersection>190 0</intersection>
<intersection>210.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210.5,267.5,210.5,273</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>267.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>273,276,282,276</points>
<connection>
<GID>261</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>256</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,266,263.5,286.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>266 3</intersection>
<intersection>277 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,277,267,277</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263.5,266,284,266</points>
<intersection>263.5 0</intersection>
<intersection>284 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>284,266,284,273</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>266 3</intersection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364,274.5,373.5,274.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<connection>
<GID>264</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,266,355,286.5</points>
<intersection>266 3</intersection>
<intersection>275.5 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,275.5,358,275.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,286.5,355,286.5</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>355,266,375.5,266</points>
<intersection>355 0</intersection>
<intersection>375.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375.5,266,375.5,271.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>266 3</intersection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>438,274.5,447,274.5</points>
<connection>
<GID>267</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>262</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,266,428.5,286.5</points>
<intersection>266 3</intersection>
<intersection>275.5 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,275.5,432,275.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,286.5,428.5,286.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428.5,266,449,266</points>
<intersection>428.5 0</intersection>
<intersection>449 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>449,266,449,271.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>266 3</intersection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,272.5,531.5,272.5</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<connection>
<GID>270</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,266.5,513,286.5</points>
<intersection>266.5 3</intersection>
<intersection>273.5 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513,273.5,516,273.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>512,286.5,513,286.5</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>513,266.5,533.5,266.5</points>
<intersection>513 0</intersection>
<intersection>533.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533.5,266.5,533.5,269.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>266.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>596,272.5,605,272.5</points>
<connection>
<GID>273</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>268</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,266.5,586.5,286.5</points>
<intersection>266.5 3</intersection>
<intersection>273.5 1</intersection>
<intersection>286.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586.5,273.5,590,273.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585.5,286.5,586.5,286.5</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586.5,266.5,607,266.5</points>
<intersection>586.5 0</intersection>
<intersection>607 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>607,266.5,607,269.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>266.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,283.5,579.5,283.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<connection>
<GID>272</GID>
<name>clock</name></connection>
<connection>
<GID>269</GID>
<name>clock</name></connection>
<connection>
<GID>266</GID>
<name>clock</name></connection>
<connection>
<GID>263</GID>
<name>clock</name></connection>
<connection>
<GID>260</GID>
<name>clock</name></connection>
<connection>
<GID>257</GID>
<name>clock</name></connection>
<connection>
<GID>254</GID>
<name>clock</name></connection>
<connection>
<GID>251</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,42.5,-109,374.5</points>
<intersection>42.5 2</intersection>
<intersection>356.5 3</intersection>
<intersection>374.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,374.5,-9.5,374.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,42.5,-109,42.5</points>
<connection>
<GID>459</GID>
<name>OUT_7</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,356.5,-28,356.5</points>
<connection>
<GID>301</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25.5,354.5,587,354.5</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>32 38</intersection>
<intersection>106 43</intersection>
<intersection>190 42</intersection>
<intersection>264 45</intersection>
<intersection>355 47</intersection>
<intersection>429 49</intersection>
<intersection>513 51</intersection>
<intersection>587 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32,354.5,32,367</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190,354.5,190,365</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106,354.5,106,367</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264,354.5,264,365</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355,354.5,355,363.5</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429,354.5,429,363.5</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513,354.5,513,361.5</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587,354.5,587,361.5</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>354.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,368,47.5,368</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>278</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,359.5,29,376.5</points>
<intersection>359.5 3</intersection>
<intersection>369 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,369,32,369</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,376.5,29,376.5</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,359.5,49.5,359.5</points>
<intersection>29 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,359.5,49.5,365</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>359.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112,368,121,368</points>
<connection>
<GID>281</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>276</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,358,102.5,376.5</points>
<intersection>358 3</intersection>
<intersection>369 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,369,106,369</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,376.5,102.5,376.5</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,358,123,358</points>
<intersection>102.5 0</intersection>
<intersection>123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123,358,123,365</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>358 3</intersection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,366,205.5,366</points>
<connection>
<GID>285</GID>
<name>OUT</name></connection>
<connection>
<GID>284</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,357.5,187,376.5</points>
<intersection>357.5 3</intersection>
<intersection>367 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,367,190,367</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,376.5,187,376.5</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,357.5,207.5,357.5</points>
<intersection>187 0</intersection>
<intersection>207.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207.5,357.5,207.5,363</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>357.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270,366,279,366</points>
<connection>
<GID>287</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>282</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,356,260.5,376.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>356 3</intersection>
<intersection>367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,367,264,367</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,356,281,356</points>
<intersection>260.5 0</intersection>
<intersection>281 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281,356,281,363</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>356 3</intersection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,364.5,370.5,364.5</points>
<connection>
<GID>291</GID>
<name>OUT</name></connection>
<connection>
<GID>290</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,356,352,376.5</points>
<intersection>356 3</intersection>
<intersection>365.5 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,365.5,355,365.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,376.5,352,376.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352,356,372.5,356</points>
<intersection>352 0</intersection>
<intersection>372.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372.5,356,372.5,361.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>356 3</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435,364.5,444,364.5</points>
<connection>
<GID>293</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>288</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,356,425.5,376.5</points>
<intersection>356 3</intersection>
<intersection>365.5 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,365.5,429,365.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,376.5,425.5,376.5</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,356,446,356</points>
<intersection>425.5 0</intersection>
<intersection>446 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446,356,446,361.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>356 3</intersection></vsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,362.5,528.5,362.5</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<connection>
<GID>296</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,356.5,510,376.5</points>
<intersection>356.5 3</intersection>
<intersection>363.5 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,363.5,513,363.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509,376.5,510,376.5</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510,356.5,530.5,356.5</points>
<intersection>510 0</intersection>
<intersection>530.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530.5,356.5,530.5,359.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>356.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593,362.5,602,362.5</points>
<connection>
<GID>299</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>294</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,356.5,583.5,376.5</points>
<intersection>356.5 3</intersection>
<intersection>363.5 1</intersection>
<intersection>376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,363.5,587,363.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,376.5,583.5,376.5</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583.5,356.5,604,356.5</points>
<intersection>583.5 0</intersection>
<intersection>604 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604,356.5,604,359.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>356.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,375,576.5,375</points>
<intersection>-3.5 2</intersection>
<intersection>22 10</intersection>
<intersection>95.5 9</intersection>
<intersection>180 8</intersection>
<intersection>254.5 7</intersection>
<intersection>345 6</intersection>
<intersection>418.5 5</intersection>
<intersection>503 4</intersection>
<intersection>576.5 3</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-3.5,373.5,-3.5,375</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>576.5,373.5,576.5,375</points>
<connection>
<GID>298</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>503,373.5,503,375</points>
<connection>
<GID>295</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>418.5,373.5,418.5,375</points>
<connection>
<GID>292</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>345,373.5,345,375</points>
<connection>
<GID>289</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>254.5,373.5,254.5,375</points>
<connection>
<GID>286</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>180,373.5,180,375</points>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>95.5,373.5,95.5,375</points>
<connection>
<GID>280</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>22,373.5,22,375</points>
<connection>
<GID>277</GID>
<name>clock</name></connection>
<intersection>375 1</intersection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,39.5,-84.5,116.5</points>
<intersection>39.5 2</intersection>
<intersection>98.5 3</intersection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84.5,116.5,-2.5,116.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,39.5,-84.5,39.5</points>
<connection>
<GID>459</GID>
<name>OUT_4</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-84.5,98.5,-21,98.5</points>
<connection>
<GID>327</GID>
<name>ENABLE_0</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-18.5,96.5,594,96.5</points>
<connection>
<GID>327</GID>
<name>OUT_0</name></connection>
<intersection>39 38</intersection>
<intersection>113 43</intersection>
<intersection>197 42</intersection>
<intersection>271 45</intersection>
<intersection>362 47</intersection>
<intersection>436 49</intersection>
<intersection>520 51</intersection>
<intersection>594 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>39,96.5,39,109</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>197,96.5,197,107</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>113,96.5,113,109</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>271,96.5,271,107</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>362,96.5,362,105.5</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>436,96.5,436,105.5</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>520,96.5,520,103.5</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>594,96.5,594,103.5</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>96.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,110,54.5,110</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<connection>
<GID>304</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,101.5,36,118.5</points>
<intersection>101.5 3</intersection>
<intersection>111 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,111,39,111</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,118.5,36,118.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,101.5,56.5,101.5</points>
<intersection>36 0</intersection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56.5,101.5,56.5,107</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>101.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,110,128,110</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>307</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,100,109.5,118.5</points>
<intersection>100 3</intersection>
<intersection>111 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,111,113,111</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,118.5,109.5,118.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>109.5,100,130,100</points>
<intersection>109.5 0</intersection>
<intersection>130 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130,100,130,107</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>100 3</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,108,212.5,108</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<connection>
<GID>310</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,99.5,194,118.5</points>
<intersection>99.5 3</intersection>
<intersection>109 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,109,197,109</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>193,118.5,194,118.5</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>194,99.5,214.5,99.5</points>
<intersection>194 0</intersection>
<intersection>214.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>214.5,99.5,214.5,105</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>99.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>277,108,286,108</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<connection>
<GID>313</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,98,267.5,118.5</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>98 3</intersection>
<intersection>109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,109,271,109</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>267.5,98,288,98</points>
<intersection>267.5 0</intersection>
<intersection>288 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>288,98,288,105</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>98 3</intersection></vsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,106,384,106</points>
<connection>
<GID>316</GID>
<name>ENABLE_0</name></connection>
<intersection>368 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>368,106,368,106.5</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<intersection>106 1</intersection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,98,359,118.5</points>
<intersection>98 3</intersection>
<intersection>107.5 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,107.5,362,107.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>358,118.5,359,118.5</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>359,98,386,98</points>
<intersection>359 0</intersection>
<intersection>386 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>386,98,386,103</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>98 3</intersection></vsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>442,106.5,451,106.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<connection>
<GID>319</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,98,432.5,118.5</points>
<intersection>98 3</intersection>
<intersection>107.5 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,107.5,436,107.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,118.5,432.5,118.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432.5,98,453,98</points>
<intersection>432.5 0</intersection>
<intersection>453 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>453,98,453,103.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>98 3</intersection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>526,104.5,535.5,104.5</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<connection>
<GID>322</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,98.5,517,118.5</points>
<intersection>98.5 3</intersection>
<intersection>105.5 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,105.5,520,105.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>516,118.5,517,118.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>517,98.5,537.5,98.5</points>
<intersection>517 0</intersection>
<intersection>537.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>537.5,98.5,537.5,101.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>98.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>600,104.5,609,104.5</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<connection>
<GID>325</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,98.5,590.5,118.5</points>
<intersection>98.5 3</intersection>
<intersection>105.5 1</intersection>
<intersection>118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,105.5,594,105.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,118.5,590.5,118.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>590.5,98.5,611,98.5</points>
<intersection>590.5 0</intersection>
<intersection>611 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>611,98.5,611,101.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>98.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,115.5,583.5,115.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<connection>
<GID>321</GID>
<name>clock</name></connection>
<connection>
<GID>318</GID>
<name>clock</name></connection>
<connection>
<GID>315</GID>
<name>clock</name></connection>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<connection>
<GID>303</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107,40.5,-107,206.5</points>
<intersection>40.5 2</intersection>
<intersection>188.5 3</intersection>
<intersection>206.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-107,206.5,-5.5,206.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,40.5,-107,40.5</points>
<connection>
<GID>459</GID>
<name>OUT_5</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-107,188.5,-24,188.5</points>
<connection>
<GID>353</GID>
<name>ENABLE_0</name></connection>
<intersection>-107 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21.5,186.5,591,186.5</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>36 38</intersection>
<intersection>110 43</intersection>
<intersection>194 42</intersection>
<intersection>268 45</intersection>
<intersection>359 47</intersection>
<intersection>433 49</intersection>
<intersection>517 51</intersection>
<intersection>591 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36,186.5,36,199</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194,186.5,194,197</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110,186.5,110,199</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268,186.5,268,197</points>
<connection>
<GID>334</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359,186.5,359,195.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433,186.5,433,195.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517,186.5,517,193.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591,186.5,591,193.5</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>186.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,200,51.5,200</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<connection>
<GID>330</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,191.5,33,208.5</points>
<intersection>191.5 3</intersection>
<intersection>201 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,201,36,201</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,208.5,33,208.5</points>
<connection>
<GID>329</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,191.5,53.5,191.5</points>
<intersection>33 0</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,191.5,53.5,197</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>191.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116,200,125,200</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<connection>
<GID>333</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,190,106.5,208.5</points>
<intersection>190 3</intersection>
<intersection>201 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,201,110,201</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,208.5,106.5,208.5</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,190,127,190</points>
<intersection>106.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,190,127,197</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>190 3</intersection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,198,209.5,198</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<connection>
<GID>336</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,189.5,191,208.5</points>
<intersection>189.5 3</intersection>
<intersection>199 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,199,194,199</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,208.5,191,208.5</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191,189.5,211.5,189.5</points>
<intersection>191 0</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211.5,189.5,211.5,195</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>189.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274,198,283,198</points>
<connection>
<GID>334</GID>
<name>OUT</name></connection>
<connection>
<GID>339</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,188,264.5,208.5</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>188 3</intersection>
<intersection>199 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,199,268,199</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264.5,188,285,188</points>
<intersection>264.5 0</intersection>
<intersection>285 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285,188,285,195</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>188 3</intersection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365,196.5,374.5,196.5</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<connection>
<GID>342</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,188,356,208.5</points>
<intersection>188 3</intersection>
<intersection>197.5 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,197.5,359,197.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355,208.5,356,208.5</points>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356,188,376.5,188</points>
<intersection>356 0</intersection>
<intersection>376.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376.5,188,376.5,193.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>188 3</intersection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439,196.5,448,196.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<connection>
<GID>345</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,188,429.5,208.5</points>
<intersection>188 3</intersection>
<intersection>197.5 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,197.5,433,197.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,208.5,429.5,208.5</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,188,450,188</points>
<intersection>429.5 0</intersection>
<intersection>450 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450,188,450,193.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>188 3</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523,194.5,532.5,194.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<connection>
<GID>348</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,188.5,514,208.5</points>
<intersection>188.5 3</intersection>
<intersection>195.5 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,195.5,517,195.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,208.5,514,208.5</points>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514,188.5,534.5,188.5</points>
<intersection>514 0</intersection>
<intersection>534.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534.5,188.5,534.5,191.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>188.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597,194.5,606,194.5</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<connection>
<GID>351</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,188.5,587.5,208.5</points>
<intersection>188.5 3</intersection>
<intersection>195.5 1</intersection>
<intersection>208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,195.5,591,195.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586.5,208.5,587.5,208.5</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587.5,188.5,608,188.5</points>
<intersection>587.5 0</intersection>
<intersection>608 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608,188.5,608,191.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>188.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,205.5,580.5,205.5</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<connection>
<GID>350</GID>
<name>clock</name></connection>
<connection>
<GID>347</GID>
<name>clock</name></connection>
<connection>
<GID>344</GID>
<name>clock</name></connection>
<connection>
<GID>341</GID>
<name>clock</name></connection>
<connection>
<GID>338</GID>
<name>clock</name></connection>
<connection>
<GID>335</GID>
<name>clock</name></connection>
<connection>
<GID>332</GID>
<name>clock</name></connection>
<connection>
<GID>329</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107,-109.5,-107,37.5</points>
<intersection>-109.5 3</intersection>
<intersection>-91.5 1</intersection>
<intersection>37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-107,-91.5,-4.5,-91.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,37.5,-107,37.5</points>
<connection>
<GID>459</GID>
<name>OUT_2</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-107,-109.5,-23,-109.5</points>
<connection>
<GID>379</GID>
<name>ENABLE_0</name></connection>
<intersection>-107 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-20.5,-111.5,592,-111.5</points>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection>
<intersection>37 38</intersection>
<intersection>111 43</intersection>
<intersection>195 42</intersection>
<intersection>269 45</intersection>
<intersection>360 47</intersection>
<intersection>434 49</intersection>
<intersection>518 51</intersection>
<intersection>592 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>37,-111.5,37,-99</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>195,-111.5,195,-101</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>111,-111.5,111,-99</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>269,-111.5,269,-101</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>360,-111.5,360,-102.5</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>434,-111.5,434,-102.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>518,-111.5,518,-104.5</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>592,-111.5,592,-104.5</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>-111.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-98,52.5,-98</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<connection>
<GID>356</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-106.5,34,-89.5</points>
<intersection>-106.5 3</intersection>
<intersection>-97 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-97,37,-97</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-89.5,34,-89.5</points>
<connection>
<GID>355</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-106.5,54.5,-106.5</points>
<intersection>34 0</intersection>
<intersection>54.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54.5,-106.5,54.5,-101</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>117,-98,126,-98</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<connection>
<GID>359</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-108,107.5,-89.5</points>
<intersection>-108 3</intersection>
<intersection>-97 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-97,111,-97</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-89.5,107.5,-89.5</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-108,128,-108</points>
<intersection>107.5 0</intersection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-108,128,-101</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>-108 3</intersection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201,-100,210.5,-100</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<connection>
<GID>362</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-108.5,192,-89.5</points>
<intersection>-108.5 3</intersection>
<intersection>-99 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-99,195,-99</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-89.5,192,-89.5</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>192,-108.5,212.5,-108.5</points>
<intersection>192 0</intersection>
<intersection>212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>212.5,-108.5,212.5,-103</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-108.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>275,-100,284,-100</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<connection>
<GID>365</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-110,265.5,-89.5</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<intersection>-110 3</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,-99,269,-99</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>265.5,-110,286,-110</points>
<intersection>265.5 0</intersection>
<intersection>286 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>286,-110,286,-103</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-110 3</intersection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366,-101.5,375.5,-101.5</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<connection>
<GID>368</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-110,357,-89.5</points>
<intersection>-110 3</intersection>
<intersection>-100.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-100.5,360,-100.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356,-89.5,357,-89.5</points>
<connection>
<GID>367</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-110,377.5,-110</points>
<intersection>357 0</intersection>
<intersection>377.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>377.5,-110,377.5,-104.5</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>-110 3</intersection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>440,-101.5,449,-101.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<connection>
<GID>371</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,-110,430.5,-89.5</points>
<intersection>-110 3</intersection>
<intersection>-100.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430.5,-100.5,434,-100.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>429.5,-89.5,430.5,-89.5</points>
<connection>
<GID>370</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>430.5,-110,451,-110</points>
<intersection>430.5 0</intersection>
<intersection>451 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>451,-110,451,-104.5</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-110 3</intersection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524,-103.5,533.5,-103.5</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<connection>
<GID>374</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-109.5,515,-89.5</points>
<intersection>-109.5 3</intersection>
<intersection>-102.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515,-102.5,518,-102.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,-89.5,515,-89.5</points>
<connection>
<GID>373</GID>
<name>OUT_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>515,-109.5,535.5,-109.5</points>
<intersection>515 0</intersection>
<intersection>535.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535.5,-109.5,535.5,-106.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-109.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>598,-103.5,607,-103.5</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<connection>
<GID>377</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588.5,-109.5,588.5,-89.5</points>
<intersection>-109.5 3</intersection>
<intersection>-102.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588.5,-102.5,592,-102.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-89.5,588.5,-89.5</points>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>588.5,-109.5,609,-109.5</points>
<intersection>588.5 0</intersection>
<intersection>609 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>609,-109.5,609,-106.5</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-109.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-92.5,581.5,-92.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<connection>
<GID>376</GID>
<name>clock</name></connection>
<connection>
<GID>373</GID>
<name>clock</name></connection>
<connection>
<GID>370</GID>
<name>clock</name></connection>
<connection>
<GID>367</GID>
<name>clock</name></connection>
<connection>
<GID>364</GID>
<name>clock</name></connection>
<connection>
<GID>361</GID>
<name>clock</name></connection>
<connection>
<GID>355</GID>
<name>clock</name></connection>
<connection>
<GID>358</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-19.5,-106,38.5</points>
<intersection>-19.5 3</intersection>
<intersection>-1.5 1</intersection>
<intersection>38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106,-1.5,-7.5,-1.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,38.5,-106,38.5</points>
<connection>
<GID>459</GID>
<name>OUT_3</name></connection>
<intersection>-106 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-106,-19.5,-26,-19.5</points>
<connection>
<GID>405</GID>
<name>ENABLE_0</name></connection>
<intersection>-106 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-21.5,589,-21.5</points>
<connection>
<GID>405</GID>
<name>OUT_0</name></connection>
<intersection>34 38</intersection>
<intersection>108 43</intersection>
<intersection>192 42</intersection>
<intersection>266 45</intersection>
<intersection>357 47</intersection>
<intersection>431 49</intersection>
<intersection>515 51</intersection>
<intersection>589 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34,-21.5,34,-9</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192,-21.5,192,-11</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108,-21.5,108,-9</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266,-21.5,266,-11</points>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357,-21.5,357,-12.5</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431,-21.5,431,-12.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515,-21.5,515,-14.5</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589,-21.5,589,-14.5</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<intersection>-21.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-8,49.5,-8</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<connection>
<GID>382</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-16.5,31,0.5</points>
<intersection>-16.5 3</intersection>
<intersection>-7 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-7,34,-7</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,0.5,31,0.5</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-16.5,51.5,-16.5</points>
<intersection>31 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-16.5,51.5,-11</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-16.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114,-8,123,-8</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<connection>
<GID>385</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-18,104.5,0.5</points>
<intersection>-18 3</intersection>
<intersection>-7 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-7,108,-7</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,0.5,104.5,0.5</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-18,125,-18</points>
<intersection>104.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-18,125,-11</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>-18 3</intersection></vsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-10,207.5,-10</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<connection>
<GID>388</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-18.5,189,0.5</points>
<intersection>-18.5 3</intersection>
<intersection>-9 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-9,192,-9</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188,0.5,189,0.5</points>
<connection>
<GID>387</GID>
<name>OUT_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189,-18.5,209.5,-18.5</points>
<intersection>189 0</intersection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,-18.5,209.5,-13</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-18.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272,-10,281,-10</points>
<connection>
<GID>386</GID>
<name>OUT</name></connection>
<connection>
<GID>391</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-20,262.5,0.5</points>
<connection>
<GID>390</GID>
<name>OUT_0</name></connection>
<intersection>-20 3</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-9,266,-9</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262.5,-20,283,-20</points>
<intersection>262.5 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-20,283,-13</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-20 3</intersection></vsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363,-11.5,372.5,-11.5</points>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<connection>
<GID>394</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-20,354,0.5</points>
<intersection>-20 3</intersection>
<intersection>-10.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-10.5,357,-10.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,0.5,354,0.5</points>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354,-20,374.5,-20</points>
<intersection>354 0</intersection>
<intersection>374.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374.5,-20,374.5,-14.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-20 3</intersection></vsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437,-11.5,446,-11.5</points>
<connection>
<GID>392</GID>
<name>OUT</name></connection>
<connection>
<GID>397</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-20,427.5,0.5</points>
<intersection>-20 3</intersection>
<intersection>-10.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-10.5,431,-10.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426.5,0.5,427.5,0.5</points>
<connection>
<GID>396</GID>
<name>OUT_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-20,448,-20</points>
<intersection>427.5 0</intersection>
<intersection>448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448,-20,448,-14.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-20 3</intersection></vsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521,-13.5,530.5,-13.5</points>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<connection>
<GID>400</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,-19.5,512,0.5</points>
<intersection>-19.5 3</intersection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-12.5,515,-12.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,0.5,512,0.5</points>
<connection>
<GID>399</GID>
<name>OUT_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512,-19.5,532.5,-19.5</points>
<intersection>512 0</intersection>
<intersection>532.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532.5,-19.5,532.5,-16.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>-19.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595,-13.5,604,-13.5</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<connection>
<GID>403</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-19.5,585.5,0.5</points>
<intersection>-19.5 3</intersection>
<intersection>-12.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-12.5,589,-12.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,0.5,585.5,0.5</points>
<connection>
<GID>402</GID>
<name>OUT_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-19.5,606,-19.5</points>
<intersection>585.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-19.5,606,-16.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>-19.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-2.5,578.5,-2.5</points>
<connection>
<GID>387</GID>
<name>clock</name></connection>
<connection>
<GID>384</GID>
<name>clock</name></connection>
<connection>
<GID>381</GID>
<name>clock</name></connection>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<connection>
<GID>402</GID>
<name>clock</name></connection>
<connection>
<GID>399</GID>
<name>clock</name></connection>
<connection>
<GID>396</GID>
<name>clock</name></connection>
<connection>
<GID>393</GID>
<name>clock</name></connection>
<connection>
<GID>390</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-277.5,-110,35.5</points>
<intersection>-277.5 3</intersection>
<intersection>-259.5 1</intersection>
<intersection>35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-259.5,-0.5,-259.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,35.5,-110,35.5</points>
<connection>
<GID>459</GID>
<name>OUT_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-277.5,-19,-277.5</points>
<connection>
<GID>431</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-16.5,-279.5,596,-279.5</points>
<connection>
<GID>431</GID>
<name>OUT_0</name></connection>
<intersection>41 38</intersection>
<intersection>115 43</intersection>
<intersection>199 42</intersection>
<intersection>273 45</intersection>
<intersection>364 47</intersection>
<intersection>438 49</intersection>
<intersection>522 51</intersection>
<intersection>596 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>41,-279.5,41,-267</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>199,-279.5,199,-269</points>
<connection>
<GID>415</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>115,-279.5,115,-267</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>273,-279.5,273,-269</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>364,-279.5,364,-270.5</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>438,-279.5,438,-270.5</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>522,-279.5,522,-272.5</points>
<connection>
<GID>427</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>596,-279.5,596,-272.5</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>-279.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-266,56.5,-266</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<connection>
<GID>408</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-274.5,38,-257.5</points>
<intersection>-274.5 3</intersection>
<intersection>-265 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-265,41,-265</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-257.5,38,-257.5</points>
<connection>
<GID>407</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-274.5,58.5,-274.5</points>
<intersection>38 0</intersection>
<intersection>58.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>58.5,-274.5,58.5,-269</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>-274.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>121,-266,130,-266</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<connection>
<GID>411</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-276,111.5,-257.5</points>
<intersection>-276 3</intersection>
<intersection>-265 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-265,115,-265</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-257.5,111.5,-257.5</points>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>111.5,-276,132,-276</points>
<intersection>111.5 0</intersection>
<intersection>132 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132,-276,132,-269</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>-276 3</intersection></vsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-268,214.5,-268</points>
<connection>
<GID>415</GID>
<name>OUT</name></connection>
<connection>
<GID>414</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-276.5,196,-257.5</points>
<intersection>-276.5 3</intersection>
<intersection>-267 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196,-267,199,-267</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,-257.5,196,-257.5</points>
<connection>
<GID>413</GID>
<name>OUT_0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>196,-276.5,216.5,-276.5</points>
<intersection>196 0</intersection>
<intersection>216.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>216.5,-276.5,216.5,-271</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>-276.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>279,-268,288,-268</points>
<connection>
<GID>412</GID>
<name>OUT</name></connection>
<connection>
<GID>417</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-278,269.5,-257.5</points>
<connection>
<GID>416</GID>
<name>OUT_0</name></connection>
<intersection>-278 3</intersection>
<intersection>-267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,-267,273,-267</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>269.5,-278,290,-278</points>
<intersection>269.5 0</intersection>
<intersection>290 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>290,-278,290,-271</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>-278 3</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>370,-269.5,379.5,-269.5</points>
<connection>
<GID>421</GID>
<name>OUT</name></connection>
<connection>
<GID>420</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-278,361,-257.5</points>
<intersection>-278 3</intersection>
<intersection>-268.5 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-268.5,364,-268.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>360,-257.5,361,-257.5</points>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>361,-278,381.5,-278</points>
<intersection>361 0</intersection>
<intersection>381.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>381.5,-278,381.5,-272.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>-278 3</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>444,-269.5,453,-269.5</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<connection>
<GID>423</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-278,434.5,-257.5</points>
<intersection>-278 3</intersection>
<intersection>-268.5 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-268.5,438,-268.5</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-257.5,434.5,-257.5</points>
<connection>
<GID>422</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>434.5,-278,455,-278</points>
<intersection>434.5 0</intersection>
<intersection>455 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>455,-278,455,-272.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>-278 3</intersection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>528,-271.5,537.5,-271.5</points>
<connection>
<GID>427</GID>
<name>OUT</name></connection>
<connection>
<GID>426</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519,-277.5,519,-257.5</points>
<intersection>-277.5 3</intersection>
<intersection>-270.5 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>519,-270.5,522,-270.5</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>519 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>518,-257.5,519,-257.5</points>
<connection>
<GID>425</GID>
<name>OUT_0</name></connection>
<intersection>519 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>519,-277.5,539.5,-277.5</points>
<intersection>519 0</intersection>
<intersection>539.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>539.5,-277.5,539.5,-274.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>-277.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>602,-271.5,611,-271.5</points>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<connection>
<GID>429</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-277.5,592.5,-257.5</points>
<intersection>-277.5 3</intersection>
<intersection>-270.5 1</intersection>
<intersection>-257.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-270.5,596,-270.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>591.5,-257.5,592.5,-257.5</points>
<connection>
<GID>428</GID>
<name>OUT_0</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>592.5,-277.5,613,-277.5</points>
<intersection>592.5 0</intersection>
<intersection>613 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>613,-277.5,613,-274.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>-277.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-260.5,585.5,-260.5</points>
<connection>
<GID>430</GID>
<name>OUT</name></connection>
<connection>
<GID>428</GID>
<name>clock</name></connection>
<connection>
<GID>425</GID>
<name>clock</name></connection>
<connection>
<GID>422</GID>
<name>clock</name></connection>
<connection>
<GID>419</GID>
<name>clock</name></connection>
<connection>
<GID>416</GID>
<name>clock</name></connection>
<connection>
<GID>413</GID>
<name>clock</name></connection>
<connection>
<GID>410</GID>
<name>clock</name></connection>
<connection>
<GID>407</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-187.5,-108,36.5</points>
<intersection>-187.5 3</intersection>
<intersection>-169.5 1</intersection>
<intersection>36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-169.5,-3.5,-169.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,36.5,-108,36.5</points>
<connection>
<GID>459</GID>
<name>OUT_1</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-187.5,-22,-187.5</points>
<connection>
<GID>457</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-19.5,-189.5,593,-189.5</points>
<connection>
<GID>457</GID>
<name>OUT_0</name></connection>
<intersection>38 38</intersection>
<intersection>112 43</intersection>
<intersection>196 42</intersection>
<intersection>270 45</intersection>
<intersection>361 47</intersection>
<intersection>435 49</intersection>
<intersection>519 51</intersection>
<intersection>593 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>38,-189.5,38,-177</points>
<connection>
<GID>435</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>196,-189.5,196,-179</points>
<connection>
<GID>441</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>112,-189.5,112,-177</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>270,-189.5,270,-179</points>
<connection>
<GID>438</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>361,-189.5,361,-180.5</points>
<connection>
<GID>447</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>435,-189.5,435,-180.5</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>519,-189.5,519,-182.5</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>593,-189.5,593,-182.5</points>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>-189.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-176,53.5,-176</points>
<connection>
<GID>435</GID>
<name>OUT</name></connection>
<connection>
<GID>434</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-184.5,35,-167.5</points>
<intersection>-184.5 3</intersection>
<intersection>-175 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-175,38,-175</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-167.5,35,-167.5</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-184.5,55.5,-184.5</points>
<intersection>35 0</intersection>
<intersection>55.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55.5,-184.5,55.5,-179</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>-184.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>118,-176,127,-176</points>
<connection>
<GID>432</GID>
<name>OUT</name></connection>
<connection>
<GID>437</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-186,108.5,-167.5</points>
<intersection>-186 3</intersection>
<intersection>-175 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-175,112,-175</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-167.5,108.5,-167.5</points>
<connection>
<GID>436</GID>
<name>OUT_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108.5,-186,129,-186</points>
<intersection>108.5 0</intersection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-186,129,-179</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>-186 3</intersection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-178,211.5,-178</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<connection>
<GID>440</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-186.5,193,-167.5</points>
<intersection>-186.5 3</intersection>
<intersection>-177 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-177,196,-177</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>192,-167.5,193,-167.5</points>
<connection>
<GID>439</GID>
<name>OUT_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>193,-186.5,213.5,-186.5</points>
<intersection>193 0</intersection>
<intersection>213.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>213.5,-186.5,213.5,-181</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>-186.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>276,-178,285,-178</points>
<connection>
<GID>438</GID>
<name>OUT</name></connection>
<connection>
<GID>443</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-188,266.5,-167.5</points>
<connection>
<GID>442</GID>
<name>OUT_0</name></connection>
<intersection>-188 3</intersection>
<intersection>-177 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-177,270,-177</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-188,287,-188</points>
<intersection>266.5 0</intersection>
<intersection>287 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>287,-188,287,-181</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-188 3</intersection></vsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367,-179.5,376.5,-179.5</points>
<connection>
<GID>447</GID>
<name>OUT</name></connection>
<connection>
<GID>446</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358,-188,358,-167.5</points>
<intersection>-188 3</intersection>
<intersection>-178.5 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358,-178.5,361,-178.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-167.5,358,-167.5</points>
<connection>
<GID>445</GID>
<name>OUT_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>358,-188,378.5,-188</points>
<intersection>358 0</intersection>
<intersection>378.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>378.5,-188,378.5,-182.5</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>-188 3</intersection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>441,-179.5,450,-179.5</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<connection>
<GID>449</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,-188,431.5,-167.5</points>
<intersection>-188 3</intersection>
<intersection>-178.5 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,-178.5,435,-178.5</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>430.5,-167.5,431.5,-167.5</points>
<connection>
<GID>448</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>431.5,-188,452,-188</points>
<intersection>431.5 0</intersection>
<intersection>452 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>452,-188,452,-182.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>-188 3</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,-187.5,516,-167.5</points>
<intersection>-187.5 3</intersection>
<intersection>-180.5 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,-180.5,519,-180.5</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515,-167.5,516,-167.5</points>
<connection>
<GID>451</GID>
<name>OUT_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>516,-187.5,536.5,-187.5</points>
<intersection>516 0</intersection>
<intersection>536.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>536.5,-187.5,536.5,-184.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>-187.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>599,-181.5,608,-181.5</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<connection>
<GID>455</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-187.5,589.5,-167.5</points>
<intersection>-187.5 3</intersection>
<intersection>-180.5 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589.5,-180.5,593,-180.5</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-167.5,589.5,-167.5</points>
<connection>
<GID>454</GID>
<name>OUT_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>589.5,-187.5,610,-187.5</points>
<intersection>589.5 0</intersection>
<intersection>610 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>610,-187.5,610,-184.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>-187.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-170.5,582.5,-170.5</points>
<connection>
<GID>456</GID>
<name>OUT</name></connection>
<connection>
<GID>454</GID>
<name>clock</name></connection>
<connection>
<GID>451</GID>
<name>clock</name></connection>
<connection>
<GID>448</GID>
<name>clock</name></connection>
<connection>
<GID>445</GID>
<name>clock</name></connection>
<connection>
<GID>442</GID>
<name>clock</name></connection>
<connection>
<GID>439</GID>
<name>clock</name></connection>
<connection>
<GID>436</GID>
<name>clock</name></connection>
<connection>
<GID>433</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-784,-108,-541</points>
<intersection>-784 2</intersection>
<intersection>-559 3</intersection>
<intersection>-541 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-541,-6.5,-541</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-784,-108,-784</points>
<connection>
<GID>529</GID>
<name>OUT_6</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-559,-25,-559</points>
<connection>
<GID>555</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-22.5,-561,590,-561</points>
<connection>
<GID>555</GID>
<name>OUT_0</name></connection>
<intersection>35 38</intersection>
<intersection>109 43</intersection>
<intersection>193 42</intersection>
<intersection>267 45</intersection>
<intersection>358 47</intersection>
<intersection>432 49</intersection>
<intersection>516 51</intersection>
<intersection>590 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>35,-561,35,-548.5</points>
<connection>
<GID>533</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>193,-561,193,-550.5</points>
<connection>
<GID>539</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>109,-561,109,-548.5</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>267,-561,267,-550.5</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>358,-561,358,-552</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>432,-561,432,-552</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>516,-561,516,-554</points>
<connection>
<GID>551</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>590,-561,590,-554</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<intersection>-561 33</intersection></vsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-547.5,50.5,-547.5</points>
<connection>
<GID>533</GID>
<name>OUT</name></connection>
<connection>
<GID>532</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-556,32,-539</points>
<intersection>-556 3</intersection>
<intersection>-546.5 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-546.5,35,-546.5</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-539,32,-539</points>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-556,52.5,-556</points>
<intersection>32 0</intersection>
<intersection>52.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52.5,-556,52.5,-550.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>-556 3</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115,-547.5,124,-547.5</points>
<connection>
<GID>530</GID>
<name>OUT</name></connection>
<connection>
<GID>535</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-557.5,105.5,-539</points>
<intersection>-557.5 3</intersection>
<intersection>-546.5 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-546.5,109,-546.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-539,105.5,-539</points>
<connection>
<GID>534</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105.5,-557.5,126,-557.5</points>
<intersection>105.5 0</intersection>
<intersection>126 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,-557.5,126,-550.5</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>-557.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-549.5,208.5,-549.5</points>
<connection>
<GID>539</GID>
<name>OUT</name></connection>
<connection>
<GID>538</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-558,190,-539</points>
<intersection>-558 3</intersection>
<intersection>-548.5 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-548.5,193,-548.5</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,-539,190,-539</points>
<connection>
<GID>537</GID>
<name>OUT_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>190,-558,210.5,-558</points>
<intersection>190 0</intersection>
<intersection>210.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210.5,-558,210.5,-552.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>-558 3</intersection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>273,-549.5,282,-549.5</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<connection>
<GID>541</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,-559.5,263.5,-539</points>
<connection>
<GID>540</GID>
<name>OUT_0</name></connection>
<intersection>-559.5 3</intersection>
<intersection>-548.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,-548.5,267,-548.5</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263.5,-559.5,284,-559.5</points>
<intersection>263.5 0</intersection>
<intersection>284 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>284,-559.5,284,-552.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>-559.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364,-551,373.5,-551</points>
<connection>
<GID>545</GID>
<name>OUT</name></connection>
<connection>
<GID>544</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-559.5,355,-539</points>
<intersection>-559.5 3</intersection>
<intersection>-550 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-550,358,-550</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-539,355,-539</points>
<connection>
<GID>543</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>355,-559.5,375.5,-559.5</points>
<intersection>355 0</intersection>
<intersection>375.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375.5,-559.5,375.5,-554</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>-559.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>438,-551,447,-551</points>
<connection>
<GID>542</GID>
<name>OUT</name></connection>
<connection>
<GID>547</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,-559.5,428.5,-539</points>
<intersection>-559.5 3</intersection>
<intersection>-550 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,-550,432,-550</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,-539,428.5,-539</points>
<connection>
<GID>546</GID>
<name>OUT_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428.5,-559.5,449,-559.5</points>
<intersection>428.5 0</intersection>
<intersection>449 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>449,-559.5,449,-554</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>-559.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,-553,531.5,-553</points>
<connection>
<GID>551</GID>
<name>OUT</name></connection>
<connection>
<GID>550</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,-559,513,-539</points>
<intersection>-559 3</intersection>
<intersection>-552 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513,-552,516,-552</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>512,-539,513,-539</points>
<connection>
<GID>549</GID>
<name>OUT_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>513,-559,533.5,-559</points>
<intersection>513 0</intersection>
<intersection>533.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533.5,-559,533.5,-556</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<intersection>-559 3</intersection></vsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>596,-553,605,-553</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<connection>
<GID>553</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,-559,586.5,-539</points>
<intersection>-559 3</intersection>
<intersection>-552 1</intersection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586.5,-552,590,-552</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585.5,-539,586.5,-539</points>
<connection>
<GID>552</GID>
<name>OUT_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586.5,-559,607,-559</points>
<intersection>586.5 0</intersection>
<intersection>607 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>607,-559,607,-556</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>-559 3</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-542,579.5,-542</points>
<connection>
<GID>554</GID>
<name>OUT</name></connection>
<connection>
<GID>552</GID>
<name>clock</name></connection>
<connection>
<GID>549</GID>
<name>clock</name></connection>
<connection>
<GID>546</GID>
<name>clock</name></connection>
<connection>
<GID>543</GID>
<name>clock</name></connection>
<connection>
<GID>540</GID>
<name>clock</name></connection>
<connection>
<GID>537</GID>
<name>clock</name></connection>
<connection>
<GID>534</GID>
<name>clock</name></connection>
<connection>
<GID>531</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-783,-109,-451</points>
<intersection>-783 2</intersection>
<intersection>-469 3</intersection>
<intersection>-451 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-451,-9.5,-451</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-783,-109,-783</points>
<connection>
<GID>529</GID>
<name>OUT_7</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-469,-28,-469</points>
<connection>
<GID>581</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25.5,-471,587,-471</points>
<connection>
<GID>581</GID>
<name>OUT_0</name></connection>
<intersection>32 38</intersection>
<intersection>106 43</intersection>
<intersection>190 42</intersection>
<intersection>264 45</intersection>
<intersection>355 47</intersection>
<intersection>429 49</intersection>
<intersection>513 51</intersection>
<intersection>587 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32,-471,32,-458.5</points>
<connection>
<GID>559</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190,-471,190,-460.5</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106,-471,106,-458.5</points>
<connection>
<GID>556</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264,-471,264,-460.5</points>
<connection>
<GID>562</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355,-471,355,-462</points>
<connection>
<GID>571</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429,-471,429,-462</points>
<connection>
<GID>568</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513,-471,513,-464</points>
<connection>
<GID>577</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587,-471,587,-464</points>
<connection>
<GID>574</GID>
<name>IN_1</name></connection>
<intersection>-471 33</intersection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-457.5,47.5,-457.5</points>
<connection>
<GID>559</GID>
<name>OUT</name></connection>
<connection>
<GID>558</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-466,29,-449</points>
<intersection>-466 3</intersection>
<intersection>-456.5 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-456.5,32,-456.5</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-449,29,-449</points>
<connection>
<GID>557</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-466,49.5,-466</points>
<intersection>29 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-466,49.5,-460.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>-466 3</intersection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112,-457.5,121,-457.5</points>
<connection>
<GID>556</GID>
<name>OUT</name></connection>
<connection>
<GID>561</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-467.5,102.5,-449</points>
<intersection>-467.5 3</intersection>
<intersection>-456.5 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-456.5,106,-456.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-449,102.5,-449</points>
<connection>
<GID>560</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-467.5,123,-467.5</points>
<intersection>102.5 0</intersection>
<intersection>123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123,-467.5,123,-460.5</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>-467.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,-459.5,205.5,-459.5</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<connection>
<GID>564</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-468,187,-449</points>
<intersection>-468 3</intersection>
<intersection>-458.5 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-458.5,190,-458.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-449,187,-449</points>
<connection>
<GID>563</GID>
<name>OUT_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,-468,207.5,-468</points>
<intersection>187 0</intersection>
<intersection>207.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207.5,-468,207.5,-462.5</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>-468 3</intersection></vsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270,-459.5,279,-459.5</points>
<connection>
<GID>562</GID>
<name>OUT</name></connection>
<connection>
<GID>567</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-469.5,260.5,-449</points>
<connection>
<GID>566</GID>
<name>OUT_0</name></connection>
<intersection>-469.5 3</intersection>
<intersection>-458.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-458.5,264,-458.5</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-469.5,281,-469.5</points>
<intersection>260.5 0</intersection>
<intersection>281 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281,-469.5,281,-462.5</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>-469.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-461,370.5,-461</points>
<connection>
<GID>571</GID>
<name>OUT</name></connection>
<connection>
<GID>570</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-469.5,352,-449</points>
<intersection>-469.5 3</intersection>
<intersection>-460 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-460,355,-460</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-449,352,-449</points>
<connection>
<GID>569</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352,-469.5,372.5,-469.5</points>
<intersection>352 0</intersection>
<intersection>372.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372.5,-469.5,372.5,-464</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>-469.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435,-461,444,-461</points>
<connection>
<GID>568</GID>
<name>OUT</name></connection>
<connection>
<GID>573</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-469.5,425.5,-449</points>
<intersection>-469.5 3</intersection>
<intersection>-460 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,-460,429,-460</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,-449,425.5,-449</points>
<connection>
<GID>572</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,-469.5,446,-469.5</points>
<intersection>425.5 0</intersection>
<intersection>446 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446,-469.5,446,-464</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>-469.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-463,528.5,-463</points>
<connection>
<GID>577</GID>
<name>OUT</name></connection>
<connection>
<GID>576</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,-469,510,-449</points>
<intersection>-469 3</intersection>
<intersection>-462 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,-462,513,-462</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509,-449,510,-449</points>
<connection>
<GID>575</GID>
<name>OUT_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510,-469,530.5,-469</points>
<intersection>510 0</intersection>
<intersection>530.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530.5,-469,530.5,-466</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>-469 3</intersection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593,-463,602,-463</points>
<connection>
<GID>574</GID>
<name>OUT</name></connection>
<connection>
<GID>579</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-469,583.5,-449</points>
<intersection>-469 3</intersection>
<intersection>-462 1</intersection>
<intersection>-449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,-462,587,-462</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,-449,583.5,-449</points>
<connection>
<GID>578</GID>
<name>OUT_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583.5,-469,604,-469</points>
<intersection>583.5 0</intersection>
<intersection>604 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604,-469,604,-466</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>-469 3</intersection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,-452,576.5,-452</points>
<connection>
<GID>580</GID>
<name>OUT</name></connection>
<connection>
<GID>578</GID>
<name>clock</name></connection>
<connection>
<GID>575</GID>
<name>clock</name></connection>
<connection>
<GID>572</GID>
<name>clock</name></connection>
<connection>
<GID>569</GID>
<name>clock</name></connection>
<connection>
<GID>566</GID>
<name>clock</name></connection>
<connection>
<GID>563</GID>
<name>clock</name></connection>
<connection>
<GID>560</GID>
<name>clock</name></connection>
<connection>
<GID>557</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-786,-106,-709</points>
<intersection>-786 2</intersection>
<intersection>-727 3</intersection>
<intersection>-709 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106,-709,-2.5,-709</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-786,-106,-786</points>
<connection>
<GID>529</GID>
<name>OUT_4</name></connection>
<intersection>-106 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-106,-727,-21,-727</points>
<connection>
<GID>607</GID>
<name>ENABLE_0</name></connection>
<intersection>-106 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-18.5,-729,594,-729</points>
<connection>
<GID>607</GID>
<name>OUT_0</name></connection>
<intersection>39 38</intersection>
<intersection>113 43</intersection>
<intersection>197 42</intersection>
<intersection>271 45</intersection>
<intersection>362 47</intersection>
<intersection>436 49</intersection>
<intersection>520 51</intersection>
<intersection>594 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>39,-729,39,-716.5</points>
<connection>
<GID>585</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>197,-729,197,-718.5</points>
<connection>
<GID>591</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>113,-729,113,-716.5</points>
<connection>
<GID>582</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>271,-729,271,-718.5</points>
<connection>
<GID>588</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>362,-729,362,-720</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>436,-729,436,-720</points>
<connection>
<GID>594</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>520,-729,520,-722</points>
<connection>
<GID>603</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>594,-729,594,-722</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>-729 33</intersection></vsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-715.5,54.5,-715.5</points>
<connection>
<GID>585</GID>
<name>OUT</name></connection>
<connection>
<GID>584</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-724,36,-707</points>
<intersection>-724 3</intersection>
<intersection>-714.5 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-714.5,39,-714.5</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-707,36,-707</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-724,56.5,-724</points>
<intersection>36 0</intersection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56.5,-724,56.5,-718.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>-724 3</intersection></vsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,-715.5,128,-715.5</points>
<connection>
<GID>582</GID>
<name>OUT</name></connection>
<connection>
<GID>587</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-725.5,109.5,-707</points>
<intersection>-725.5 3</intersection>
<intersection>-714.5 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-714.5,113,-714.5</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-707,109.5,-707</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-725.5,130,-725.5</points>
<intersection>109.5 0</intersection>
<intersection>130 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130,-725.5,130,-718.5</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>-725.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,-717.5,212.5,-717.5</points>
<connection>
<GID>591</GID>
<name>OUT</name></connection>
<connection>
<GID>590</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-726,194,-707</points>
<intersection>-726 3</intersection>
<intersection>-716.5 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,-716.5,197,-716.5</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>193,-707,194,-707</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>194,-726,214.5,-726</points>
<intersection>194 0</intersection>
<intersection>214.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>214.5,-726,214.5,-720.5</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>-726 3</intersection></vsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>277,-717.5,286,-717.5</points>
<connection>
<GID>588</GID>
<name>OUT</name></connection>
<connection>
<GID>593</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-727.5,267.5,-707</points>
<connection>
<GID>592</GID>
<name>OUT_0</name></connection>
<intersection>-727.5 3</intersection>
<intersection>-716.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-716.5,271,-716.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>267.5,-727.5,288,-727.5</points>
<intersection>267.5 0</intersection>
<intersection>288 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>288,-727.5,288,-720.5</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<intersection>-727.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-719,377.5,-719</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<connection>
<GID>596</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-727.5,359,-707</points>
<intersection>-727.5 3</intersection>
<intersection>-718 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-718,362,-718</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>358,-707,359,-707</points>
<connection>
<GID>595</GID>
<name>OUT_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>359,-727.5,379.5,-727.5</points>
<intersection>359 0</intersection>
<intersection>379.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>379.5,-727.5,379.5,-722</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>-727.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>442,-719,451,-719</points>
<connection>
<GID>594</GID>
<name>OUT</name></connection>
<connection>
<GID>599</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,-727.5,432.5,-707</points>
<intersection>-727.5 3</intersection>
<intersection>-718 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,-718,436,-718</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-707,432.5,-707</points>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432.5,-727.5,453,-727.5</points>
<intersection>432.5 0</intersection>
<intersection>453 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>453,-727.5,453,-722</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>-727.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>526,-721,535.5,-721</points>
<connection>
<GID>603</GID>
<name>OUT</name></connection>
<connection>
<GID>602</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,-727,517,-707</points>
<intersection>-727 3</intersection>
<intersection>-720 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,-720,520,-720</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>516,-707,517,-707</points>
<connection>
<GID>601</GID>
<name>OUT_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>517,-727,537.5,-727</points>
<intersection>517 0</intersection>
<intersection>537.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>537.5,-727,537.5,-724</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>-727 3</intersection></vsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>600,-721,609,-721</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<connection>
<GID>605</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,-727,590.5,-707</points>
<intersection>-727 3</intersection>
<intersection>-720 1</intersection>
<intersection>-707 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,-720,594,-720</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,-707,590.5,-707</points>
<connection>
<GID>604</GID>
<name>OUT_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>590.5,-727,611,-727</points>
<intersection>590.5 0</intersection>
<intersection>611 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>611,-727,611,-724</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>-727 3</intersection></vsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-710,583.5,-710</points>
<connection>
<GID>606</GID>
<name>OUT</name></connection>
<connection>
<GID>604</GID>
<name>clock</name></connection>
<connection>
<GID>601</GID>
<name>clock</name></connection>
<connection>
<GID>598</GID>
<name>clock</name></connection>
<connection>
<GID>595</GID>
<name>clock</name></connection>
<connection>
<GID>592</GID>
<name>clock</name></connection>
<connection>
<GID>589</GID>
<name>clock</name></connection>
<connection>
<GID>586</GID>
<name>clock</name></connection>
<connection>
<GID>583</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107,-785,-107,-619</points>
<intersection>-785 2</intersection>
<intersection>-637 3</intersection>
<intersection>-619 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-107,-619,-5.5,-619</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-785,-107,-785</points>
<connection>
<GID>529</GID>
<name>OUT_5</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-107,-637,-24,-637</points>
<connection>
<GID>633</GID>
<name>ENABLE_0</name></connection>
<intersection>-107 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21.5,-639,591,-639</points>
<connection>
<GID>633</GID>
<name>OUT_0</name></connection>
<intersection>36 38</intersection>
<intersection>110 43</intersection>
<intersection>194 42</intersection>
<intersection>268 45</intersection>
<intersection>359 47</intersection>
<intersection>433 49</intersection>
<intersection>517 51</intersection>
<intersection>591 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36,-639,36,-626.5</points>
<connection>
<GID>611</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194,-639,194,-628.5</points>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110,-639,110,-626.5</points>
<connection>
<GID>608</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268,-639,268,-628.5</points>
<connection>
<GID>614</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359,-639,359,-630</points>
<connection>
<GID>623</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433,-639,433,-630</points>
<connection>
<GID>620</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517,-639,517,-632</points>
<connection>
<GID>629</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591,-639,591,-632</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<intersection>-639 33</intersection></vsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-625.5,51.5,-625.5</points>
<connection>
<GID>611</GID>
<name>OUT</name></connection>
<connection>
<GID>610</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-634,33,-617</points>
<intersection>-634 3</intersection>
<intersection>-624.5 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-624.5,36,-624.5</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-617,33,-617</points>
<connection>
<GID>609</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-634,53.5,-634</points>
<intersection>33 0</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-634,53.5,-628.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>-634 3</intersection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116,-625.5,125,-625.5</points>
<connection>
<GID>608</GID>
<name>OUT</name></connection>
<connection>
<GID>613</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-635.5,106.5,-617</points>
<intersection>-635.5 3</intersection>
<intersection>-624.5 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-624.5,110,-624.5</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-617,106.5,-617</points>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,-635.5,127,-635.5</points>
<intersection>106.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-635.5,127,-628.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>-635.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-627.5,209.5,-627.5</points>
<connection>
<GID>617</GID>
<name>OUT</name></connection>
<connection>
<GID>616</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-636,191,-617</points>
<intersection>-636 3</intersection>
<intersection>-626.5 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-626.5,194,-626.5</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,-617,191,-617</points>
<connection>
<GID>615</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191,-636,211.5,-636</points>
<intersection>191 0</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211.5,-636,211.5,-630.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>-636 3</intersection></vsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274,-627.5,283,-627.5</points>
<connection>
<GID>614</GID>
<name>OUT</name></connection>
<connection>
<GID>619</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-637.5,264.5,-617</points>
<connection>
<GID>618</GID>
<name>OUT_0</name></connection>
<intersection>-637.5 3</intersection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-626.5,268,-626.5</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264.5,-637.5,285,-637.5</points>
<intersection>264.5 0</intersection>
<intersection>285 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285,-637.5,285,-630.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>-637.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365,-629,374.5,-629</points>
<connection>
<GID>623</GID>
<name>OUT</name></connection>
<connection>
<GID>622</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-637.5,356,-617</points>
<intersection>-637.5 3</intersection>
<intersection>-628 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-628,359,-628</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355,-617,356,-617</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356,-637.5,376.5,-637.5</points>
<intersection>356 0</intersection>
<intersection>376.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376.5,-637.5,376.5,-632</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-637.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439,-629,448,-629</points>
<connection>
<GID>620</GID>
<name>OUT</name></connection>
<connection>
<GID>625</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-637.5,429.5,-617</points>
<intersection>-637.5 3</intersection>
<intersection>-628 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,-628,433,-628</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,-617,429.5,-617</points>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,-637.5,450,-637.5</points>
<intersection>429.5 0</intersection>
<intersection>450 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450,-637.5,450,-632</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>-637.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523,-631,532.5,-631</points>
<connection>
<GID>629</GID>
<name>OUT</name></connection>
<connection>
<GID>628</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-637,514,-617</points>
<intersection>-637 3</intersection>
<intersection>-630 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-630,517,-630</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,-617,514,-617</points>
<connection>
<GID>627</GID>
<name>OUT_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514,-637,534.5,-637</points>
<intersection>514 0</intersection>
<intersection>534.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534.5,-637,534.5,-634</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>-637 3</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597,-631,606,-631</points>
<connection>
<GID>626</GID>
<name>OUT</name></connection>
<connection>
<GID>631</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,-637,587.5,-617</points>
<intersection>-637 3</intersection>
<intersection>-630 1</intersection>
<intersection>-617 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,-630,591,-630</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586.5,-617,587.5,-617</points>
<connection>
<GID>630</GID>
<name>OUT_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587.5,-637,608,-637</points>
<intersection>587.5 0</intersection>
<intersection>608 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608,-637,608,-634</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>-637 3</intersection></vsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-620,580.5,-620</points>
<connection>
<GID>632</GID>
<name>OUT</name></connection>
<connection>
<GID>630</GID>
<name>clock</name></connection>
<connection>
<GID>627</GID>
<name>clock</name></connection>
<connection>
<GID>624</GID>
<name>clock</name></connection>
<connection>
<GID>621</GID>
<name>clock</name></connection>
<connection>
<GID>618</GID>
<name>clock</name></connection>
<connection>
<GID>615</GID>
<name>clock</name></connection>
<connection>
<GID>612</GID>
<name>clock</name></connection>
<connection>
<GID>609</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107,-935,-107,-788</points>
<intersection>-935 3</intersection>
<intersection>-917 1</intersection>
<intersection>-788 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-107,-917,-4.5,-917</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-788,-107,-788</points>
<connection>
<GID>529</GID>
<name>OUT_2</name></connection>
<intersection>-107 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-107,-935,-23,-935</points>
<connection>
<GID>659</GID>
<name>ENABLE_0</name></connection>
<intersection>-107 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-20.5,-937,592,-937</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>37 38</intersection>
<intersection>111 43</intersection>
<intersection>195 42</intersection>
<intersection>269 45</intersection>
<intersection>360 47</intersection>
<intersection>434 49</intersection>
<intersection>518 51</intersection>
<intersection>592 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>37,-937,37,-924.5</points>
<connection>
<GID>637</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>195,-937,195,-926.5</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>111,-937,111,-924.5</points>
<connection>
<GID>634</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>269,-937,269,-926.5</points>
<connection>
<GID>640</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>360,-937,360,-928</points>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>434,-937,434,-928</points>
<connection>
<GID>646</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>518,-937,518,-930</points>
<connection>
<GID>655</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>592,-937,592,-930</points>
<connection>
<GID>652</GID>
<name>IN_1</name></connection>
<intersection>-937 33</intersection></vsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-923.5,52.5,-923.5</points>
<connection>
<GID>637</GID>
<name>OUT</name></connection>
<connection>
<GID>636</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-932,34,-915</points>
<intersection>-932 3</intersection>
<intersection>-922.5 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-922.5,37,-922.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-915,34,-915</points>
<connection>
<GID>635</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-932,54.5,-932</points>
<intersection>34 0</intersection>
<intersection>54.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54.5,-932,54.5,-926.5</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>-932 3</intersection></vsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>117,-923.5,127,-923.5</points>
<connection>
<GID>634</GID>
<name>OUT</name></connection>
<connection>
<GID>639</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-933.5,107.5,-915</points>
<intersection>-933.5 3</intersection>
<intersection>-922.5 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-922.5,111,-922.5</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-915,107.5,-915</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-933.5,129,-933.5</points>
<intersection>107.5 0</intersection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-933.5,129,-926.5</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>-933.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201,-925.5,210.5,-925.5</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<connection>
<GID>642</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-934,192,-915</points>
<intersection>-934 3</intersection>
<intersection>-924.5 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-924.5,195,-924.5</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-915,192,-915</points>
<connection>
<GID>641</GID>
<name>OUT_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>192,-934,212.5,-934</points>
<intersection>192 0</intersection>
<intersection>212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>212.5,-934,212.5,-928.5</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>-934 3</intersection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>275,-925.5,284,-925.5</points>
<connection>
<GID>640</GID>
<name>OUT</name></connection>
<connection>
<GID>645</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-935.5,265.5,-915</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>-935.5 3</intersection>
<intersection>-924.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,-924.5,269,-924.5</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>265.5,-935.5,286,-935.5</points>
<intersection>265.5 0</intersection>
<intersection>286 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>286,-935.5,286,-928.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>-935.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366,-927,375.5,-927</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<connection>
<GID>648</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-935.5,357,-915</points>
<intersection>-935.5 3</intersection>
<intersection>-926 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-926,360,-926</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356,-915,357,-915</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-935.5,377.5,-935.5</points>
<intersection>357 0</intersection>
<intersection>377.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>377.5,-935.5,377.5,-930</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-935.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>440,-927,449,-927</points>
<connection>
<GID>646</GID>
<name>OUT</name></connection>
<connection>
<GID>651</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,-935.5,430.5,-915</points>
<intersection>-935.5 3</intersection>
<intersection>-926 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430.5,-926,434,-926</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>429.5,-915,430.5,-915</points>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>430.5,-935.5,451,-935.5</points>
<intersection>430.5 0</intersection>
<intersection>451 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>451,-935.5,451,-930</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-935.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524,-929,533.5,-929</points>
<connection>
<GID>655</GID>
<name>OUT</name></connection>
<connection>
<GID>654</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-935,515,-915</points>
<intersection>-935 3</intersection>
<intersection>-928 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515,-928,518,-928</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,-915,515,-915</points>
<connection>
<GID>653</GID>
<name>OUT_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>515,-935,535.5,-935</points>
<intersection>515 0</intersection>
<intersection>535.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535.5,-935,535.5,-932</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>-935 3</intersection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>598,-929,607,-929</points>
<connection>
<GID>652</GID>
<name>OUT</name></connection>
<connection>
<GID>657</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588.5,-935,588.5,-915</points>
<intersection>-935 3</intersection>
<intersection>-928 1</intersection>
<intersection>-915 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588.5,-928,592,-928</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-915,588.5,-915</points>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>588.5,-935,609,-935</points>
<intersection>588.5 0</intersection>
<intersection>609 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>609,-935,609,-932</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>-935 3</intersection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-918,581.5,-918</points>
<connection>
<GID>658</GID>
<name>OUT</name></connection>
<connection>
<GID>656</GID>
<name>clock</name></connection>
<connection>
<GID>653</GID>
<name>clock</name></connection>
<connection>
<GID>650</GID>
<name>clock</name></connection>
<connection>
<GID>647</GID>
<name>clock</name></connection>
<connection>
<GID>644</GID>
<name>clock</name></connection>
<connection>
<GID>641</GID>
<name>clock</name></connection>
<connection>
<GID>638</GID>
<name>clock</name></connection>
<connection>
<GID>635</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-845,-106,-787</points>
<intersection>-845 3</intersection>
<intersection>-827 1</intersection>
<intersection>-787 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106,-827,-7.5,-827</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>-106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-787,-106,-787</points>
<connection>
<GID>529</GID>
<name>OUT_3</name></connection>
<intersection>-106 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-106,-845,-26,-845</points>
<connection>
<GID>476</GID>
<name>ENABLE_0</name></connection>
<intersection>-106 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-847,589,-847</points>
<connection>
<GID>476</GID>
<name>OUT_0</name></connection>
<intersection>34 38</intersection>
<intersection>108 43</intersection>
<intersection>192 42</intersection>
<intersection>266 45</intersection>
<intersection>357 47</intersection>
<intersection>431 49</intersection>
<intersection>515 51</intersection>
<intersection>589 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34,-847,34,-834.5</points>
<connection>
<GID>663</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192,-847,192,-836.5</points>
<connection>
<GID>460</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108,-847,108,-834.5</points>
<connection>
<GID>660</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266,-847,266,-836.5</points>
<connection>
<GID>666</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357,-847,357,-838</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431,-847,431,-838</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515,-847,515,-840</points>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589,-847,589,-840</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>-847 33</intersection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-833.5,49.5,-833.5</points>
<connection>
<GID>663</GID>
<name>OUT</name></connection>
<connection>
<GID>662</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-842,31,-825</points>
<intersection>-842 3</intersection>
<intersection>-832.5 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-832.5,34,-832.5</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-825,31,-825</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-842,51.5,-842</points>
<intersection>31 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-842,51.5,-836.5</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>-842 3</intersection></vsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114,-833.5,123,-833.5</points>
<connection>
<GID>660</GID>
<name>OUT</name></connection>
<connection>
<GID>665</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-843.5,104.5,-825</points>
<intersection>-843.5 3</intersection>
<intersection>-832.5 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-832.5,108,-832.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-825,104.5,-825</points>
<connection>
<GID>664</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-843.5,125,-843.5</points>
<intersection>104.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-843.5,125,-836.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>-843.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-835.5,207.5,-835.5</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<connection>
<GID>668</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-844,189,-825</points>
<intersection>-844 3</intersection>
<intersection>-834.5 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-834.5,192,-834.5</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188,-825,189,-825</points>
<connection>
<GID>667</GID>
<name>OUT_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189,-844,209.5,-844</points>
<intersection>189 0</intersection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,-844,209.5,-838.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-844 3</intersection></vsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272,-835.5,281,-835.5</points>
<connection>
<GID>666</GID>
<name>OUT</name></connection>
<connection>
<GID>462</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-845.5,262.5,-825</points>
<connection>
<GID>461</GID>
<name>OUT_0</name></connection>
<intersection>-845.5 3</intersection>
<intersection>-834.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-834.5,266,-834.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262.5,-845.5,283,-845.5</points>
<intersection>262.5 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-845.5,283,-838.5</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>-845.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363,-837,372.5,-837</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<connection>
<GID>465</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-845.5,354,-825</points>
<intersection>-845.5 3</intersection>
<intersection>-836 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-836,357,-836</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-825,354,-825</points>
<connection>
<GID>464</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354,-845.5,374.5,-845.5</points>
<intersection>354 0</intersection>
<intersection>374.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374.5,-845.5,374.5,-840</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-845.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437,-837,446,-837</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<connection>
<GID>468</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-845.5,427.5,-825</points>
<intersection>-845.5 3</intersection>
<intersection>-836 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-836,431,-836</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426.5,-825,427.5,-825</points>
<connection>
<GID>467</GID>
<name>OUT_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-845.5,448,-845.5</points>
<intersection>427.5 0</intersection>
<intersection>448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448,-845.5,448,-840</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>-845.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521,-839,530.5,-839</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<connection>
<GID>471</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,-845,512,-825</points>
<intersection>-845 3</intersection>
<intersection>-838 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-838,515,-838</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,-825,512,-825</points>
<connection>
<GID>470</GID>
<name>OUT_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512,-845,532.5,-845</points>
<intersection>512 0</intersection>
<intersection>532.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532.5,-845,532.5,-842</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>-845 3</intersection></vsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595,-839,604,-839</points>
<connection>
<GID>469</GID>
<name>OUT</name></connection>
<connection>
<GID>474</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-845,585.5,-825</points>
<intersection>-845 3</intersection>
<intersection>-838 1</intersection>
<intersection>-825 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-838,589,-838</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,-825,585.5,-825</points>
<connection>
<GID>473</GID>
<name>OUT_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-845,606,-845</points>
<intersection>585.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-845,606,-842</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>-845 3</intersection></vsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-828,578.5,-828</points>
<connection>
<GID>667</GID>
<name>clock</name></connection>
<connection>
<GID>664</GID>
<name>clock</name></connection>
<connection>
<GID>661</GID>
<name>clock</name></connection>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<connection>
<GID>473</GID>
<name>clock</name></connection>
<connection>
<GID>470</GID>
<name>clock</name></connection>
<connection>
<GID>467</GID>
<name>clock</name></connection>
<connection>
<GID>464</GID>
<name>clock</name></connection>
<connection>
<GID>461</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-1103,-110,-790</points>
<intersection>-1103 3</intersection>
<intersection>-1085 1</intersection>
<intersection>-790 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-1085,-0.5,-1085</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-790,-110,-790</points>
<connection>
<GID>529</GID>
<name>OUT_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-1103,-19,-1103</points>
<connection>
<GID>502</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-16.5,-1105,596,-1105</points>
<connection>
<GID>502</GID>
<name>OUT_0</name></connection>
<intersection>41 38</intersection>
<intersection>115 43</intersection>
<intersection>199 42</intersection>
<intersection>273 45</intersection>
<intersection>364 47</intersection>
<intersection>438 49</intersection>
<intersection>522 51</intersection>
<intersection>596 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>41,-1105,41,-1092.5</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>199,-1105,199,-1094.5</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>115,-1105,115,-1092.5</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>273,-1105,273,-1094.5</points>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>364,-1105,364,-1096</points>
<connection>
<GID>492</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>438,-1105,438,-1096</points>
<connection>
<GID>489</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>522,-1105,522,-1098</points>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>596,-1105,596,-1098</points>
<connection>
<GID>495</GID>
<name>IN_1</name></connection>
<intersection>-1105 33</intersection></vsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-1091.5,56.5,-1091.5</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>479</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-1100,38,-1083</points>
<intersection>-1100 3</intersection>
<intersection>-1090.5 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-1090.5,41,-1090.5</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-1083,38,-1083</points>
<connection>
<GID>478</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-1100,58.5,-1100</points>
<intersection>38 0</intersection>
<intersection>58.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>58.5,-1100,58.5,-1094.5</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>-1100 3</intersection></vsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>121,-1091.5,130,-1091.5</points>
<connection>
<GID>477</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-1101.5,111.5,-1083</points>
<intersection>-1101.5 3</intersection>
<intersection>-1090.5 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-1090.5,115,-1090.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-1083,111.5,-1083</points>
<connection>
<GID>481</GID>
<name>OUT_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>111.5,-1101.5,132,-1101.5</points>
<intersection>111.5 0</intersection>
<intersection>132 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132,-1101.5,132,-1094.5</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>-1101.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-1093.5,214.5,-1093.5</points>
<connection>
<GID>486</GID>
<name>OUT</name></connection>
<connection>
<GID>485</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-1102,196,-1083</points>
<intersection>-1102 3</intersection>
<intersection>-1092.5 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196,-1092.5,199,-1092.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,-1083,196,-1083</points>
<connection>
<GID>484</GID>
<name>OUT_0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>196,-1102,216.5,-1102</points>
<intersection>196 0</intersection>
<intersection>216.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>216.5,-1102,216.5,-1096.5</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>-1102 3</intersection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>279,-1093.5,288,-1093.5</points>
<connection>
<GID>483</GID>
<name>OUT</name></connection>
<connection>
<GID>488</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-1103.5,269.5,-1083</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<intersection>-1103.5 3</intersection>
<intersection>-1092.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,-1092.5,273,-1092.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>269.5,-1103.5,290,-1103.5</points>
<intersection>269.5 0</intersection>
<intersection>290 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>290,-1103.5,290,-1096.5</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-1103.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>370,-1095,379.5,-1095</points>
<connection>
<GID>492</GID>
<name>OUT</name></connection>
<connection>
<GID>491</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-1103.5,361,-1083</points>
<intersection>-1103.5 3</intersection>
<intersection>-1094 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-1094,364,-1094</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>360,-1083,361,-1083</points>
<connection>
<GID>490</GID>
<name>OUT_0</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>361,-1103.5,381.5,-1103.5</points>
<intersection>361 0</intersection>
<intersection>381.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>381.5,-1103.5,381.5,-1098</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>-1103.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>444,-1095,453,-1095</points>
<connection>
<GID>489</GID>
<name>OUT</name></connection>
<connection>
<GID>494</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-1103.5,434.5,-1083</points>
<intersection>-1103.5 3</intersection>
<intersection>-1094 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-1094,438,-1094</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-1083,434.5,-1083</points>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>434.5,-1103.5,455,-1103.5</points>
<intersection>434.5 0</intersection>
<intersection>455 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>455,-1103.5,455,-1098</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>-1103.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>528,-1097,537.5,-1097</points>
<connection>
<GID>498</GID>
<name>OUT</name></connection>
<connection>
<GID>497</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519,-1103,519,-1083</points>
<intersection>-1103 3</intersection>
<intersection>-1096 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>519,-1096,522,-1096</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>519 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>518,-1083,519,-1083</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<intersection>519 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>519,-1103,539.5,-1103</points>
<intersection>519 0</intersection>
<intersection>539.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>539.5,-1103,539.5,-1100</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>-1103 3</intersection></vsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>602,-1097,611,-1097</points>
<connection>
<GID>495</GID>
<name>OUT</name></connection>
<connection>
<GID>500</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-1103,592.5,-1083</points>
<intersection>-1103 3</intersection>
<intersection>-1096 1</intersection>
<intersection>-1083 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-1096,596,-1096</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>591.5,-1083,592.5,-1083</points>
<connection>
<GID>499</GID>
<name>OUT_0</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>592.5,-1103,613,-1103</points>
<intersection>592.5 0</intersection>
<intersection>613 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>613,-1103,613,-1100</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-1103 3</intersection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-1086,585.5,-1086</points>
<connection>
<GID>501</GID>
<name>OUT</name></connection>
<connection>
<GID>499</GID>
<name>clock</name></connection>
<connection>
<GID>496</GID>
<name>clock</name></connection>
<connection>
<GID>493</GID>
<name>clock</name></connection>
<connection>
<GID>490</GID>
<name>clock</name></connection>
<connection>
<GID>487</GID>
<name>clock</name></connection>
<connection>
<GID>484</GID>
<name>clock</name></connection>
<connection>
<GID>481</GID>
<name>clock</name></connection>
<connection>
<GID>478</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-1013,-108,-789</points>
<intersection>-1013 3</intersection>
<intersection>-995 1</intersection>
<intersection>-789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-995,-3.5,-995</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-789,-108,-789</points>
<connection>
<GID>529</GID>
<name>OUT_1</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-1013,-22,-1013</points>
<connection>
<GID>528</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-19.5,-1015,593,-1015</points>
<connection>
<GID>528</GID>
<name>OUT_0</name></connection>
<intersection>38 38</intersection>
<intersection>112 43</intersection>
<intersection>196 42</intersection>
<intersection>270 45</intersection>
<intersection>361 47</intersection>
<intersection>435 49</intersection>
<intersection>519 51</intersection>
<intersection>593 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>38,-1015,38,-1002.5</points>
<connection>
<GID>506</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>196,-1015,196,-1004.5</points>
<connection>
<GID>512</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>112,-1015,112,-1002.5</points>
<connection>
<GID>503</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>270,-1015,270,-1004.5</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>361,-1015,361,-1006</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>435,-1015,435,-1006</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>519,-1015,519,-1008</points>
<connection>
<GID>524</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>593,-1015,593,-1008</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>-1015 33</intersection></vsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-1001.5,53.5,-1001.5</points>
<connection>
<GID>506</GID>
<name>OUT</name></connection>
<connection>
<GID>505</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-1010,35,-993</points>
<intersection>-1010 3</intersection>
<intersection>-1000.5 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-1000.5,38,-1000.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-993,35,-993</points>
<connection>
<GID>504</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-1010,55.5,-1010</points>
<intersection>35 0</intersection>
<intersection>55.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55.5,-1010,55.5,-1004.5</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>-1010 3</intersection></vsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>118,-1001.5,127,-1001.5</points>
<connection>
<GID>503</GID>
<name>OUT</name></connection>
<connection>
<GID>508</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-1011.5,108.5,-993</points>
<intersection>-1011.5 3</intersection>
<intersection>-1000.5 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-1000.5,112,-1000.5</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-993,108.5,-993</points>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108.5,-1011.5,129,-1011.5</points>
<intersection>108.5 0</intersection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-1011.5,129,-1004.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>-1011.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-1003.5,211.5,-1003.5</points>
<connection>
<GID>512</GID>
<name>OUT</name></connection>
<connection>
<GID>511</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-1012,193,-993</points>
<intersection>-1012 3</intersection>
<intersection>-1002.5 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-1002.5,196,-1002.5</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>192,-993,193,-993</points>
<connection>
<GID>510</GID>
<name>OUT_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>193,-1012,213.5,-1012</points>
<intersection>193 0</intersection>
<intersection>213.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>213.5,-1012,213.5,-1006.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>-1012 3</intersection></vsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>276,-1003.5,285,-1003.5</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<connection>
<GID>514</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-1013.5,266.5,-993</points>
<connection>
<GID>513</GID>
<name>OUT_0</name></connection>
<intersection>-1013.5 3</intersection>
<intersection>-1002.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-1002.5,270,-1002.5</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-1013.5,287,-1013.5</points>
<intersection>266.5 0</intersection>
<intersection>287 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>287,-1013.5,287,-1006.5</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>-1013.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367,-1005,376.5,-1005</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<connection>
<GID>517</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358,-1013.5,358,-993</points>
<intersection>-1013.5 3</intersection>
<intersection>-1004 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358,-1004,361,-1004</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-993,358,-993</points>
<connection>
<GID>516</GID>
<name>OUT_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>358,-1013.5,378.5,-1013.5</points>
<intersection>358 0</intersection>
<intersection>378.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>378.5,-1013.5,378.5,-1008</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>-1013.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>441,-1005,450,-1005</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<connection>
<GID>520</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,-1013.5,431.5,-993</points>
<intersection>-1013.5 3</intersection>
<intersection>-1004 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,-1004,435,-1004</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>430.5,-993,431.5,-993</points>
<connection>
<GID>519</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>431.5,-1013.5,452,-1013.5</points>
<intersection>431.5 0</intersection>
<intersection>452 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>452,-1013.5,452,-1008</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>-1013.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>525,-1007,534.5,-1007</points>
<connection>
<GID>524</GID>
<name>OUT</name></connection>
<connection>
<GID>523</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,-1013,516,-993</points>
<intersection>-1013 3</intersection>
<intersection>-1006 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,-1006,519,-1006</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515,-993,516,-993</points>
<connection>
<GID>522</GID>
<name>OUT_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>516,-1013,536.5,-1013</points>
<intersection>516 0</intersection>
<intersection>536.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>536.5,-1013,536.5,-1010</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>-1013 3</intersection></vsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>599,-1007,608,-1007</points>
<connection>
<GID>521</GID>
<name>OUT</name></connection>
<connection>
<GID>526</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-1013,589.5,-993</points>
<intersection>-1013 3</intersection>
<intersection>-1006 1</intersection>
<intersection>-993 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589.5,-1006,593,-1006</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-993,589.5,-993</points>
<connection>
<GID>525</GID>
<name>OUT_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>589.5,-1013,610,-1013</points>
<intersection>589.5 0</intersection>
<intersection>610 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>610,-1013,610,-1010</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>-1013 3</intersection></vsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-996,582.5,-996</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<connection>
<GID>525</GID>
<name>clock</name></connection>
<connection>
<GID>522</GID>
<name>clock</name></connection>
<connection>
<GID>519</GID>
<name>clock</name></connection>
<connection>
<GID>516</GID>
<name>clock</name></connection>
<connection>
<GID>513</GID>
<name>clock</name></connection>
<connection>
<GID>510</GID>
<name>clock</name></connection>
<connection>
<GID>507</GID>
<name>clock</name></connection>
<connection>
<GID>504</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110.5,-1708.5,-110.5,-1465.5</points>
<intersection>-1708.5 2</intersection>
<intersection>-1483.5 3</intersection>
<intersection>-1465.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-1465.5,-9,-1465.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1708.5,-110.5,-1708.5</points>
<connection>
<GID>738</GID>
<name>OUT_6</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110.5,-1483.5,-27.5,-1483.5</points>
<connection>
<GID>764</GID>
<name>ENABLE_0</name></connection>
<intersection>-110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25,-1485.5,587.5,-1485.5</points>
<connection>
<GID>764</GID>
<name>OUT_0</name></connection>
<intersection>32.5 38</intersection>
<intersection>106.5 43</intersection>
<intersection>190.5 42</intersection>
<intersection>264.5 45</intersection>
<intersection>355.5 47</intersection>
<intersection>429.5 49</intersection>
<intersection>513.5 51</intersection>
<intersection>587.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32.5,-1485.5,32.5,-1473</points>
<connection>
<GID>742</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190.5,-1485.5,190.5,-1475</points>
<connection>
<GID>748</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106.5,-1485.5,106.5,-1473</points>
<connection>
<GID>739</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264.5,-1485.5,264.5,-1475</points>
<connection>
<GID>745</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355.5,-1485.5,355.5,-1476.5</points>
<connection>
<GID>754</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429.5,-1485.5,429.5,-1476.5</points>
<connection>
<GID>751</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513.5,-1485.5,513.5,-1478.5</points>
<connection>
<GID>760</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587.5,-1485.5,587.5,-1478.5</points>
<connection>
<GID>757</GID>
<name>IN_1</name></connection>
<intersection>-1485.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-1472,48,-1472</points>
<connection>
<GID>742</GID>
<name>OUT</name></connection>
<connection>
<GID>741</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-1480.5,29.5,-1463.5</points>
<intersection>-1480.5 3</intersection>
<intersection>-1471 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-1471,32.5,-1471</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-1463.5,29.5,-1463.5</points>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-1480.5,50,-1480.5</points>
<intersection>29.5 0</intersection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,-1480.5,50,-1475</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-1480.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112.5,-1472,121.5,-1472</points>
<connection>
<GID>744</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>739</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-1482,103,-1463.5</points>
<intersection>-1482 3</intersection>
<intersection>-1471 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-1471,106.5,-1471</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-1463.5,103,-1463.5</points>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,-1482,123.5,-1482</points>
<intersection>103 0</intersection>
<intersection>123.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123.5,-1482,123.5,-1475</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>-1482 3</intersection></vsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,-1474,206,-1474</points>
<connection>
<GID>748</GID>
<name>OUT</name></connection>
<connection>
<GID>747</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-1482.5,187.5,-1463.5</points>
<intersection>-1482.5 3</intersection>
<intersection>-1473 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,-1473,190.5,-1473</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186.5,-1463.5,187.5,-1463.5</points>
<connection>
<GID>746</GID>
<name>OUT_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-1482.5,208,-1482.5</points>
<intersection>187.5 0</intersection>
<intersection>208 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208,-1482.5,208,-1477</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>-1482.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270.5,-1474,279.5,-1474</points>
<connection>
<GID>750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>745</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-1484,261,-1463.5</points>
<connection>
<GID>749</GID>
<name>OUT_0</name></connection>
<intersection>-1484 3</intersection>
<intersection>-1473 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-1473,264.5,-1473</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>261,-1484,281.5,-1484</points>
<intersection>261 0</intersection>
<intersection>281.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281.5,-1484,281.5,-1477</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>-1484 3</intersection></vsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361.5,-1475.5,371,-1475.5</points>
<connection>
<GID>754</GID>
<name>OUT</name></connection>
<connection>
<GID>753</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352.5,-1484,352.5,-1463.5</points>
<intersection>-1484 3</intersection>
<intersection>-1474.5 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352.5,-1474.5,355.5,-1474.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>352.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351.5,-1463.5,352.5,-1463.5</points>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection>
<intersection>352.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352.5,-1484,373,-1484</points>
<intersection>352.5 0</intersection>
<intersection>373 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>373,-1484,373,-1478.5</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>-1484 3</intersection></vsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435.5,-1475.5,444.5,-1475.5</points>
<connection>
<GID>756</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>751</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,-1484,426,-1463.5</points>
<intersection>-1484 3</intersection>
<intersection>-1474.5 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426,-1474.5,429.5,-1474.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425,-1463.5,426,-1463.5</points>
<connection>
<GID>755</GID>
<name>OUT_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426,-1484,446.5,-1484</points>
<intersection>426 0</intersection>
<intersection>446.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446.5,-1484,446.5,-1478.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>-1484 3</intersection></vsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519.5,-1477.5,529,-1477.5</points>
<connection>
<GID>760</GID>
<name>OUT</name></connection>
<connection>
<GID>759</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510.5,-1483.5,510.5,-1463.5</points>
<intersection>-1483.5 3</intersection>
<intersection>-1476.5 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,-1476.5,513.5,-1476.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>510.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509.5,-1463.5,510.5,-1463.5</points>
<connection>
<GID>758</GID>
<name>OUT_0</name></connection>
<intersection>510.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510.5,-1483.5,531,-1483.5</points>
<intersection>510.5 0</intersection>
<intersection>531 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531,-1483.5,531,-1480.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>-1483.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593.5,-1477.5,602.5,-1477.5</points>
<connection>
<GID>762</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>757</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584,-1483.5,584,-1463.5</points>
<intersection>-1483.5 3</intersection>
<intersection>-1476.5 1</intersection>
<intersection>-1463.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584,-1476.5,587.5,-1476.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>584 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583,-1463.5,584,-1463.5</points>
<connection>
<GID>761</GID>
<name>OUT_0</name></connection>
<intersection>584 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>584,-1483.5,604.5,-1483.5</points>
<intersection>584 0</intersection>
<intersection>604.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604.5,-1483.5,604.5,-1480.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>-1483.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3,-1466.5,577,-1466.5</points>
<connection>
<GID>763</GID>
<name>OUT</name></connection>
<connection>
<GID>761</GID>
<name>clock</name></connection>
<connection>
<GID>758</GID>
<name>clock</name></connection>
<connection>
<GID>755</GID>
<name>clock</name></connection>
<connection>
<GID>752</GID>
<name>clock</name></connection>
<connection>
<GID>749</GID>
<name>clock</name></connection>
<connection>
<GID>746</GID>
<name>clock</name></connection>
<connection>
<GID>743</GID>
<name>clock</name></connection>
<connection>
<GID>740</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111.5,-1707.5,-111.5,-1375.5</points>
<intersection>-1707.5 2</intersection>
<intersection>-1393.5 3</intersection>
<intersection>-1375.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111.5,-1375.5,-12,-1375.5</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1707.5,-111.5,-1707.5</points>
<connection>
<GID>738</GID>
<name>OUT_7</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111.5,-1393.5,-26,-1393.5</points>
<intersection>-111.5 0</intersection>
<intersection>-26 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-26,-1394,-26,-1393.5</points>
<connection>
<GID>790</GID>
<name>ENABLE_0</name></connection>
<intersection>-1393.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-1396,584.5,-1396</points>
<connection>
<GID>790</GID>
<name>OUT_0</name></connection>
<intersection>29.5 38</intersection>
<intersection>103.5 43</intersection>
<intersection>187.5 42</intersection>
<intersection>261.5 45</intersection>
<intersection>352.5 47</intersection>
<intersection>426.5 49</intersection>
<intersection>510.5 51</intersection>
<intersection>584.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>29.5,-1396,29.5,-1383</points>
<connection>
<GID>768</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>187.5,-1396,187.5,-1385</points>
<connection>
<GID>774</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>103.5,-1396,103.5,-1383</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>261.5,-1396,261.5,-1385</points>
<connection>
<GID>771</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>352.5,-1396,352.5,-1386.5</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>426.5,-1396,426.5,-1386.5</points>
<connection>
<GID>777</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>510.5,-1396,510.5,-1388.5</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>584.5,-1396,584.5,-1388.5</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>-1396 33</intersection></vsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-1382,45,-1382</points>
<connection>
<GID>768</GID>
<name>OUT</name></connection>
<connection>
<GID>767</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-1390.5,26.5,-1373.5</points>
<intersection>-1390.5 3</intersection>
<intersection>-1381 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-1381,29.5,-1381</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-1373.5,26.5,-1373.5</points>
<connection>
<GID>766</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-1390.5,47,-1390.5</points>
<intersection>26.5 0</intersection>
<intersection>47 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>47,-1390.5,47,-1385</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>-1390.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>109.5,-1382,118.5,-1382</points>
<connection>
<GID>765</GID>
<name>OUT</name></connection>
<connection>
<GID>770</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-1392,100,-1373.5</points>
<intersection>-1392 3</intersection>
<intersection>-1381 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-1381,103.5,-1381</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-1373.5,100,-1373.5</points>
<connection>
<GID>769</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100,-1392,120.5,-1392</points>
<intersection>100 0</intersection>
<intersection>120.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>120.5,-1392,120.5,-1385</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-1392 3</intersection></vsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>193.5,-1384,203,-1384</points>
<connection>
<GID>774</GID>
<name>OUT</name></connection>
<connection>
<GID>773</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-1392.5,184.5,-1373.5</points>
<intersection>-1392.5 3</intersection>
<intersection>-1383 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-1383,187.5,-1383</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-1373.5,184.5,-1373.5</points>
<connection>
<GID>772</GID>
<name>OUT_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184.5,-1392.5,205,-1392.5</points>
<intersection>184.5 0</intersection>
<intersection>205 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>205,-1392.5,205,-1387</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>-1392.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>267.5,-1384,276.5,-1384</points>
<connection>
<GID>776</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>771</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-1394,258,-1373.5</points>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection>
<intersection>-1394 3</intersection>
<intersection>-1383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-1383,261.5,-1383</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258,-1394,278.5,-1394</points>
<intersection>258 0</intersection>
<intersection>278.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>278.5,-1394,278.5,-1387</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-1394 3</intersection></vsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358.5,-1385.5,368,-1385.5</points>
<connection>
<GID>780</GID>
<name>OUT</name></connection>
<connection>
<GID>779</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-1394,349.5,-1373.5</points>
<intersection>-1394 3</intersection>
<intersection>-1384.5 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349.5,-1384.5,352.5,-1384.5</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,-1373.5,349.5,-1373.5</points>
<connection>
<GID>778</GID>
<name>OUT_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>349.5,-1394,370,-1394</points>
<intersection>349.5 0</intersection>
<intersection>370 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>370,-1394,370,-1388.5</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-1394 3</intersection></vsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>432.5,-1385.5,441.5,-1385.5</points>
<connection>
<GID>782</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>777</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423,-1394,423,-1373.5</points>
<intersection>-1394 3</intersection>
<intersection>-1384.5 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,-1384.5,426.5,-1384.5</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>423 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422,-1373.5,423,-1373.5</points>
<connection>
<GID>781</GID>
<name>OUT_0</name></connection>
<intersection>423 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>423,-1394,443.5,-1394</points>
<intersection>423 0</intersection>
<intersection>443.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>443.5,-1394,443.5,-1388.5</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-1394 3</intersection></vsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>516.5,-1387.5,526,-1387.5</points>
<connection>
<GID>786</GID>
<name>OUT</name></connection>
<connection>
<GID>785</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507.5,-1393.5,507.5,-1373.5</points>
<intersection>-1393.5 3</intersection>
<intersection>-1386.5 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507.5,-1386.5,510.5,-1386.5</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>507.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>506.5,-1373.5,507.5,-1373.5</points>
<connection>
<GID>784</GID>
<name>OUT_0</name></connection>
<intersection>507.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>507.5,-1393.5,528,-1393.5</points>
<intersection>507.5 0</intersection>
<intersection>528 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>528,-1393.5,528,-1390.5</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>-1393.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>590.5,-1387.5,599.5,-1387.5</points>
<connection>
<GID>788</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>783</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,-1393.5,581,-1373.5</points>
<intersection>-1393.5 3</intersection>
<intersection>-1386.5 1</intersection>
<intersection>-1373.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581,-1386.5,584.5,-1386.5</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>581 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>580,-1373.5,581,-1373.5</points>
<connection>
<GID>787</GID>
<name>OUT_0</name></connection>
<intersection>581 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>581,-1393.5,601.5,-1393.5</points>
<intersection>581 0</intersection>
<intersection>601.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>601.5,-1393.5,601.5,-1390.5</points>
<connection>
<GID>788</GID>
<name>IN_0</name></connection>
<intersection>-1393.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-1376.5,574,-1376.5</points>
<connection>
<GID>766</GID>
<name>clock</name></connection>
<connection>
<GID>789</GID>
<name>OUT</name></connection>
<connection>
<GID>787</GID>
<name>clock</name></connection>
<connection>
<GID>784</GID>
<name>clock</name></connection>
<connection>
<GID>781</GID>
<name>clock</name></connection>
<connection>
<GID>778</GID>
<name>clock</name></connection>
<connection>
<GID>775</GID>
<name>clock</name></connection>
<connection>
<GID>772</GID>
<name>clock</name></connection>
<connection>
<GID>769</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108.5,-1710.5,-108.5,-1633.5</points>
<intersection>-1710.5 2</intersection>
<intersection>-1651.5 3</intersection>
<intersection>-1633.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108.5,-1633.5,-5,-1633.5</points>
<connection>
<GID>815</GID>
<name>IN_0</name></connection>
<intersection>-108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1710.5,-108.5,-1710.5</points>
<connection>
<GID>738</GID>
<name>OUT_4</name></connection>
<intersection>-108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108.5,-1651.5,-23.5,-1651.5</points>
<connection>
<GID>816</GID>
<name>ENABLE_0</name></connection>
<intersection>-108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21,-1653.5,591.5,-1653.5</points>
<connection>
<GID>816</GID>
<name>OUT_0</name></connection>
<intersection>36.5 38</intersection>
<intersection>110.5 43</intersection>
<intersection>194.5 42</intersection>
<intersection>268.5 45</intersection>
<intersection>359.5 47</intersection>
<intersection>433.5 49</intersection>
<intersection>517.5 51</intersection>
<intersection>591.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36.5,-1653.5,36.5,-1641</points>
<connection>
<GID>794</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194.5,-1653.5,194.5,-1643</points>
<connection>
<GID>800</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110.5,-1653.5,110.5,-1641</points>
<connection>
<GID>791</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268.5,-1653.5,268.5,-1643</points>
<connection>
<GID>797</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359.5,-1653.5,359.5,-1644.5</points>
<connection>
<GID>806</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433.5,-1653.5,433.5,-1644.5</points>
<connection>
<GID>803</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517.5,-1653.5,517.5,-1646.5</points>
<connection>
<GID>812</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591.5,-1653.5,591.5,-1646.5</points>
<connection>
<GID>809</GID>
<name>IN_1</name></connection>
<intersection>-1653.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-1640,52,-1640</points>
<connection>
<GID>794</GID>
<name>OUT</name></connection>
<connection>
<GID>793</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-1648.5,33.5,-1631.5</points>
<intersection>-1648.5 3</intersection>
<intersection>-1639 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-1639,36.5,-1639</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-1631.5,33.5,-1631.5</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-1648.5,54,-1648.5</points>
<intersection>33.5 0</intersection>
<intersection>54 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54,-1648.5,54,-1643</points>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>-1648.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116.5,-1640,125.5,-1640</points>
<connection>
<GID>796</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>791</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-1650,107,-1631.5</points>
<intersection>-1650 3</intersection>
<intersection>-1639 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-1639,110.5,-1639</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,-1631.5,107,-1631.5</points>
<connection>
<GID>795</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107,-1650,127.5,-1650</points>
<intersection>107 0</intersection>
<intersection>127.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127.5,-1650,127.5,-1643</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>-1650 3</intersection></vsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,-1642,210,-1642</points>
<connection>
<GID>800</GID>
<name>OUT</name></connection>
<connection>
<GID>799</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-1650.5,191.5,-1631.5</points>
<intersection>-1650.5 3</intersection>
<intersection>-1641 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-1641,194.5,-1641</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190.5,-1631.5,191.5,-1631.5</points>
<connection>
<GID>798</GID>
<name>OUT_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191.5,-1650.5,212,-1650.5</points>
<intersection>191.5 0</intersection>
<intersection>212 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>212,-1650.5,212,-1645</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>-1650.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274.5,-1642,283.5,-1642</points>
<connection>
<GID>797</GID>
<name>OUT</name></connection>
<connection>
<GID>802</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265,-1652,265,-1631.5</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<intersection>-1652 3</intersection>
<intersection>-1641 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265,-1641,268.5,-1641</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>265 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>265,-1652,285.5,-1652</points>
<intersection>265 0</intersection>
<intersection>285.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285.5,-1652,285.5,-1645</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<intersection>-1652 3</intersection></vsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365.5,-1643.5,375,-1643.5</points>
<connection>
<GID>806</GID>
<name>OUT</name></connection>
<connection>
<GID>805</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,-1652,356.5,-1631.5</points>
<intersection>-1652 3</intersection>
<intersection>-1642.5 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356.5,-1642.5,359.5,-1642.5</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355.5,-1631.5,356.5,-1631.5</points>
<connection>
<GID>804</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356.5,-1652,377,-1652</points>
<intersection>356.5 0</intersection>
<intersection>377 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>377,-1652,377,-1646.5</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>-1652 3</intersection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439.5,-1643.5,448.5,-1643.5</points>
<connection>
<GID>808</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>803</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,-1652,430,-1631.5</points>
<intersection>-1652 3</intersection>
<intersection>-1642.5 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430,-1642.5,433.5,-1642.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>429,-1631.5,430,-1631.5</points>
<connection>
<GID>807</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>430,-1652,450.5,-1652</points>
<intersection>430 0</intersection>
<intersection>450.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450.5,-1652,450.5,-1646.5</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<intersection>-1652 3</intersection></vsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523.5,-1645.5,533,-1645.5</points>
<connection>
<GID>812</GID>
<name>OUT</name></connection>
<connection>
<GID>811</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514.5,-1651.5,514.5,-1631.5</points>
<intersection>-1651.5 3</intersection>
<intersection>-1644.5 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514.5,-1644.5,517.5,-1644.5</points>
<connection>
<GID>812</GID>
<name>IN_0</name></connection>
<intersection>514.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513.5,-1631.5,514.5,-1631.5</points>
<connection>
<GID>810</GID>
<name>OUT_0</name></connection>
<intersection>514.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514.5,-1651.5,535,-1651.5</points>
<intersection>514.5 0</intersection>
<intersection>535 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535,-1651.5,535,-1648.5</points>
<connection>
<GID>811</GID>
<name>IN_0</name></connection>
<intersection>-1651.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597.5,-1645.5,606.5,-1645.5</points>
<connection>
<GID>814</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>809</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588,-1651.5,588,-1631.5</points>
<intersection>-1651.5 3</intersection>
<intersection>-1644.5 1</intersection>
<intersection>-1631.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588,-1644.5,591.5,-1644.5</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>588 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587,-1631.5,588,-1631.5</points>
<connection>
<GID>813</GID>
<name>OUT_0</name></connection>
<intersection>588 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>588,-1651.5,608.5,-1651.5</points>
<intersection>588 0</intersection>
<intersection>608.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608.5,-1651.5,608.5,-1648.5</points>
<connection>
<GID>814</GID>
<name>IN_0</name></connection>
<intersection>-1651.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-1634.5,581,-1634.5</points>
<connection>
<GID>815</GID>
<name>OUT</name></connection>
<connection>
<GID>813</GID>
<name>clock</name></connection>
<connection>
<GID>810</GID>
<name>clock</name></connection>
<connection>
<GID>807</GID>
<name>clock</name></connection>
<connection>
<GID>804</GID>
<name>clock</name></connection>
<connection>
<GID>801</GID>
<name>clock</name></connection>
<connection>
<GID>798</GID>
<name>clock</name></connection>
<connection>
<GID>795</GID>
<name>clock</name></connection>
<connection>
<GID>792</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-1709.5,-109.5,-1543.5</points>
<intersection>-1709.5 2</intersection>
<intersection>-1561.5 3</intersection>
<intersection>-1543.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109.5,-1543.5,-8,-1543.5</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1709.5,-109.5,-1709.5</points>
<connection>
<GID>738</GID>
<name>OUT_5</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109.5,-1561.5,-26.5,-1561.5</points>
<connection>
<GID>842</GID>
<name>ENABLE_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-24,-1563.5,588.5,-1563.5</points>
<connection>
<GID>842</GID>
<name>OUT_0</name></connection>
<intersection>33.5 38</intersection>
<intersection>107.5 43</intersection>
<intersection>191.5 42</intersection>
<intersection>265.5 45</intersection>
<intersection>356.5 47</intersection>
<intersection>430.5 49</intersection>
<intersection>514.5 51</intersection>
<intersection>588.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>33.5,-1563.5,33.5,-1551</points>
<connection>
<GID>820</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>191.5,-1563.5,191.5,-1553</points>
<connection>
<GID>826</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>107.5,-1563.5,107.5,-1551</points>
<connection>
<GID>817</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>265.5,-1563.5,265.5,-1553</points>
<connection>
<GID>823</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>356.5,-1563.5,356.5,-1554.5</points>
<connection>
<GID>832</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>430.5,-1563.5,430.5,-1554.5</points>
<connection>
<GID>829</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>514.5,-1563.5,514.5,-1556.5</points>
<connection>
<GID>838</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>588.5,-1563.5,588.5,-1556.5</points>
<connection>
<GID>835</GID>
<name>IN_1</name></connection>
<intersection>-1563.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-1550,49,-1550</points>
<connection>
<GID>820</GID>
<name>OUT</name></connection>
<connection>
<GID>819</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-1558.5,30.5,-1541.5</points>
<intersection>-1558.5 3</intersection>
<intersection>-1549 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-1549,33.5,-1549</points>
<connection>
<GID>820</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-1541.5,30.5,-1541.5</points>
<connection>
<GID>818</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-1558.5,51,-1558.5</points>
<intersection>30.5 0</intersection>
<intersection>51 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51,-1558.5,51,-1553</points>
<connection>
<GID>819</GID>
<name>IN_0</name></connection>
<intersection>-1558.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113.5,-1550,122.5,-1550</points>
<connection>
<GID>822</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>817</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-1560,104,-1541.5</points>
<intersection>-1560 3</intersection>
<intersection>-1549 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-1549,107.5,-1549</points>
<connection>
<GID>817</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-1541.5,104,-1541.5</points>
<connection>
<GID>821</GID>
<name>OUT_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-1560,124.5,-1560</points>
<intersection>104 0</intersection>
<intersection>124.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124.5,-1560,124.5,-1553</points>
<connection>
<GID>822</GID>
<name>IN_0</name></connection>
<intersection>-1560 3</intersection></vsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197.5,-1552,207,-1552</points>
<connection>
<GID>826</GID>
<name>OUT</name></connection>
<connection>
<GID>825</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-1560.5,188.5,-1541.5</points>
<intersection>-1560.5 3</intersection>
<intersection>-1551 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-1551,191.5,-1551</points>
<connection>
<GID>826</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-1541.5,188.5,-1541.5</points>
<connection>
<GID>824</GID>
<name>OUT_0</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188.5,-1560.5,209,-1560.5</points>
<intersection>188.5 0</intersection>
<intersection>209 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209,-1560.5,209,-1555</points>
<connection>
<GID>825</GID>
<name>IN_0</name></connection>
<intersection>-1560.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>271.5,-1552,280.5,-1552</points>
<connection>
<GID>828</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>823</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-1562,262,-1541.5</points>
<connection>
<GID>827</GID>
<name>OUT_0</name></connection>
<intersection>-1562 3</intersection>
<intersection>-1551 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-1551,265.5,-1551</points>
<connection>
<GID>823</GID>
<name>IN_0</name></connection>
<intersection>262 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262,-1562,282.5,-1562</points>
<intersection>262 0</intersection>
<intersection>282.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282.5,-1562,282.5,-1555</points>
<connection>
<GID>828</GID>
<name>IN_0</name></connection>
<intersection>-1562 3</intersection></vsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362.5,-1553.5,372,-1553.5</points>
<connection>
<GID>832</GID>
<name>OUT</name></connection>
<connection>
<GID>831</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353.5,-1562,353.5,-1541.5</points>
<intersection>-1562 3</intersection>
<intersection>-1552.5 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353.5,-1552.5,356.5,-1552.5</points>
<connection>
<GID>832</GID>
<name>IN_0</name></connection>
<intersection>353.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352.5,-1541.5,353.5,-1541.5</points>
<connection>
<GID>830</GID>
<name>OUT_0</name></connection>
<intersection>353.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353.5,-1562,374,-1562</points>
<intersection>353.5 0</intersection>
<intersection>374 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374,-1562,374,-1556.5</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>-1562 3</intersection></vsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>436.5,-1553.5,445.5,-1553.5</points>
<connection>
<GID>834</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>829</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427,-1562,427,-1541.5</points>
<intersection>-1562 3</intersection>
<intersection>-1552.5 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427,-1552.5,430.5,-1552.5</points>
<connection>
<GID>829</GID>
<name>IN_0</name></connection>
<intersection>427 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426,-1541.5,427,-1541.5</points>
<connection>
<GID>833</GID>
<name>OUT_0</name></connection>
<intersection>427 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427,-1562,447.5,-1562</points>
<intersection>427 0</intersection>
<intersection>447.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447.5,-1562,447.5,-1556.5</points>
<connection>
<GID>834</GID>
<name>IN_0</name></connection>
<intersection>-1562 3</intersection></vsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520.5,-1555.5,530,-1555.5</points>
<connection>
<GID>838</GID>
<name>OUT</name></connection>
<connection>
<GID>837</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-1561.5,511.5,-1541.5</points>
<intersection>-1561.5 3</intersection>
<intersection>-1554.5 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511.5,-1554.5,514.5,-1554.5</points>
<connection>
<GID>838</GID>
<name>IN_0</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>510.5,-1541.5,511.5,-1541.5</points>
<connection>
<GID>836</GID>
<name>OUT_0</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511.5,-1561.5,532,-1561.5</points>
<intersection>511.5 0</intersection>
<intersection>532 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532,-1561.5,532,-1558.5</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<intersection>-1561.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>594.5,-1555.5,603.5,-1555.5</points>
<connection>
<GID>840</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>835</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585,-1561.5,585,-1541.5</points>
<intersection>-1561.5 3</intersection>
<intersection>-1554.5 1</intersection>
<intersection>-1541.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585,-1554.5,588.5,-1554.5</points>
<connection>
<GID>835</GID>
<name>IN_0</name></connection>
<intersection>585 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584,-1541.5,585,-1541.5</points>
<connection>
<GID>839</GID>
<name>OUT_0</name></connection>
<intersection>585 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585,-1561.5,605.5,-1561.5</points>
<intersection>585 0</intersection>
<intersection>605.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>605.5,-1561.5,605.5,-1558.5</points>
<connection>
<GID>840</GID>
<name>IN_0</name></connection>
<intersection>-1561.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-1544.5,578,-1544.5</points>
<connection>
<GID>841</GID>
<name>OUT</name></connection>
<connection>
<GID>839</GID>
<name>clock</name></connection>
<connection>
<GID>836</GID>
<name>clock</name></connection>
<connection>
<GID>833</GID>
<name>clock</name></connection>
<connection>
<GID>830</GID>
<name>clock</name></connection>
<connection>
<GID>827</GID>
<name>clock</name></connection>
<connection>
<GID>824</GID>
<name>clock</name></connection>
<connection>
<GID>821</GID>
<name>clock</name></connection>
<connection>
<GID>818</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,-1859.5,-109.5,-1712.5</points>
<intersection>-1859.5 3</intersection>
<intersection>-1841.5 1</intersection>
<intersection>-1712.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109.5,-1841.5,-7,-1841.5</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1712.5,-109.5,-1712.5</points>
<connection>
<GID>738</GID>
<name>OUT_2</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109.5,-1859.5,-25.5,-1859.5</points>
<connection>
<GID>868</GID>
<name>ENABLE_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23,-1861.5,589.5,-1861.5</points>
<connection>
<GID>868</GID>
<name>OUT_0</name></connection>
<intersection>34.5 38</intersection>
<intersection>108.5 43</intersection>
<intersection>192.5 42</intersection>
<intersection>266.5 45</intersection>
<intersection>357.5 47</intersection>
<intersection>431.5 49</intersection>
<intersection>515.5 51</intersection>
<intersection>589.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34.5,-1861.5,34.5,-1849</points>
<connection>
<GID>846</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192.5,-1861.5,192.5,-1851</points>
<connection>
<GID>852</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108.5,-1861.5,108.5,-1849</points>
<connection>
<GID>843</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266.5,-1861.5,266.5,-1851</points>
<connection>
<GID>849</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357.5,-1861.5,357.5,-1852.5</points>
<connection>
<GID>858</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431.5,-1861.5,431.5,-1852.5</points>
<connection>
<GID>855</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515.5,-1861.5,515.5,-1854.5</points>
<connection>
<GID>864</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589.5,-1861.5,589.5,-1854.5</points>
<connection>
<GID>861</GID>
<name>IN_1</name></connection>
<intersection>-1861.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-1848,50,-1848</points>
<connection>
<GID>846</GID>
<name>OUT</name></connection>
<connection>
<GID>845</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-1856.5,31.5,-1839.5</points>
<intersection>-1856.5 3</intersection>
<intersection>-1847 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-1847,34.5,-1847</points>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-1839.5,31.5,-1839.5</points>
<connection>
<GID>844</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-1856.5,52,-1856.5</points>
<intersection>31.5 0</intersection>
<intersection>52 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52,-1856.5,52,-1851</points>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<intersection>-1856.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114.5,-1848,123.5,-1848</points>
<connection>
<GID>848</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>843</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-1858,105,-1839.5</points>
<intersection>-1858 3</intersection>
<intersection>-1847 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-1847,108.5,-1847</points>
<connection>
<GID>843</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-1839.5,105,-1839.5</points>
<connection>
<GID>847</GID>
<name>OUT_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105,-1858,125.5,-1858</points>
<intersection>105 0</intersection>
<intersection>125.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125.5,-1858,125.5,-1851</points>
<connection>
<GID>848</GID>
<name>IN_0</name></connection>
<intersection>-1858 3</intersection></vsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198.5,-1850,208,-1850</points>
<connection>
<GID>852</GID>
<name>OUT</name></connection>
<connection>
<GID>851</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-1858.5,189.5,-1839.5</points>
<intersection>-1858.5 3</intersection>
<intersection>-1849 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,-1849,192.5,-1849</points>
<connection>
<GID>852</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,-1839.5,189.5,-1839.5</points>
<connection>
<GID>850</GID>
<name>OUT_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189.5,-1858.5,210,-1858.5</points>
<intersection>189.5 0</intersection>
<intersection>210 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210,-1858.5,210,-1853</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<intersection>-1858.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272.5,-1850,281.5,-1850</points>
<connection>
<GID>854</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>849</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-1860,263,-1839.5</points>
<connection>
<GID>853</GID>
<name>OUT_0</name></connection>
<intersection>-1860 3</intersection>
<intersection>-1849 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-1849,266.5,-1849</points>
<connection>
<GID>849</GID>
<name>IN_0</name></connection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263,-1860,283.5,-1860</points>
<intersection>263 0</intersection>
<intersection>283.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283.5,-1860,283.5,-1853</points>
<connection>
<GID>854</GID>
<name>IN_0</name></connection>
<intersection>-1860 3</intersection></vsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363.5,-1851.5,373,-1851.5</points>
<connection>
<GID>858</GID>
<name>OUT</name></connection>
<connection>
<GID>857</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-1860,354.5,-1839.5</points>
<intersection>-1860 3</intersection>
<intersection>-1850.5 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354.5,-1850.5,357.5,-1850.5</points>
<connection>
<GID>858</GID>
<name>IN_0</name></connection>
<intersection>354.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353.5,-1839.5,354.5,-1839.5</points>
<connection>
<GID>856</GID>
<name>OUT_0</name></connection>
<intersection>354.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354.5,-1860,375,-1860</points>
<intersection>354.5 0</intersection>
<intersection>375 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375,-1860,375,-1854.5</points>
<connection>
<GID>857</GID>
<name>IN_0</name></connection>
<intersection>-1860 3</intersection></vsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437.5,-1851.5,446.5,-1851.5</points>
<connection>
<GID>860</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>855</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,-1860,428,-1839.5</points>
<intersection>-1860 3</intersection>
<intersection>-1850.5 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428,-1850.5,431.5,-1850.5</points>
<connection>
<GID>855</GID>
<name>IN_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427,-1839.5,428,-1839.5</points>
<connection>
<GID>859</GID>
<name>OUT_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428,-1860,448.5,-1860</points>
<intersection>428 0</intersection>
<intersection>448.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448.5,-1860,448.5,-1854.5</points>
<connection>
<GID>860</GID>
<name>IN_0</name></connection>
<intersection>-1860 3</intersection></vsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521.5,-1853.5,531,-1853.5</points>
<connection>
<GID>864</GID>
<name>OUT</name></connection>
<connection>
<GID>863</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512.5,-1859.5,512.5,-1839.5</points>
<intersection>-1859.5 3</intersection>
<intersection>-1852.5 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512.5,-1852.5,515.5,-1852.5</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<intersection>512.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511.5,-1839.5,512.5,-1839.5</points>
<connection>
<GID>862</GID>
<name>OUT_0</name></connection>
<intersection>512.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512.5,-1859.5,533,-1859.5</points>
<intersection>512.5 0</intersection>
<intersection>533 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533,-1859.5,533,-1856.5</points>
<connection>
<GID>863</GID>
<name>IN_0</name></connection>
<intersection>-1859.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595.5,-1853.5,604.5,-1853.5</points>
<connection>
<GID>866</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>861</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586,-1859.5,586,-1839.5</points>
<intersection>-1859.5 3</intersection>
<intersection>-1852.5 1</intersection>
<intersection>-1839.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586,-1852.5,589.5,-1852.5</points>
<connection>
<GID>861</GID>
<name>IN_0</name></connection>
<intersection>586 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585,-1839.5,586,-1839.5</points>
<connection>
<GID>865</GID>
<name>OUT_0</name></connection>
<intersection>586 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586,-1859.5,606.5,-1859.5</points>
<intersection>586 0</intersection>
<intersection>606.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606.5,-1859.5,606.5,-1856.5</points>
<connection>
<GID>866</GID>
<name>IN_0</name></connection>
<intersection>-1859.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-1842.5,579,-1842.5</points>
<connection>
<GID>867</GID>
<name>OUT</name></connection>
<connection>
<GID>865</GID>
<name>clock</name></connection>
<connection>
<GID>862</GID>
<name>clock</name></connection>
<connection>
<GID>859</GID>
<name>clock</name></connection>
<connection>
<GID>856</GID>
<name>clock</name></connection>
<connection>
<GID>853</GID>
<name>clock</name></connection>
<connection>
<GID>850</GID>
<name>clock</name></connection>
<connection>
<GID>847</GID>
<name>clock</name></connection>
<connection>
<GID>844</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108.5,-1769.5,-108.5,-1711.5</points>
<intersection>-1769.5 3</intersection>
<intersection>-1751.5 1</intersection>
<intersection>-1711.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108.5,-1751.5,-10,-1751.5</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>-108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1711.5,-108.5,-1711.5</points>
<connection>
<GID>738</GID>
<name>OUT_3</name></connection>
<intersection>-108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108.5,-1769.5,-28.5,-1769.5</points>
<connection>
<GID>685</GID>
<name>ENABLE_0</name></connection>
<intersection>-108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-26,-1771.5,586.5,-1771.5</points>
<connection>
<GID>685</GID>
<name>OUT_0</name></connection>
<intersection>31.5 38</intersection>
<intersection>105.5 43</intersection>
<intersection>189.5 42</intersection>
<intersection>263.5 45</intersection>
<intersection>354.5 47</intersection>
<intersection>428.5 49</intersection>
<intersection>512.5 51</intersection>
<intersection>586.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>31.5,-1771.5,31.5,-1759</points>
<connection>
<GID>872</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>189.5,-1771.5,189.5,-1761</points>
<connection>
<GID>669</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>105.5,-1771.5,105.5,-1759</points>
<connection>
<GID>869</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>263.5,-1771.5,263.5,-1761</points>
<connection>
<GID>875</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>354.5,-1771.5,354.5,-1762.5</points>
<connection>
<GID>675</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>428.5,-1771.5,428.5,-1762.5</points>
<connection>
<GID>672</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>512.5,-1771.5,512.5,-1764.5</points>
<connection>
<GID>681</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>586.5,-1771.5,586.5,-1764.5</points>
<connection>
<GID>678</GID>
<name>IN_1</name></connection>
<intersection>-1771.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-1758,47,-1758</points>
<connection>
<GID>872</GID>
<name>OUT</name></connection>
<connection>
<GID>871</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-1766.5,28.5,-1749.5</points>
<intersection>-1766.5 3</intersection>
<intersection>-1757 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-1757,31.5,-1757</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-1749.5,28.5,-1749.5</points>
<connection>
<GID>870</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28.5,-1766.5,49,-1766.5</points>
<intersection>28.5 0</intersection>
<intersection>49 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49,-1766.5,49,-1761</points>
<connection>
<GID>871</GID>
<name>IN_0</name></connection>
<intersection>-1766.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>111.5,-1758,120.5,-1758</points>
<connection>
<GID>874</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>869</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-1768,102,-1749.5</points>
<intersection>-1768 3</intersection>
<intersection>-1757 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-1757,105.5,-1757</points>
<connection>
<GID>869</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-1749.5,102,-1749.5</points>
<connection>
<GID>873</GID>
<name>OUT_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,-1768,122.5,-1768</points>
<intersection>102 0</intersection>
<intersection>122.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122.5,-1768,122.5,-1761</points>
<connection>
<GID>874</GID>
<name>IN_0</name></connection>
<intersection>-1768 3</intersection></vsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195.5,-1760,205,-1760</points>
<connection>
<GID>669</GID>
<name>OUT</name></connection>
<connection>
<GID>877</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-1768.5,186.5,-1749.5</points>
<intersection>-1768.5 3</intersection>
<intersection>-1759 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,-1759,189.5,-1759</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185.5,-1749.5,186.5,-1749.5</points>
<connection>
<GID>876</GID>
<name>OUT_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>186.5,-1768.5,207,-1768.5</points>
<intersection>186.5 0</intersection>
<intersection>207 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207,-1768.5,207,-1763</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<intersection>-1768.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>269.5,-1760,278.5,-1760</points>
<connection>
<GID>671</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>875</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-1770,260,-1749.5</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>-1770 3</intersection>
<intersection>-1759 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-1759,263.5,-1759</points>
<connection>
<GID>875</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260,-1770,280.5,-1770</points>
<intersection>260 0</intersection>
<intersection>280.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>280.5,-1770,280.5,-1763</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>-1770 3</intersection></vsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360.5,-1761.5,370,-1761.5</points>
<connection>
<GID>675</GID>
<name>OUT</name></connection>
<connection>
<GID>674</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,-1770,351.5,-1749.5</points>
<intersection>-1770 3</intersection>
<intersection>-1760.5 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,-1760.5,354.5,-1760.5</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350.5,-1749.5,351.5,-1749.5</points>
<connection>
<GID>673</GID>
<name>OUT_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>351.5,-1770,372,-1770</points>
<intersection>351.5 0</intersection>
<intersection>372 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372,-1770,372,-1764.5</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>-1770 3</intersection></vsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>434.5,-1761.5,443.5,-1761.5</points>
<connection>
<GID>677</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>672</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425,-1770,425,-1749.5</points>
<intersection>-1770 3</intersection>
<intersection>-1760.5 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425,-1760.5,428.5,-1760.5</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>425 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424,-1749.5,425,-1749.5</points>
<connection>
<GID>676</GID>
<name>OUT_0</name></connection>
<intersection>425 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425,-1770,445.5,-1770</points>
<intersection>425 0</intersection>
<intersection>445.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>445.5,-1770,445.5,-1764.5</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>-1770 3</intersection></vsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>518.5,-1763.5,528,-1763.5</points>
<connection>
<GID>681</GID>
<name>OUT</name></connection>
<connection>
<GID>680</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509.5,-1769.5,509.5,-1749.5</points>
<intersection>-1769.5 3</intersection>
<intersection>-1762.5 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,-1762.5,512.5,-1762.5</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>509.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>508.5,-1749.5,509.5,-1749.5</points>
<connection>
<GID>679</GID>
<name>OUT_0</name></connection>
<intersection>509.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>509.5,-1769.5,530,-1769.5</points>
<intersection>509.5 0</intersection>
<intersection>530 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530,-1769.5,530,-1766.5</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>-1769.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>592.5,-1763.5,601.5,-1763.5</points>
<connection>
<GID>683</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>678</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583,-1769.5,583,-1749.5</points>
<intersection>-1769.5 3</intersection>
<intersection>-1762.5 1</intersection>
<intersection>-1749.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583,-1762.5,586.5,-1762.5</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582,-1749.5,583,-1749.5</points>
<connection>
<GID>682</GID>
<name>OUT_0</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583,-1769.5,603.5,-1769.5</points>
<intersection>583 0</intersection>
<intersection>603.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>603.5,-1769.5,603.5,-1766.5</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>-1769.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-1752.5,576,-1752.5</points>
<connection>
<GID>684</GID>
<name>OUT</name></connection>
<connection>
<GID>682</GID>
<name>clock</name></connection>
<connection>
<GID>679</GID>
<name>clock</name></connection>
<connection>
<GID>676</GID>
<name>clock</name></connection>
<connection>
<GID>673</GID>
<name>clock</name></connection>
<connection>
<GID>670</GID>
<name>clock</name></connection>
<connection>
<GID>876</GID>
<name>clock</name></connection>
<connection>
<GID>873</GID>
<name>clock</name></connection>
<connection>
<GID>870</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112.5,-2027.5,-112.5,-1714.5</points>
<intersection>-2027.5 3</intersection>
<intersection>-2009.5 1</intersection>
<intersection>-1714.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112.5,-2009.5,-3,-2009.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1714.5,-112.5,-1714.5</points>
<connection>
<GID>738</GID>
<name>OUT_0</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112.5,-2027.5,-21.5,-2027.5</points>
<connection>
<GID>711</GID>
<name>ENABLE_0</name></connection>
<intersection>-112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-19,-2029.5,593.5,-2029.5</points>
<connection>
<GID>711</GID>
<name>OUT_0</name></connection>
<intersection>38.5 38</intersection>
<intersection>112.5 43</intersection>
<intersection>196.5 42</intersection>
<intersection>270.5 45</intersection>
<intersection>361.5 47</intersection>
<intersection>435.5 49</intersection>
<intersection>519.5 51</intersection>
<intersection>593.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>38.5,-2029.5,38.5,-2017</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>196.5,-2029.5,196.5,-2019</points>
<connection>
<GID>695</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>112.5,-2029.5,112.5,-2017</points>
<connection>
<GID>686</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>270.5,-2029.5,270.5,-2019</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>361.5,-2029.5,361.5,-2020.5</points>
<connection>
<GID>701</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>435.5,-2029.5,435.5,-2020.5</points>
<connection>
<GID>698</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>519.5,-2029.5,519.5,-2022.5</points>
<connection>
<GID>707</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>593.5,-2029.5,593.5,-2022.5</points>
<connection>
<GID>704</GID>
<name>IN_1</name></connection>
<intersection>-2029.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-2016,54,-2016</points>
<connection>
<GID>689</GID>
<name>OUT</name></connection>
<connection>
<GID>688</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-2024.5,35.5,-2007.5</points>
<intersection>-2024.5 3</intersection>
<intersection>-2015 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-2015,38.5,-2015</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-2007.5,35.5,-2007.5</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35.5,-2024.5,56,-2024.5</points>
<intersection>35.5 0</intersection>
<intersection>56 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56,-2024.5,56,-2019</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>-2024.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>118.5,-2016,127.5,-2016</points>
<connection>
<GID>691</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>686</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-2026,109,-2007.5</points>
<intersection>-2026 3</intersection>
<intersection>-2015 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-2015,112.5,-2015</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,-2007.5,109,-2007.5</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>109,-2026,129.5,-2026</points>
<intersection>109 0</intersection>
<intersection>129.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129.5,-2026,129.5,-2019</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>-2026 3</intersection></vsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202.5,-2018,212,-2018</points>
<connection>
<GID>695</GID>
<name>OUT</name></connection>
<connection>
<GID>694</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-2026.5,193.5,-2007.5</points>
<intersection>-2026.5 3</intersection>
<intersection>-2017 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-2017,196.5,-2017</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>192.5,-2007.5,193.5,-2007.5</points>
<connection>
<GID>693</GID>
<name>OUT_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>193.5,-2026.5,214,-2026.5</points>
<intersection>193.5 0</intersection>
<intersection>214 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>214,-2026.5,214,-2021</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>-2026.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>276.5,-2018,285.5,-2018</points>
<connection>
<GID>697</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>692</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267,-2028,267,-2007.5</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>-2028 3</intersection>
<intersection>-2017 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267,-2017,270.5,-2017</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>267,-2028,287.5,-2028</points>
<intersection>267 0</intersection>
<intersection>287.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>287.5,-2028,287.5,-2021</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>-2028 3</intersection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367.5,-2019.5,377,-2019.5</points>
<connection>
<GID>701</GID>
<name>OUT</name></connection>
<connection>
<GID>700</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358.5,-2028,358.5,-2007.5</points>
<intersection>-2028 3</intersection>
<intersection>-2018.5 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358.5,-2018.5,361.5,-2018.5</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>358.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357.5,-2007.5,358.5,-2007.5</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>358.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>358.5,-2028,379,-2028</points>
<intersection>358.5 0</intersection>
<intersection>379 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>379,-2028,379,-2022.5</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-2028 3</intersection></vsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>441.5,-2019.5,450.5,-2019.5</points>
<connection>
<GID>703</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>698</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,-2028,432,-2007.5</points>
<intersection>-2028 3</intersection>
<intersection>-2018.5 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432,-2018.5,435.5,-2018.5</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431,-2007.5,432,-2007.5</points>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432,-2028,452.5,-2028</points>
<intersection>432 0</intersection>
<intersection>452.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>452.5,-2028,452.5,-2022.5</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-2028 3</intersection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>525.5,-2021.5,535,-2021.5</points>
<connection>
<GID>707</GID>
<name>OUT</name></connection>
<connection>
<GID>706</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516.5,-2027.5,516.5,-2007.5</points>
<intersection>-2027.5 3</intersection>
<intersection>-2020.5 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516.5,-2020.5,519.5,-2020.5</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>516.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515.5,-2007.5,516.5,-2007.5</points>
<connection>
<GID>705</GID>
<name>OUT_0</name></connection>
<intersection>516.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>516.5,-2027.5,537,-2027.5</points>
<intersection>516.5 0</intersection>
<intersection>537 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>537,-2027.5,537,-2024.5</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>-2027.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>599.5,-2021.5,608.5,-2021.5</points>
<connection>
<GID>709</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>704</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590,-2027.5,590,-2007.5</points>
<intersection>-2027.5 3</intersection>
<intersection>-2020.5 1</intersection>
<intersection>-2007.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590,-2020.5,593.5,-2020.5</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>590 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589,-2007.5,590,-2007.5</points>
<connection>
<GID>708</GID>
<name>OUT_0</name></connection>
<intersection>590 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>590,-2027.5,610.5,-2027.5</points>
<intersection>590 0</intersection>
<intersection>610.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>610.5,-2027.5,610.5,-2024.5</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>-2027.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-2010.5,583,-2010.5</points>
<connection>
<GID>710</GID>
<name>OUT</name></connection>
<connection>
<GID>708</GID>
<name>clock</name></connection>
<connection>
<GID>705</GID>
<name>clock</name></connection>
<connection>
<GID>702</GID>
<name>clock</name></connection>
<connection>
<GID>699</GID>
<name>clock</name></connection>
<connection>
<GID>696</GID>
<name>clock</name></connection>
<connection>
<GID>693</GID>
<name>clock</name></connection>
<connection>
<GID>690</GID>
<name>clock</name></connection>
<connection>
<GID>687</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110.5,-1937.5,-110.5,-1713.5</points>
<intersection>-1937.5 3</intersection>
<intersection>-1919.5 1</intersection>
<intersection>-1713.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-1919.5,-6,-1919.5</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119,-1713.5,-110.5,-1713.5</points>
<connection>
<GID>738</GID>
<name>OUT_1</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110.5,-1937.5,-24.5,-1937.5</points>
<connection>
<GID>737</GID>
<name>ENABLE_0</name></connection>
<intersection>-110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-22,-1939.5,590.5,-1939.5</points>
<connection>
<GID>737</GID>
<name>OUT_0</name></connection>
<intersection>35.5 38</intersection>
<intersection>109.5 43</intersection>
<intersection>193.5 42</intersection>
<intersection>267.5 45</intersection>
<intersection>358.5 47</intersection>
<intersection>432.5 49</intersection>
<intersection>516.5 51</intersection>
<intersection>590.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>35.5,-1939.5,35.5,-1927</points>
<connection>
<GID>715</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>193.5,-1939.5,193.5,-1929</points>
<connection>
<GID>721</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>109.5,-1939.5,109.5,-1927</points>
<connection>
<GID>712</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>267.5,-1939.5,267.5,-1929</points>
<connection>
<GID>718</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>358.5,-1939.5,358.5,-1930.5</points>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>432.5,-1939.5,432.5,-1930.5</points>
<connection>
<GID>724</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>516.5,-1939.5,516.5,-1932.5</points>
<connection>
<GID>733</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>590.5,-1939.5,590.5,-1932.5</points>
<connection>
<GID>730</GID>
<name>IN_1</name></connection>
<intersection>-1939.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-1926,51,-1926</points>
<connection>
<GID>715</GID>
<name>OUT</name></connection>
<connection>
<GID>714</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-1934.5,32.5,-1917.5</points>
<intersection>-1934.5 3</intersection>
<intersection>-1925 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-1925,35.5,-1925</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-1917.5,32.5,-1917.5</points>
<connection>
<GID>713</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-1934.5,53,-1934.5</points>
<intersection>32.5 0</intersection>
<intersection>53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53,-1934.5,53,-1929</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>-1934.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115.5,-1926,124.5,-1926</points>
<connection>
<GID>717</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>712</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-1936,106,-1917.5</points>
<intersection>-1936 3</intersection>
<intersection>-1925 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-1925,109.5,-1925</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,-1917.5,106,-1917.5</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106,-1936,126.5,-1936</points>
<intersection>106 0</intersection>
<intersection>126.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126.5,-1936,126.5,-1929</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>-1936 3</intersection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199.5,-1928,209,-1928</points>
<connection>
<GID>721</GID>
<name>OUT</name></connection>
<connection>
<GID>720</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-1936.5,190.5,-1917.5</points>
<intersection>-1936.5 3</intersection>
<intersection>-1927 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190.5,-1927,193.5,-1927</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189.5,-1917.5,190.5,-1917.5</points>
<connection>
<GID>719</GID>
<name>OUT_0</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>190.5,-1936.5,211,-1936.5</points>
<intersection>190.5 0</intersection>
<intersection>211 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211,-1936.5,211,-1931</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-1936.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>273.5,-1928,282.5,-1928</points>
<connection>
<GID>723</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>718</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-1938,264,-1917.5</points>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection>
<intersection>-1938 3</intersection>
<intersection>-1927 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264,-1927,267.5,-1927</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>264 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264,-1938,284.5,-1938</points>
<intersection>264 0</intersection>
<intersection>284.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>284.5,-1938,284.5,-1931</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>-1938 3</intersection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364.5,-1929.5,374,-1929.5</points>
<connection>
<GID>727</GID>
<name>OUT</name></connection>
<connection>
<GID>726</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355.5,-1938,355.5,-1917.5</points>
<intersection>-1938 3</intersection>
<intersection>-1928.5 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355.5,-1928.5,358.5,-1928.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>355.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354.5,-1917.5,355.5,-1917.5</points>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection>
<intersection>355.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>355.5,-1938,376,-1938</points>
<intersection>355.5 0</intersection>
<intersection>376 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376,-1938,376,-1932.5</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>-1938 3</intersection></vsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>438.5,-1929.5,447.5,-1929.5</points>
<connection>
<GID>729</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>724</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429,-1938,429,-1917.5</points>
<intersection>-1938 3</intersection>
<intersection>-1928.5 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429,-1928.5,432.5,-1928.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>429 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428,-1917.5,429,-1917.5</points>
<connection>
<GID>728</GID>
<name>OUT_0</name></connection>
<intersection>429 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429,-1938,449.5,-1938</points>
<intersection>429 0</intersection>
<intersection>449.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>449.5,-1938,449.5,-1932.5</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>-1938 3</intersection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522.5,-1931.5,532,-1931.5</points>
<connection>
<GID>733</GID>
<name>OUT</name></connection>
<connection>
<GID>732</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513.5,-1937.5,513.5,-1917.5</points>
<intersection>-1937.5 3</intersection>
<intersection>-1930.5 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-1930.5,516.5,-1930.5</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>513.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>512.5,-1917.5,513.5,-1917.5</points>
<connection>
<GID>731</GID>
<name>OUT_0</name></connection>
<intersection>513.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>513.5,-1937.5,534,-1937.5</points>
<intersection>513.5 0</intersection>
<intersection>534 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534,-1937.5,534,-1934.5</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>-1937.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>596.5,-1931.5,605.5,-1931.5</points>
<connection>
<GID>735</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>730</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587,-1937.5,587,-1917.5</points>
<intersection>-1937.5 3</intersection>
<intersection>-1930.5 1</intersection>
<intersection>-1917.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587,-1930.5,590.5,-1930.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>587 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586,-1917.5,587,-1917.5</points>
<connection>
<GID>734</GID>
<name>OUT_0</name></connection>
<intersection>587 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587,-1937.5,607.5,-1937.5</points>
<intersection>587 0</intersection>
<intersection>607.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>607.5,-1937.5,607.5,-1934.5</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>-1937.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-1920.5,580,-1920.5</points>
<connection>
<GID>736</GID>
<name>OUT</name></connection>
<connection>
<GID>734</GID>
<name>clock</name></connection>
<connection>
<GID>731</GID>
<name>clock</name></connection>
<connection>
<GID>728</GID>
<name>clock</name></connection>
<connection>
<GID>725</GID>
<name>clock</name></connection>
<connection>
<GID>722</GID>
<name>clock</name></connection>
<connection>
<GID>719</GID>
<name>clock</name></connection>
<connection>
<GID>716</GID>
<name>clock</name></connection>
<connection>
<GID>713</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-2580,-111,-2337</points>
<intersection>-2580 2</intersection>
<intersection>-2355 3</intersection>
<intersection>-2337 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-2337,-9.5,-2337</points>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2580,-111,-2580</points>
<connection>
<GID>947</GID>
<name>OUT_6</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111,-2355,-28,-2355</points>
<connection>
<GID>973</GID>
<name>ENABLE_0</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25.5,-2357,587,-2357</points>
<connection>
<GID>973</GID>
<name>OUT_0</name></connection>
<intersection>32 38</intersection>
<intersection>106 43</intersection>
<intersection>190 42</intersection>
<intersection>264 45</intersection>
<intersection>355 47</intersection>
<intersection>429 49</intersection>
<intersection>513 51</intersection>
<intersection>587 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32,-2357,32,-2344.5</points>
<connection>
<GID>951</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190,-2357,190,-2346.5</points>
<connection>
<GID>957</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106,-2357,106,-2344.5</points>
<connection>
<GID>948</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264,-2357,264,-2346.5</points>
<connection>
<GID>954</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355,-2357,355,-2348</points>
<connection>
<GID>963</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429,-2357,429,-2348</points>
<connection>
<GID>960</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513,-2357,513,-2350</points>
<connection>
<GID>969</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587,-2357,587,-2350</points>
<connection>
<GID>966</GID>
<name>IN_1</name></connection>
<intersection>-2357 33</intersection></vsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-2343.5,47.5,-2343.5</points>
<connection>
<GID>951</GID>
<name>OUT</name></connection>
<connection>
<GID>950</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-2352,29,-2335</points>
<intersection>-2352 3</intersection>
<intersection>-2342.5 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-2342.5,32,-2342.5</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-2335,29,-2335</points>
<connection>
<GID>949</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-2352,49.5,-2352</points>
<intersection>29 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-2352,49.5,-2346.5</points>
<connection>
<GID>950</GID>
<name>IN_0</name></connection>
<intersection>-2352 3</intersection></vsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112,-2343.5,121,-2343.5</points>
<connection>
<GID>953</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>948</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-2353.5,102.5,-2335</points>
<intersection>-2353.5 3</intersection>
<intersection>-2342.5 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-2342.5,106,-2342.5</points>
<connection>
<GID>948</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-2335,102.5,-2335</points>
<connection>
<GID>952</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-2353.5,123,-2353.5</points>
<intersection>102.5 0</intersection>
<intersection>123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123,-2353.5,123,-2346.5</points>
<connection>
<GID>953</GID>
<name>IN_0</name></connection>
<intersection>-2353.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,-2345.5,205.5,-2345.5</points>
<connection>
<GID>957</GID>
<name>OUT</name></connection>
<connection>
<GID>956</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-2354,187,-2335</points>
<intersection>-2354 3</intersection>
<intersection>-2344.5 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-2344.5,190,-2344.5</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-2335,187,-2335</points>
<connection>
<GID>955</GID>
<name>OUT_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,-2354,207.5,-2354</points>
<intersection>187 0</intersection>
<intersection>207.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207.5,-2354,207.5,-2348.5</points>
<connection>
<GID>956</GID>
<name>IN_0</name></connection>
<intersection>-2354 3</intersection></vsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270,-2345.5,279,-2345.5</points>
<connection>
<GID>959</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>954</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-2355.5,260.5,-2335</points>
<connection>
<GID>958</GID>
<name>OUT_0</name></connection>
<intersection>-2355.5 3</intersection>
<intersection>-2344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-2344.5,264,-2344.5</points>
<connection>
<GID>954</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-2355.5,281,-2355.5</points>
<intersection>260.5 0</intersection>
<intersection>281 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281,-2355.5,281,-2348.5</points>
<connection>
<GID>959</GID>
<name>IN_0</name></connection>
<intersection>-2355.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-2347,370.5,-2347</points>
<connection>
<GID>963</GID>
<name>OUT</name></connection>
<connection>
<GID>962</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-2355.5,352,-2335</points>
<intersection>-2355.5 3</intersection>
<intersection>-2346 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-2346,355,-2346</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-2335,352,-2335</points>
<connection>
<GID>961</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352,-2355.5,372.5,-2355.5</points>
<intersection>352 0</intersection>
<intersection>372.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372.5,-2355.5,372.5,-2350</points>
<connection>
<GID>962</GID>
<name>IN_0</name></connection>
<intersection>-2355.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435,-2347,444,-2347</points>
<connection>
<GID>965</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>960</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-2355.5,425.5,-2335</points>
<intersection>-2355.5 3</intersection>
<intersection>-2346 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,-2346,429,-2346</points>
<connection>
<GID>960</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,-2335,425.5,-2335</points>
<connection>
<GID>964</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,-2355.5,446,-2355.5</points>
<intersection>425.5 0</intersection>
<intersection>446 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446,-2355.5,446,-2350</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>-2355.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-2349,528.5,-2349</points>
<connection>
<GID>969</GID>
<name>OUT</name></connection>
<connection>
<GID>968</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,-2355,510,-2335</points>
<intersection>-2355 3</intersection>
<intersection>-2348 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,-2348,513,-2348</points>
<connection>
<GID>969</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509,-2335,510,-2335</points>
<connection>
<GID>967</GID>
<name>OUT_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510,-2355,530.5,-2355</points>
<intersection>510 0</intersection>
<intersection>530.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530.5,-2355,530.5,-2352</points>
<connection>
<GID>968</GID>
<name>IN_0</name></connection>
<intersection>-2355 3</intersection></vsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593,-2349,602,-2349</points>
<connection>
<GID>971</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>966</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-2355,583.5,-2335</points>
<intersection>-2355 3</intersection>
<intersection>-2348 1</intersection>
<intersection>-2335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,-2348,587,-2348</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,-2335,583.5,-2335</points>
<connection>
<GID>970</GID>
<name>OUT_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583.5,-2355,604,-2355</points>
<intersection>583.5 0</intersection>
<intersection>604 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604,-2355,604,-2352</points>
<connection>
<GID>971</GID>
<name>IN_0</name></connection>
<intersection>-2355 3</intersection></vsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,-2338,576.5,-2338</points>
<connection>
<GID>972</GID>
<name>OUT</name></connection>
<connection>
<GID>970</GID>
<name>clock</name></connection>
<connection>
<GID>967</GID>
<name>clock</name></connection>
<connection>
<GID>964</GID>
<name>clock</name></connection>
<connection>
<GID>961</GID>
<name>clock</name></connection>
<connection>
<GID>958</GID>
<name>clock</name></connection>
<connection>
<GID>955</GID>
<name>clock</name></connection>
<connection>
<GID>952</GID>
<name>clock</name></connection>
<connection>
<GID>949</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-2579,-112,-2247</points>
<intersection>-2579 2</intersection>
<intersection>-2265 3</intersection>
<intersection>-2247 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112,-2247,-12.5,-2247</points>
<connection>
<GID>998</GID>
<name>IN_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2579,-112,-2579</points>
<connection>
<GID>947</GID>
<name>OUT_7</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112,-2265,-31,-2265</points>
<connection>
<GID>999</GID>
<name>ENABLE_0</name></connection>
<intersection>-112 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-28.5,-2267,584,-2267</points>
<connection>
<GID>999</GID>
<name>OUT_0</name></connection>
<intersection>29 38</intersection>
<intersection>103 43</intersection>
<intersection>187 42</intersection>
<intersection>261 45</intersection>
<intersection>352 47</intersection>
<intersection>426 49</intersection>
<intersection>510 51</intersection>
<intersection>584 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>29,-2267,29,-2254.5</points>
<connection>
<GID>977</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>187,-2267,187,-2256.5</points>
<connection>
<GID>983</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>103,-2267,103,-2254.5</points>
<connection>
<GID>974</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>261,-2267,261,-2256.5</points>
<connection>
<GID>980</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>352,-2267,352,-2258</points>
<connection>
<GID>989</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>426,-2267,426,-2258</points>
<connection>
<GID>986</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>510,-2267,510,-2260</points>
<connection>
<GID>995</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>584,-2267,584,-2260</points>
<connection>
<GID>992</GID>
<name>IN_1</name></connection>
<intersection>-2267 33</intersection></vsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-2253.5,44.5,-2253.5</points>
<connection>
<GID>977</GID>
<name>OUT</name></connection>
<connection>
<GID>976</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-2262,26,-2245</points>
<intersection>-2262 3</intersection>
<intersection>-2252.5 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-2252.5,29,-2252.5</points>
<connection>
<GID>977</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-2245,26,-2245</points>
<connection>
<GID>975</GID>
<name>OUT_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-2262,46.5,-2262</points>
<intersection>26 0</intersection>
<intersection>46.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46.5,-2262,46.5,-2256.5</points>
<connection>
<GID>976</GID>
<name>IN_0</name></connection>
<intersection>-2262 3</intersection></vsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>109,-2253.5,118,-2253.5</points>
<connection>
<GID>979</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>974</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-2263.5,99.5,-2245</points>
<intersection>-2263.5 3</intersection>
<intersection>-2252.5 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-2252.5,103,-2252.5</points>
<connection>
<GID>974</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-2245,99.5,-2245</points>
<connection>
<GID>978</GID>
<name>OUT_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-2263.5,120,-2263.5</points>
<intersection>99.5 0</intersection>
<intersection>120 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>120,-2263.5,120,-2256.5</points>
<connection>
<GID>979</GID>
<name>IN_0</name></connection>
<intersection>-2263.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>193,-2255.5,202.5,-2255.5</points>
<connection>
<GID>983</GID>
<name>OUT</name></connection>
<connection>
<GID>982</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-2264,184,-2245</points>
<intersection>-2264 3</intersection>
<intersection>-2254.5 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-2254.5,187,-2254.5</points>
<connection>
<GID>983</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183,-2245,184,-2245</points>
<connection>
<GID>981</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184,-2264,204.5,-2264</points>
<intersection>184 0</intersection>
<intersection>204.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>204.5,-2264,204.5,-2258.5</points>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<intersection>-2264 3</intersection></vsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>267,-2255.5,276,-2255.5</points>
<connection>
<GID>985</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>980</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-2265.5,257.5,-2245</points>
<connection>
<GID>984</GID>
<name>OUT_0</name></connection>
<intersection>-2265.5 3</intersection>
<intersection>-2254.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-2254.5,261,-2254.5</points>
<connection>
<GID>980</GID>
<name>IN_0</name></connection>
<intersection>257.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,-2265.5,278,-2265.5</points>
<intersection>257.5 0</intersection>
<intersection>278 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>278,-2265.5,278,-2258.5</points>
<connection>
<GID>985</GID>
<name>IN_0</name></connection>
<intersection>-2265.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358,-2257,367.5,-2257</points>
<connection>
<GID>989</GID>
<name>OUT</name></connection>
<connection>
<GID>988</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,-2265.5,349,-2245</points>
<intersection>-2265.5 3</intersection>
<intersection>-2256 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349,-2256,352,-2256</points>
<connection>
<GID>989</GID>
<name>IN_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348,-2245,349,-2245</points>
<connection>
<GID>987</GID>
<name>OUT_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>349,-2265.5,369.5,-2265.5</points>
<intersection>349 0</intersection>
<intersection>369.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>369.5,-2265.5,369.5,-2260</points>
<connection>
<GID>988</GID>
<name>IN_0</name></connection>
<intersection>-2265.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>432,-2257,441,-2257</points>
<connection>
<GID>991</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>986</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422.5,-2265.5,422.5,-2245</points>
<intersection>-2265.5 3</intersection>
<intersection>-2256 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>422.5,-2256,426,-2256</points>
<connection>
<GID>986</GID>
<name>IN_0</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,-2245,422.5,-2245</points>
<connection>
<GID>990</GID>
<name>OUT_0</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>422.5,-2265.5,443,-2265.5</points>
<intersection>422.5 0</intersection>
<intersection>443 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>443,-2265.5,443,-2260</points>
<connection>
<GID>991</GID>
<name>IN_0</name></connection>
<intersection>-2265.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>516,-2259,525.5,-2259</points>
<connection>
<GID>995</GID>
<name>OUT</name></connection>
<connection>
<GID>994</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,-2265,507,-2245</points>
<intersection>-2265 3</intersection>
<intersection>-2258 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507,-2258,510,-2258</points>
<connection>
<GID>995</GID>
<name>IN_0</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>506,-2245,507,-2245</points>
<connection>
<GID>993</GID>
<name>OUT_0</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>507,-2265,527.5,-2265</points>
<intersection>507 0</intersection>
<intersection>527.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>527.5,-2265,527.5,-2262</points>
<connection>
<GID>994</GID>
<name>IN_0</name></connection>
<intersection>-2265 3</intersection></vsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>590,-2259,599,-2259</points>
<connection>
<GID>997</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>992</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>580.5,-2265,580.5,-2245</points>
<intersection>-2265 3</intersection>
<intersection>-2258 1</intersection>
<intersection>-2245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>580.5,-2258,584,-2258</points>
<connection>
<GID>992</GID>
<name>IN_0</name></connection>
<intersection>580.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>579.5,-2245,580.5,-2245</points>
<connection>
<GID>996</GID>
<name>OUT_0</name></connection>
<intersection>580.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>580.5,-2265,601,-2265</points>
<intersection>580.5 0</intersection>
<intersection>601 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>601,-2265,601,-2262</points>
<connection>
<GID>997</GID>
<name>IN_0</name></connection>
<intersection>-2265 3</intersection></vsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-2248,573.5,-2248</points>
<connection>
<GID>998</GID>
<name>OUT</name></connection>
<connection>
<GID>996</GID>
<name>clock</name></connection>
<connection>
<GID>993</GID>
<name>clock</name></connection>
<connection>
<GID>990</GID>
<name>clock</name></connection>
<connection>
<GID>987</GID>
<name>clock</name></connection>
<connection>
<GID>984</GID>
<name>clock</name></connection>
<connection>
<GID>981</GID>
<name>clock</name></connection>
<connection>
<GID>978</GID>
<name>clock</name></connection>
<connection>
<GID>975</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-2582,-109,-2505</points>
<intersection>-2582 2</intersection>
<intersection>-2523 3</intersection>
<intersection>-2505 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-2505,-5.5,-2505</points>
<connection>
<GID>1024</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2582,-109,-2582</points>
<connection>
<GID>947</GID>
<name>OUT_4</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-2523,-24,-2523</points>
<connection>
<GID>1025</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21.5,-2525,591,-2525</points>
<connection>
<GID>1025</GID>
<name>OUT_0</name></connection>
<intersection>36 38</intersection>
<intersection>110 43</intersection>
<intersection>194 42</intersection>
<intersection>268 45</intersection>
<intersection>359 47</intersection>
<intersection>433 49</intersection>
<intersection>517 51</intersection>
<intersection>591 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36,-2525,36,-2512.5</points>
<connection>
<GID>1003</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194,-2525,194,-2514.5</points>
<connection>
<GID>1009</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110,-2525,110,-2512.5</points>
<connection>
<GID>1000</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268,-2525,268,-2514.5</points>
<connection>
<GID>1006</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359,-2525,359,-2516</points>
<connection>
<GID>1015</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433,-2525,433,-2516</points>
<connection>
<GID>1012</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517,-2525,517,-2518</points>
<connection>
<GID>1021</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591,-2525,591,-2518</points>
<connection>
<GID>1018</GID>
<name>IN_1</name></connection>
<intersection>-2525 33</intersection></vsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-2511.5,51.5,-2511.5</points>
<connection>
<GID>1003</GID>
<name>OUT</name></connection>
<connection>
<GID>1002</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-2520,33,-2503</points>
<intersection>-2520 3</intersection>
<intersection>-2510.5 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-2510.5,36,-2510.5</points>
<connection>
<GID>1003</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-2503,33,-2503</points>
<connection>
<GID>1001</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-2520,53.5,-2520</points>
<intersection>33 0</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-2520,53.5,-2514.5</points>
<connection>
<GID>1002</GID>
<name>IN_0</name></connection>
<intersection>-2520 3</intersection></vsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116,-2511.5,125,-2511.5</points>
<connection>
<GID>1005</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1000</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-2521.5,106.5,-2503</points>
<intersection>-2521.5 3</intersection>
<intersection>-2510.5 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-2510.5,110,-2510.5</points>
<connection>
<GID>1000</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-2503,106.5,-2503</points>
<connection>
<GID>1004</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,-2521.5,127,-2521.5</points>
<intersection>106.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-2521.5,127,-2514.5</points>
<connection>
<GID>1005</GID>
<name>IN_0</name></connection>
<intersection>-2521.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-2513.5,209.5,-2513.5</points>
<connection>
<GID>1009</GID>
<name>OUT</name></connection>
<connection>
<GID>1008</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-2522,191,-2503</points>
<intersection>-2522 3</intersection>
<intersection>-2512.5 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-2512.5,194,-2512.5</points>
<connection>
<GID>1009</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,-2503,191,-2503</points>
<connection>
<GID>1007</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191,-2522,211.5,-2522</points>
<intersection>191 0</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211.5,-2522,211.5,-2516.5</points>
<connection>
<GID>1008</GID>
<name>IN_0</name></connection>
<intersection>-2522 3</intersection></vsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274,-2513.5,283,-2513.5</points>
<connection>
<GID>1011</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1006</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-2523.5,264.5,-2503</points>
<connection>
<GID>1010</GID>
<name>OUT_0</name></connection>
<intersection>-2523.5 3</intersection>
<intersection>-2512.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-2512.5,268,-2512.5</points>
<connection>
<GID>1006</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264.5,-2523.5,285,-2523.5</points>
<intersection>264.5 0</intersection>
<intersection>285 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285,-2523.5,285,-2516.5</points>
<connection>
<GID>1011</GID>
<name>IN_0</name></connection>
<intersection>-2523.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365,-2515,374.5,-2515</points>
<connection>
<GID>1015</GID>
<name>OUT</name></connection>
<connection>
<GID>1014</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-2523.5,356,-2503</points>
<intersection>-2523.5 3</intersection>
<intersection>-2514 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-2514,359,-2514</points>
<connection>
<GID>1015</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355,-2503,356,-2503</points>
<connection>
<GID>1013</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356,-2523.5,376.5,-2523.5</points>
<intersection>356 0</intersection>
<intersection>376.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376.5,-2523.5,376.5,-2518</points>
<connection>
<GID>1014</GID>
<name>IN_0</name></connection>
<intersection>-2523.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439,-2515,448,-2515</points>
<connection>
<GID>1017</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1012</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-2523.5,429.5,-2503</points>
<intersection>-2523.5 3</intersection>
<intersection>-2514 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,-2514,433,-2514</points>
<connection>
<GID>1012</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,-2503,429.5,-2503</points>
<connection>
<GID>1016</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,-2523.5,450,-2523.5</points>
<intersection>429.5 0</intersection>
<intersection>450 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450,-2523.5,450,-2518</points>
<connection>
<GID>1017</GID>
<name>IN_0</name></connection>
<intersection>-2523.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523,-2517,532.5,-2517</points>
<connection>
<GID>1021</GID>
<name>OUT</name></connection>
<connection>
<GID>1020</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-2523,514,-2503</points>
<intersection>-2523 3</intersection>
<intersection>-2516 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-2516,517,-2516</points>
<connection>
<GID>1021</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,-2503,514,-2503</points>
<connection>
<GID>1019</GID>
<name>OUT_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514,-2523,534.5,-2523</points>
<intersection>514 0</intersection>
<intersection>534.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534.5,-2523,534.5,-2520</points>
<connection>
<GID>1020</GID>
<name>IN_0</name></connection>
<intersection>-2523 3</intersection></vsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597,-2517,606,-2517</points>
<connection>
<GID>1023</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1018</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,-2523,587.5,-2503</points>
<intersection>-2523 3</intersection>
<intersection>-2516 1</intersection>
<intersection>-2503 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,-2516,591,-2516</points>
<connection>
<GID>1018</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586.5,-2503,587.5,-2503</points>
<connection>
<GID>1022</GID>
<name>OUT_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587.5,-2523,608,-2523</points>
<intersection>587.5 0</intersection>
<intersection>608 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608,-2523,608,-2520</points>
<connection>
<GID>1023</GID>
<name>IN_0</name></connection>
<intersection>-2523 3</intersection></vsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-2506,580.5,-2506</points>
<connection>
<GID>1004</GID>
<name>clock</name></connection>
<connection>
<GID>1024</GID>
<name>OUT</name></connection>
<connection>
<GID>1022</GID>
<name>clock</name></connection>
<connection>
<GID>1019</GID>
<name>clock</name></connection>
<connection>
<GID>1016</GID>
<name>clock</name></connection>
<connection>
<GID>1010</GID>
<name>clock</name></connection>
<connection>
<GID>1007</GID>
<name>clock</name></connection>
<connection>
<GID>1001</GID>
<name>clock</name></connection>
<connection>
<GID>1013</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-2581,-110,-2415</points>
<intersection>-2581 2</intersection>
<intersection>-2433 3</intersection>
<intersection>-2415 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-2415,-8.5,-2415</points>
<connection>
<GID>1050</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2581,-110,-2581</points>
<connection>
<GID>947</GID>
<name>OUT_5</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-2433,-27,-2433</points>
<connection>
<GID>1051</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-24.5,-2435,588,-2435</points>
<connection>
<GID>1051</GID>
<name>OUT_0</name></connection>
<intersection>33 38</intersection>
<intersection>107 43</intersection>
<intersection>191 42</intersection>
<intersection>265 45</intersection>
<intersection>356 47</intersection>
<intersection>430 49</intersection>
<intersection>514 51</intersection>
<intersection>588 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>33,-2435,33,-2422.5</points>
<connection>
<GID>1029</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>191,-2435,191,-2424.5</points>
<connection>
<GID>1035</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>107,-2435,107,-2422.5</points>
<connection>
<GID>1026</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>265,-2435,265,-2424.5</points>
<connection>
<GID>1032</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>356,-2435,356,-2426</points>
<connection>
<GID>1041</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>430,-2435,430,-2426</points>
<connection>
<GID>1038</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>514,-2435,514,-2428</points>
<connection>
<GID>1047</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>588,-2435,588,-2428</points>
<connection>
<GID>1044</GID>
<name>IN_1</name></connection>
<intersection>-2435 33</intersection></vsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-2421.5,48.5,-2421.5</points>
<connection>
<GID>1029</GID>
<name>OUT</name></connection>
<connection>
<GID>1028</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-2430,30,-2413</points>
<intersection>-2430 3</intersection>
<intersection>-2420.5 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-2420.5,33,-2420.5</points>
<connection>
<GID>1029</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-2413,30,-2413</points>
<connection>
<GID>1027</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30,-2430,50.5,-2430</points>
<intersection>30 0</intersection>
<intersection>50.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50.5,-2430,50.5,-2424.5</points>
<connection>
<GID>1028</GID>
<name>IN_0</name></connection>
<intersection>-2430 3</intersection></vsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113,-2421.5,122,-2421.5</points>
<connection>
<GID>1031</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1026</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-2431.5,103.5,-2413</points>
<intersection>-2431.5 3</intersection>
<intersection>-2420.5 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-2420.5,107,-2420.5</points>
<connection>
<GID>1026</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-2413,103.5,-2413</points>
<connection>
<GID>1030</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,-2431.5,124,-2431.5</points>
<intersection>103.5 0</intersection>
<intersection>124 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124,-2431.5,124,-2424.5</points>
<connection>
<GID>1031</GID>
<name>IN_0</name></connection>
<intersection>-2431.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-2423.5,206.5,-2423.5</points>
<connection>
<GID>1035</GID>
<name>OUT</name></connection>
<connection>
<GID>1034</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-2432,188,-2413</points>
<intersection>-2432 3</intersection>
<intersection>-2422.5 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188,-2422.5,191,-2422.5</points>
<connection>
<GID>1035</GID>
<name>IN_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-2413,188,-2413</points>
<connection>
<GID>1033</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188,-2432,208.5,-2432</points>
<intersection>188 0</intersection>
<intersection>208.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208.5,-2432,208.5,-2426.5</points>
<connection>
<GID>1034</GID>
<name>IN_0</name></connection>
<intersection>-2432 3</intersection></vsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>271,-2423.5,280,-2423.5</points>
<connection>
<GID>1037</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1032</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-2433.5,261.5,-2413</points>
<connection>
<GID>1036</GID>
<name>OUT_0</name></connection>
<intersection>-2433.5 3</intersection>
<intersection>-2422.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-2422.5,265,-2422.5</points>
<connection>
<GID>1032</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-2433.5,282,-2433.5</points>
<intersection>261.5 0</intersection>
<intersection>282 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282,-2433.5,282,-2426.5</points>
<connection>
<GID>1037</GID>
<name>IN_0</name></connection>
<intersection>-2433.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362,-2425,371.5,-2425</points>
<connection>
<GID>1041</GID>
<name>OUT</name></connection>
<connection>
<GID>1040</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-2433.5,353,-2413</points>
<intersection>-2433.5 3</intersection>
<intersection>-2424 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-2424,356,-2424</points>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-2413,353,-2413</points>
<connection>
<GID>1039</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353,-2433.5,373.5,-2433.5</points>
<intersection>353 0</intersection>
<intersection>373.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>373.5,-2433.5,373.5,-2428</points>
<connection>
<GID>1040</GID>
<name>IN_0</name></connection>
<intersection>-2433.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>436,-2425,445,-2425</points>
<connection>
<GID>1043</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1038</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-2433.5,426.5,-2413</points>
<intersection>-2433.5 3</intersection>
<intersection>-2424 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426.5,-2424,430,-2424</points>
<connection>
<GID>1038</GID>
<name>IN_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425.5,-2413,426.5,-2413</points>
<connection>
<GID>1042</GID>
<name>OUT_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426.5,-2433.5,447,-2433.5</points>
<intersection>426.5 0</intersection>
<intersection>447 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447,-2433.5,447,-2428</points>
<connection>
<GID>1043</GID>
<name>IN_0</name></connection>
<intersection>-2433.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520,-2427,529.5,-2427</points>
<connection>
<GID>1047</GID>
<name>OUT</name></connection>
<connection>
<GID>1046</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,-2433,511,-2413</points>
<intersection>-2433 3</intersection>
<intersection>-2426 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,-2426,514,-2426</points>
<connection>
<GID>1047</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>510,-2413,511,-2413</points>
<connection>
<GID>1045</GID>
<name>OUT_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511,-2433,531.5,-2433</points>
<intersection>511 0</intersection>
<intersection>531.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531.5,-2433,531.5,-2430</points>
<connection>
<GID>1046</GID>
<name>IN_0</name></connection>
<intersection>-2433 3</intersection></vsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>594,-2427,603,-2427</points>
<connection>
<GID>1049</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1044</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,-2433,584.5,-2413</points>
<intersection>-2433 3</intersection>
<intersection>-2426 1</intersection>
<intersection>-2413 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584.5,-2426,588,-2426</points>
<connection>
<GID>1044</GID>
<name>IN_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583.5,-2413,584.5,-2413</points>
<connection>
<GID>1048</GID>
<name>OUT_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>584.5,-2433,605,-2433</points>
<intersection>584.5 0</intersection>
<intersection>605 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>605,-2433,605,-2430</points>
<connection>
<GID>1049</GID>
<name>IN_0</name></connection>
<intersection>-2433 3</intersection></vsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-2416,577.5,-2416</points>
<connection>
<GID>1050</GID>
<name>OUT</name></connection>
<connection>
<GID>1048</GID>
<name>clock</name></connection>
<connection>
<GID>1045</GID>
<name>clock</name></connection>
<connection>
<GID>1042</GID>
<name>clock</name></connection>
<connection>
<GID>1039</GID>
<name>clock</name></connection>
<connection>
<GID>1036</GID>
<name>clock</name></connection>
<connection>
<GID>1033</GID>
<name>clock</name></connection>
<connection>
<GID>1030</GID>
<name>clock</name></connection>
<connection>
<GID>1027</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-2731,-110,-2584</points>
<intersection>-2731 3</intersection>
<intersection>-2713 1</intersection>
<intersection>-2584 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-2713,-7.5,-2713</points>
<connection>
<GID>1076</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2584,-110,-2584</points>
<connection>
<GID>947</GID>
<name>OUT_2</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-2731,-26,-2731</points>
<connection>
<GID>1077</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-2733,589,-2733</points>
<connection>
<GID>1077</GID>
<name>OUT_0</name></connection>
<intersection>34 38</intersection>
<intersection>108 43</intersection>
<intersection>192 42</intersection>
<intersection>266 45</intersection>
<intersection>357 47</intersection>
<intersection>431 49</intersection>
<intersection>515 51</intersection>
<intersection>589 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34,-2733,34,-2720.5</points>
<connection>
<GID>1055</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192,-2733,192,-2722.5</points>
<connection>
<GID>1061</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108,-2733,108,-2720.5</points>
<connection>
<GID>1052</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266,-2733,266,-2722.5</points>
<connection>
<GID>1058</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357,-2733,357,-2724</points>
<connection>
<GID>1067</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431,-2733,431,-2724</points>
<connection>
<GID>1064</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515,-2733,515,-2726</points>
<connection>
<GID>1073</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589,-2733,589,-2726</points>
<connection>
<GID>1070</GID>
<name>IN_1</name></connection>
<intersection>-2733 33</intersection></vsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-2719.5,49.5,-2719.5</points>
<connection>
<GID>1055</GID>
<name>OUT</name></connection>
<connection>
<GID>1054</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-2728,31,-2711</points>
<intersection>-2728 3</intersection>
<intersection>-2718.5 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-2718.5,34,-2718.5</points>
<connection>
<GID>1055</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-2711,31,-2711</points>
<connection>
<GID>1053</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-2728,51.5,-2728</points>
<intersection>31 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-2728,51.5,-2722.5</points>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection>
<intersection>-2728 3</intersection></vsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114,-2719.5,123,-2719.5</points>
<connection>
<GID>1057</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1052</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-2729.5,104.5,-2711</points>
<intersection>-2729.5 3</intersection>
<intersection>-2718.5 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-2718.5,108,-2718.5</points>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-2711,104.5,-2711</points>
<connection>
<GID>1056</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-2729.5,125,-2729.5</points>
<intersection>104.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-2729.5,125,-2722.5</points>
<connection>
<GID>1057</GID>
<name>IN_0</name></connection>
<intersection>-2729.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-2721.5,207.5,-2721.5</points>
<connection>
<GID>1061</GID>
<name>OUT</name></connection>
<connection>
<GID>1060</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-2730,189,-2711</points>
<intersection>-2730 3</intersection>
<intersection>-2720.5 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-2720.5,192,-2720.5</points>
<connection>
<GID>1061</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188,-2711,189,-2711</points>
<connection>
<GID>1059</GID>
<name>OUT_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189,-2730,209.5,-2730</points>
<intersection>189 0</intersection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,-2730,209.5,-2724.5</points>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection>
<intersection>-2730 3</intersection></vsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272,-2721.5,281,-2721.5</points>
<connection>
<GID>1063</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1058</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-2731.5,262.5,-2711</points>
<connection>
<GID>1062</GID>
<name>OUT_0</name></connection>
<intersection>-2731.5 3</intersection>
<intersection>-2720.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-2720.5,266,-2720.5</points>
<connection>
<GID>1058</GID>
<name>IN_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262.5,-2731.5,283,-2731.5</points>
<intersection>262.5 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-2731.5,283,-2724.5</points>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection>
<intersection>-2731.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363,-2723,372.5,-2723</points>
<connection>
<GID>1067</GID>
<name>OUT</name></connection>
<connection>
<GID>1066</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-2731.5,354,-2711</points>
<intersection>-2731.5 3</intersection>
<intersection>-2722 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-2722,357,-2722</points>
<connection>
<GID>1067</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-2711,354,-2711</points>
<connection>
<GID>1065</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354,-2731.5,374.5,-2731.5</points>
<intersection>354 0</intersection>
<intersection>374.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374.5,-2731.5,374.5,-2726</points>
<connection>
<GID>1066</GID>
<name>IN_0</name></connection>
<intersection>-2731.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437,-2723,446,-2723</points>
<connection>
<GID>1069</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1064</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-2731.5,427.5,-2711</points>
<intersection>-2731.5 3</intersection>
<intersection>-2722 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-2722,431,-2722</points>
<connection>
<GID>1064</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426.5,-2711,427.5,-2711</points>
<connection>
<GID>1068</GID>
<name>OUT_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-2731.5,448,-2731.5</points>
<intersection>427.5 0</intersection>
<intersection>448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448,-2731.5,448,-2726</points>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection>
<intersection>-2731.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521,-2725,530.5,-2725</points>
<connection>
<GID>1073</GID>
<name>OUT</name></connection>
<connection>
<GID>1072</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,-2731,512,-2711</points>
<intersection>-2731 3</intersection>
<intersection>-2724 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-2724,515,-2724</points>
<connection>
<GID>1073</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,-2711,512,-2711</points>
<connection>
<GID>1071</GID>
<name>OUT_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512,-2731,532.5,-2731</points>
<intersection>512 0</intersection>
<intersection>532.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532.5,-2731,532.5,-2728</points>
<connection>
<GID>1072</GID>
<name>IN_0</name></connection>
<intersection>-2731 3</intersection></vsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595,-2725,604,-2725</points>
<connection>
<GID>1075</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1070</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-2731,585.5,-2711</points>
<intersection>-2731 3</intersection>
<intersection>-2724 1</intersection>
<intersection>-2711 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-2724,589,-2724</points>
<connection>
<GID>1070</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,-2711,585.5,-2711</points>
<connection>
<GID>1074</GID>
<name>OUT_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-2731,606,-2731</points>
<intersection>585.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-2731,606,-2728</points>
<connection>
<GID>1075</GID>
<name>IN_0</name></connection>
<intersection>-2731 3</intersection></vsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-2714,578.5,-2714</points>
<connection>
<GID>1076</GID>
<name>OUT</name></connection>
<connection>
<GID>1074</GID>
<name>clock</name></connection>
<connection>
<GID>1071</GID>
<name>clock</name></connection>
<connection>
<GID>1068</GID>
<name>clock</name></connection>
<connection>
<GID>1065</GID>
<name>clock</name></connection>
<connection>
<GID>1062</GID>
<name>clock</name></connection>
<connection>
<GID>1059</GID>
<name>clock</name></connection>
<connection>
<GID>1056</GID>
<name>clock</name></connection>
<connection>
<GID>1053</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-2641,-109,-2583</points>
<intersection>-2641 3</intersection>
<intersection>-2623 1</intersection>
<intersection>-2583 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-2623,-10.5,-2623</points>
<connection>
<GID>893</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2583,-109,-2583</points>
<connection>
<GID>947</GID>
<name>OUT_3</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-2641,-29,-2641</points>
<connection>
<GID>894</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-26.5,-2643,586,-2643</points>
<connection>
<GID>894</GID>
<name>OUT_0</name></connection>
<intersection>31 38</intersection>
<intersection>105 43</intersection>
<intersection>189 42</intersection>
<intersection>263 45</intersection>
<intersection>354 47</intersection>
<intersection>428 49</intersection>
<intersection>512 51</intersection>
<intersection>586 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>31,-2643,31,-2630.5</points>
<connection>
<GID>1081</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>189,-2643,189,-2632.5</points>
<connection>
<GID>878</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>105,-2643,105,-2630.5</points>
<connection>
<GID>1078</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>263,-2643,263,-2632.5</points>
<connection>
<GID>1084</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>354,-2643,354,-2634</points>
<connection>
<GID>884</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>428,-2643,428,-2634</points>
<connection>
<GID>881</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>512,-2643,512,-2636</points>
<connection>
<GID>890</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>586,-2643,586,-2636</points>
<connection>
<GID>887</GID>
<name>IN_1</name></connection>
<intersection>-2643 33</intersection></vsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-2638,28,-2621</points>
<intersection>-2638 3</intersection>
<intersection>-2628.5 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-2628.5,31,-2628.5</points>
<connection>
<GID>1081</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-2621,28,-2621</points>
<connection>
<GID>1079</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-2638,48.5,-2638</points>
<intersection>28 0</intersection>
<intersection>48.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-2638,48.5,-2632.5</points>
<connection>
<GID>1080</GID>
<name>IN_0</name></connection>
<intersection>-2638 3</intersection></vsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>111,-2629.5,120,-2629.5</points>
<connection>
<GID>1083</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1078</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-2639.5,101.5,-2621</points>
<intersection>-2639.5 3</intersection>
<intersection>-2628.5 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-2628.5,105,-2628.5</points>
<connection>
<GID>1078</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-2621,101.5,-2621</points>
<connection>
<GID>1082</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101.5,-2639.5,122,-2639.5</points>
<intersection>101.5 0</intersection>
<intersection>122 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122,-2639.5,122,-2632.5</points>
<connection>
<GID>1083</GID>
<name>IN_0</name></connection>
<intersection>-2639.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-2631.5,204.5,-2631.5</points>
<connection>
<GID>1086</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>878</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-2640,186,-2621</points>
<intersection>-2640 3</intersection>
<intersection>-2630.5 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186,-2630.5,189,-2630.5</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-2621,186,-2621</points>
<connection>
<GID>1085</GID>
<name>OUT_0</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>186,-2640,206.5,-2640</points>
<intersection>186 0</intersection>
<intersection>206.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>206.5,-2640,206.5,-2634.5</points>
<connection>
<GID>1086</GID>
<name>IN_0</name></connection>
<intersection>-2640 3</intersection></vsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>269,-2631.5,278,-2631.5</points>
<connection>
<GID>1084</GID>
<name>OUT</name></connection>
<connection>
<GID>880</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-2641.5,259.5,-2621</points>
<connection>
<GID>879</GID>
<name>OUT_0</name></connection>
<intersection>-2641.5 3</intersection>
<intersection>-2630.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-2630.5,263,-2630.5</points>
<connection>
<GID>1084</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259.5,-2641.5,280,-2641.5</points>
<intersection>259.5 0</intersection>
<intersection>280 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>280,-2641.5,280,-2634.5</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<intersection>-2641.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360,-2633,369.5,-2633</points>
<connection>
<GID>884</GID>
<name>OUT</name></connection>
<connection>
<GID>883</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-2641.5,351,-2621</points>
<intersection>-2641.5 3</intersection>
<intersection>-2632 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,-2632,354,-2632</points>
<connection>
<GID>884</GID>
<name>IN_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-2621,351,-2621</points>
<connection>
<GID>882</GID>
<name>OUT_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>351,-2641.5,371.5,-2641.5</points>
<intersection>351 0</intersection>
<intersection>371.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>371.5,-2641.5,371.5,-2636</points>
<connection>
<GID>883</GID>
<name>IN_0</name></connection>
<intersection>-2641.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>434,-2633,443,-2633</points>
<connection>
<GID>886</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>881</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,-2641.5,424.5,-2621</points>
<intersection>-2641.5 3</intersection>
<intersection>-2632 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424.5,-2632,428,-2632</points>
<connection>
<GID>881</GID>
<name>IN_0</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423.5,-2621,424.5,-2621</points>
<connection>
<GID>885</GID>
<name>OUT_0</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>424.5,-2641.5,445,-2641.5</points>
<intersection>424.5 0</intersection>
<intersection>445 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>445,-2641.5,445,-2636</points>
<connection>
<GID>886</GID>
<name>IN_0</name></connection>
<intersection>-2641.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>518,-2635,527.5,-2635</points>
<connection>
<GID>890</GID>
<name>OUT</name></connection>
<connection>
<GID>889</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,-2641,509,-2621</points>
<intersection>-2641 3</intersection>
<intersection>-2634 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509,-2634,512,-2634</points>
<connection>
<GID>890</GID>
<name>IN_0</name></connection>
<intersection>509 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>508,-2621,509,-2621</points>
<connection>
<GID>888</GID>
<name>OUT_0</name></connection>
<intersection>509 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>509,-2641,529.5,-2641</points>
<intersection>509 0</intersection>
<intersection>529.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>529.5,-2641,529.5,-2638</points>
<connection>
<GID>889</GID>
<name>IN_0</name></connection>
<intersection>-2641 3</intersection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>592,-2635,601,-2635</points>
<connection>
<GID>892</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>887</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>582.5,-2641,582.5,-2621</points>
<intersection>-2641 3</intersection>
<intersection>-2634 1</intersection>
<intersection>-2621 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>582.5,-2634,586,-2634</points>
<connection>
<GID>887</GID>
<name>IN_0</name></connection>
<intersection>582.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>581.5,-2621,582.5,-2621</points>
<connection>
<GID>891</GID>
<name>OUT_0</name></connection>
<intersection>582.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>582.5,-2641,603,-2641</points>
<intersection>582.5 0</intersection>
<intersection>603 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>603,-2641,603,-2638</points>
<connection>
<GID>892</GID>
<name>IN_0</name></connection>
<intersection>-2641 3</intersection></vsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,-2624,575.5,-2624</points>
<connection>
<GID>1085</GID>
<name>clock</name></connection>
<connection>
<GID>1082</GID>
<name>clock</name></connection>
<connection>
<GID>1079</GID>
<name>clock</name></connection>
<connection>
<GID>893</GID>
<name>OUT</name></connection>
<connection>
<GID>891</GID>
<name>clock</name></connection>
<connection>
<GID>888</GID>
<name>clock</name></connection>
<connection>
<GID>885</GID>
<name>clock</name></connection>
<connection>
<GID>882</GID>
<name>clock</name></connection>
<connection>
<GID>879</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113,-2899,-113,-2586</points>
<intersection>-2899 3</intersection>
<intersection>-2881 1</intersection>
<intersection>-2586 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-113,-2881,-3.5,-2881</points>
<connection>
<GID>919</GID>
<name>IN_0</name></connection>
<intersection>-113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2586,-113,-2586</points>
<connection>
<GID>947</GID>
<name>OUT_0</name></connection>
<intersection>-113 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-113,-2899,-22,-2899</points>
<connection>
<GID>920</GID>
<name>ENABLE_0</name></connection>
<intersection>-113 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-19.5,-2901,593,-2901</points>
<connection>
<GID>920</GID>
<name>OUT_0</name></connection>
<intersection>38 38</intersection>
<intersection>112 43</intersection>
<intersection>196 42</intersection>
<intersection>270 45</intersection>
<intersection>361 47</intersection>
<intersection>435 49</intersection>
<intersection>519 51</intersection>
<intersection>593 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>38,-2901,38,-2888.5</points>
<connection>
<GID>898</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>196,-2901,196,-2890.5</points>
<connection>
<GID>904</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>112,-2901,112,-2888.5</points>
<connection>
<GID>895</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>270,-2901,270,-2890.5</points>
<connection>
<GID>901</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>361,-2901,361,-2892</points>
<connection>
<GID>910</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>435,-2901,435,-2892</points>
<connection>
<GID>907</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>519,-2901,519,-2894</points>
<connection>
<GID>916</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>593,-2901,593,-2894</points>
<connection>
<GID>913</GID>
<name>IN_1</name></connection>
<intersection>-2901 33</intersection></vsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-2887.5,53.5,-2887.5</points>
<connection>
<GID>898</GID>
<name>OUT</name></connection>
<connection>
<GID>897</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-2896,35,-2879</points>
<intersection>-2896 3</intersection>
<intersection>-2886.5 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-2886.5,38,-2886.5</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-2879,35,-2879</points>
<connection>
<GID>896</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-2896,55.5,-2896</points>
<intersection>35 0</intersection>
<intersection>55.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55.5,-2896,55.5,-2890.5</points>
<connection>
<GID>897</GID>
<name>IN_0</name></connection>
<intersection>-2896 3</intersection></vsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>118,-2887.5,127,-2887.5</points>
<connection>
<GID>900</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>895</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-2897.5,108.5,-2879</points>
<intersection>-2897.5 3</intersection>
<intersection>-2886.5 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-2886.5,112,-2886.5</points>
<connection>
<GID>895</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-2879,108.5,-2879</points>
<connection>
<GID>899</GID>
<name>OUT_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108.5,-2897.5,129,-2897.5</points>
<intersection>108.5 0</intersection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-2897.5,129,-2890.5</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<intersection>-2897.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202,-2889.5,211.5,-2889.5</points>
<connection>
<GID>904</GID>
<name>OUT</name></connection>
<connection>
<GID>903</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-2898,193,-2879</points>
<intersection>-2898 3</intersection>
<intersection>-2888.5 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-2888.5,196,-2888.5</points>
<connection>
<GID>904</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>192,-2879,193,-2879</points>
<connection>
<GID>902</GID>
<name>OUT_0</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>193,-2898,213.5,-2898</points>
<intersection>193 0</intersection>
<intersection>213.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>213.5,-2898,213.5,-2892.5</points>
<connection>
<GID>903</GID>
<name>IN_0</name></connection>
<intersection>-2898 3</intersection></vsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>276,-2889.5,285,-2889.5</points>
<connection>
<GID>906</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>901</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-2899.5,266.5,-2879</points>
<connection>
<GID>905</GID>
<name>OUT_0</name></connection>
<intersection>-2899.5 3</intersection>
<intersection>-2888.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-2888.5,270,-2888.5</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-2899.5,287,-2899.5</points>
<intersection>266.5 0</intersection>
<intersection>287 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>287,-2899.5,287,-2892.5</points>
<connection>
<GID>906</GID>
<name>IN_0</name></connection>
<intersection>-2899.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367,-2891,376.5,-2891</points>
<connection>
<GID>910</GID>
<name>OUT</name></connection>
<connection>
<GID>909</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358,-2899.5,358,-2879</points>
<intersection>-2899.5 3</intersection>
<intersection>-2890 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358,-2890,361,-2890</points>
<connection>
<GID>910</GID>
<name>IN_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357,-2879,358,-2879</points>
<connection>
<GID>908</GID>
<name>OUT_0</name></connection>
<intersection>358 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>358,-2899.5,378.5,-2899.5</points>
<intersection>358 0</intersection>
<intersection>378.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>378.5,-2899.5,378.5,-2894</points>
<connection>
<GID>909</GID>
<name>IN_0</name></connection>
<intersection>-2899.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>441,-2891,450,-2891</points>
<connection>
<GID>912</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>907</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,-2899.5,431.5,-2879</points>
<intersection>-2899.5 3</intersection>
<intersection>-2890 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,-2890,435,-2890</points>
<connection>
<GID>907</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>430.5,-2879,431.5,-2879</points>
<connection>
<GID>911</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>431.5,-2899.5,452,-2899.5</points>
<intersection>431.5 0</intersection>
<intersection>452 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>452,-2899.5,452,-2894</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<intersection>-2899.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>525,-2893,534.5,-2893</points>
<connection>
<GID>916</GID>
<name>OUT</name></connection>
<connection>
<GID>915</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,-2899,516,-2879</points>
<intersection>-2899 3</intersection>
<intersection>-2892 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,-2892,519,-2892</points>
<connection>
<GID>916</GID>
<name>IN_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515,-2879,516,-2879</points>
<connection>
<GID>914</GID>
<name>OUT_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>516,-2899,536.5,-2899</points>
<intersection>516 0</intersection>
<intersection>536.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>536.5,-2899,536.5,-2896</points>
<connection>
<GID>915</GID>
<name>IN_0</name></connection>
<intersection>-2899 3</intersection></vsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>599,-2893,608,-2893</points>
<connection>
<GID>918</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>913</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-2899,589.5,-2879</points>
<intersection>-2899 3</intersection>
<intersection>-2892 1</intersection>
<intersection>-2879 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589.5,-2892,593,-2892</points>
<connection>
<GID>913</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-2879,589.5,-2879</points>
<connection>
<GID>917</GID>
<name>OUT_0</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>589.5,-2899,610,-2899</points>
<intersection>589.5 0</intersection>
<intersection>610 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>610,-2899,610,-2896</points>
<connection>
<GID>918</GID>
<name>IN_0</name></connection>
<intersection>-2899 3</intersection></vsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-2882,582.5,-2882</points>
<connection>
<GID>919</GID>
<name>OUT</name></connection>
<connection>
<GID>917</GID>
<name>clock</name></connection>
<connection>
<GID>914</GID>
<name>clock</name></connection>
<connection>
<GID>911</GID>
<name>clock</name></connection>
<connection>
<GID>908</GID>
<name>clock</name></connection>
<connection>
<GID>905</GID>
<name>clock</name></connection>
<connection>
<GID>902</GID>
<name>clock</name></connection>
<connection>
<GID>899</GID>
<name>clock</name></connection>
<connection>
<GID>896</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-2809,-111,-2585</points>
<intersection>-2809 3</intersection>
<intersection>-2791 1</intersection>
<intersection>-2585 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-2791,-6.5,-2791</points>
<connection>
<GID>945</GID>
<name>IN_0</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-2585,-111,-2585</points>
<connection>
<GID>947</GID>
<name>OUT_1</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111,-2809,-25,-2809</points>
<connection>
<GID>946</GID>
<name>ENABLE_0</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-22.5,-2811,590,-2811</points>
<connection>
<GID>946</GID>
<name>OUT_0</name></connection>
<intersection>35 38</intersection>
<intersection>109 43</intersection>
<intersection>193 42</intersection>
<intersection>267 45</intersection>
<intersection>358 47</intersection>
<intersection>432 49</intersection>
<intersection>516 51</intersection>
<intersection>590 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>35,-2811,35,-2798.5</points>
<connection>
<GID>924</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>193,-2811,193,-2800.5</points>
<connection>
<GID>930</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>109,-2811,109,-2798.5</points>
<connection>
<GID>921</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>267,-2811,267,-2800.5</points>
<connection>
<GID>927</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>358,-2811,358,-2802</points>
<connection>
<GID>936</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>432,-2811,432,-2802</points>
<connection>
<GID>933</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>516,-2811,516,-2804</points>
<connection>
<GID>942</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>590,-2811,590,-2804</points>
<connection>
<GID>939</GID>
<name>IN_1</name></connection>
<intersection>-2811 33</intersection></vsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-2797.5,50.5,-2797.5</points>
<connection>
<GID>924</GID>
<name>OUT</name></connection>
<connection>
<GID>923</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-2806,32,-2789</points>
<intersection>-2806 3</intersection>
<intersection>-2796.5 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-2796.5,35,-2796.5</points>
<connection>
<GID>924</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-2789,32,-2789</points>
<connection>
<GID>922</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-2806,52.5,-2806</points>
<intersection>32 0</intersection>
<intersection>52.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52.5,-2806,52.5,-2800.5</points>
<connection>
<GID>923</GID>
<name>IN_0</name></connection>
<intersection>-2806 3</intersection></vsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115,-2797.5,124,-2797.5</points>
<connection>
<GID>926</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>921</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-2807.5,105.5,-2789</points>
<intersection>-2807.5 3</intersection>
<intersection>-2796.5 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-2796.5,109,-2796.5</points>
<connection>
<GID>921</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-2789,105.5,-2789</points>
<connection>
<GID>925</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105.5,-2807.5,126,-2807.5</points>
<intersection>105.5 0</intersection>
<intersection>126 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,-2807.5,126,-2800.5</points>
<connection>
<GID>926</GID>
<name>IN_0</name></connection>
<intersection>-2807.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-2799.5,208.5,-2799.5</points>
<connection>
<GID>930</GID>
<name>OUT</name></connection>
<connection>
<GID>929</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-2808,190,-2789</points>
<intersection>-2808 3</intersection>
<intersection>-2798.5 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-2798.5,193,-2798.5</points>
<connection>
<GID>930</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,-2789,190,-2789</points>
<connection>
<GID>928</GID>
<name>OUT_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>190,-2808,210.5,-2808</points>
<intersection>190 0</intersection>
<intersection>210.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210.5,-2808,210.5,-2802.5</points>
<connection>
<GID>929</GID>
<name>IN_0</name></connection>
<intersection>-2808 3</intersection></vsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>273,-2799.5,282,-2799.5</points>
<connection>
<GID>932</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>927</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,-2809.5,263.5,-2789</points>
<connection>
<GID>931</GID>
<name>OUT_0</name></connection>
<intersection>-2809.5 3</intersection>
<intersection>-2798.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,-2798.5,267,-2798.5</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263.5,-2809.5,284,-2809.5</points>
<intersection>263.5 0</intersection>
<intersection>284 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>284,-2809.5,284,-2802.5</points>
<connection>
<GID>932</GID>
<name>IN_0</name></connection>
<intersection>-2809.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364,-2801,373.5,-2801</points>
<connection>
<GID>936</GID>
<name>OUT</name></connection>
<connection>
<GID>935</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-2809.5,355,-2789</points>
<intersection>-2809.5 3</intersection>
<intersection>-2800 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-2800,358,-2800</points>
<connection>
<GID>936</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-2789,355,-2789</points>
<connection>
<GID>934</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>355,-2809.5,375.5,-2809.5</points>
<intersection>355 0</intersection>
<intersection>375.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375.5,-2809.5,375.5,-2804</points>
<connection>
<GID>935</GID>
<name>IN_0</name></connection>
<intersection>-2809.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>438,-2801,447,-2801</points>
<connection>
<GID>938</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>933</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,-2809.5,428.5,-2789</points>
<intersection>-2809.5 3</intersection>
<intersection>-2800 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,-2800,432,-2800</points>
<connection>
<GID>933</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,-2789,428.5,-2789</points>
<connection>
<GID>937</GID>
<name>OUT_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428.5,-2809.5,449,-2809.5</points>
<intersection>428.5 0</intersection>
<intersection>449 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>449,-2809.5,449,-2804</points>
<connection>
<GID>938</GID>
<name>IN_0</name></connection>
<intersection>-2809.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>772</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,-2803,531.5,-2803</points>
<connection>
<GID>942</GID>
<name>OUT</name></connection>
<connection>
<GID>941</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,-2809,513,-2789</points>
<intersection>-2809 3</intersection>
<intersection>-2802 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513,-2802,516,-2802</points>
<connection>
<GID>942</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>512,-2789,513,-2789</points>
<connection>
<GID>940</GID>
<name>OUT_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>513,-2809,533.5,-2809</points>
<intersection>513 0</intersection>
<intersection>533.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533.5,-2809,533.5,-2806</points>
<connection>
<GID>941</GID>
<name>IN_0</name></connection>
<intersection>-2809 3</intersection></vsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>596,-2803,605,-2803</points>
<connection>
<GID>944</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>939</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,-2809,586.5,-2789</points>
<intersection>-2809 3</intersection>
<intersection>-2802 1</intersection>
<intersection>-2789 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586.5,-2802,590,-2802</points>
<connection>
<GID>939</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585.5,-2789,586.5,-2789</points>
<connection>
<GID>943</GID>
<name>OUT_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586.5,-2809,607,-2809</points>
<intersection>586.5 0</intersection>
<intersection>607 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>607,-2809,607,-2806</points>
<connection>
<GID>944</GID>
<name>IN_0</name></connection>
<intersection>-2809 3</intersection></vsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-2792,579.5,-2792</points>
<connection>
<GID>945</GID>
<name>OUT</name></connection>
<connection>
<GID>943</GID>
<name>clock</name></connection>
<connection>
<GID>940</GID>
<name>clock</name></connection>
<connection>
<GID>937</GID>
<name>clock</name></connection>
<connection>
<GID>934</GID>
<name>clock</name></connection>
<connection>
<GID>931</GID>
<name>clock</name></connection>
<connection>
<GID>928</GID>
<name>clock</name></connection>
<connection>
<GID>925</GID>
<name>clock</name></connection>
<connection>
<GID>922</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-3474,-110,-3231</points>
<intersection>-3474 2</intersection>
<intersection>-3249 3</intersection>
<intersection>-3231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-3231,-8.5,-3231</points>
<connection>
<GID>1111</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3474,-110,-3474</points>
<connection>
<GID>1295</GID>
<name>OUT_6</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-3249,-27,-3249</points>
<connection>
<GID>1112</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-24.5,-3251,588,-3251</points>
<connection>
<GID>1112</GID>
<name>OUT_0</name></connection>
<intersection>33 38</intersection>
<intersection>107 43</intersection>
<intersection>191 42</intersection>
<intersection>265 45</intersection>
<intersection>356 47</intersection>
<intersection>430 49</intersection>
<intersection>514 51</intersection>
<intersection>588 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>33,-3251,33,-3238.5</points>
<connection>
<GID>1090</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>191,-3251,191,-3240.5</points>
<connection>
<GID>1096</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>107,-3251,107,-3238.5</points>
<connection>
<GID>1087</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>265,-3251,265,-3240.5</points>
<connection>
<GID>1093</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>356,-3251,356,-3242</points>
<connection>
<GID>1102</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>430,-3251,430,-3242</points>
<connection>
<GID>1099</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>514,-3251,514,-3244</points>
<connection>
<GID>1108</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>588,-3251,588,-3244</points>
<connection>
<GID>1105</GID>
<name>IN_1</name></connection>
<intersection>-3251 33</intersection></vsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-3237.5,48.5,-3237.5</points>
<connection>
<GID>1090</GID>
<name>OUT</name></connection>
<connection>
<GID>1089</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-3246,30,-3229</points>
<intersection>-3246 3</intersection>
<intersection>-3236.5 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-3236.5,33,-3236.5</points>
<connection>
<GID>1090</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-3229,30,-3229</points>
<connection>
<GID>1088</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30,-3246,50.5,-3246</points>
<intersection>30 0</intersection>
<intersection>50.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50.5,-3246,50.5,-3240.5</points>
<connection>
<GID>1089</GID>
<name>IN_0</name></connection>
<intersection>-3246 3</intersection></vsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113,-3237.5,122,-3237.5</points>
<connection>
<GID>1087</GID>
<name>OUT</name></connection>
<connection>
<GID>1092</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-3247.5,103.5,-3229</points>
<intersection>-3247.5 3</intersection>
<intersection>-3236.5 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-3236.5,107,-3236.5</points>
<connection>
<GID>1087</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-3229,103.5,-3229</points>
<connection>
<GID>1091</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,-3247.5,124,-3247.5</points>
<intersection>103.5 0</intersection>
<intersection>124 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124,-3247.5,124,-3240.5</points>
<connection>
<GID>1092</GID>
<name>IN_0</name></connection>
<intersection>-3247.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-3239.5,206.5,-3239.5</points>
<connection>
<GID>1096</GID>
<name>OUT</name></connection>
<connection>
<GID>1095</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-3248,188,-3229</points>
<intersection>-3248 3</intersection>
<intersection>-3238.5 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188,-3238.5,191,-3238.5</points>
<connection>
<GID>1096</GID>
<name>IN_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-3229,188,-3229</points>
<connection>
<GID>1094</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188,-3248,208.5,-3248</points>
<intersection>188 0</intersection>
<intersection>208.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208.5,-3248,208.5,-3242.5</points>
<connection>
<GID>1095</GID>
<name>IN_0</name></connection>
<intersection>-3248 3</intersection></vsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>271,-3239.5,280,-3239.5</points>
<connection>
<GID>1093</GID>
<name>OUT</name></connection>
<connection>
<GID>1098</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-3249.5,261.5,-3229</points>
<connection>
<GID>1097</GID>
<name>OUT_0</name></connection>
<intersection>-3249.5 3</intersection>
<intersection>-3238.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-3238.5,265,-3238.5</points>
<connection>
<GID>1093</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-3249.5,282,-3249.5</points>
<intersection>261.5 0</intersection>
<intersection>282 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282,-3249.5,282,-3242.5</points>
<connection>
<GID>1098</GID>
<name>IN_0</name></connection>
<intersection>-3249.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362,-3241,371.5,-3241</points>
<connection>
<GID>1102</GID>
<name>OUT</name></connection>
<connection>
<GID>1101</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-3249.5,353,-3229</points>
<intersection>-3249.5 3</intersection>
<intersection>-3240 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-3240,356,-3240</points>
<connection>
<GID>1102</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-3229,353,-3229</points>
<connection>
<GID>1100</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353,-3249.5,373.5,-3249.5</points>
<intersection>353 0</intersection>
<intersection>373.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>373.5,-3249.5,373.5,-3244</points>
<connection>
<GID>1101</GID>
<name>IN_0</name></connection>
<intersection>-3249.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>436,-3241,445,-3241</points>
<connection>
<GID>1099</GID>
<name>OUT</name></connection>
<connection>
<GID>1104</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-3249.5,426.5,-3229</points>
<intersection>-3249.5 3</intersection>
<intersection>-3240 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426.5,-3240,430,-3240</points>
<connection>
<GID>1099</GID>
<name>IN_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425.5,-3229,426.5,-3229</points>
<connection>
<GID>1103</GID>
<name>OUT_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426.5,-3249.5,447,-3249.5</points>
<intersection>426.5 0</intersection>
<intersection>447 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447,-3249.5,447,-3244</points>
<connection>
<GID>1104</GID>
<name>IN_0</name></connection>
<intersection>-3249.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520,-3243,529.5,-3243</points>
<connection>
<GID>1108</GID>
<name>OUT</name></connection>
<connection>
<GID>1107</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,-3249,511,-3229</points>
<intersection>-3249 3</intersection>
<intersection>-3242 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,-3242,514,-3242</points>
<connection>
<GID>1108</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>510,-3229,511,-3229</points>
<connection>
<GID>1106</GID>
<name>OUT_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511,-3249,531.5,-3249</points>
<intersection>511 0</intersection>
<intersection>531.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531.5,-3249,531.5,-3246</points>
<connection>
<GID>1107</GID>
<name>IN_0</name></connection>
<intersection>-3249 3</intersection></vsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>594,-3243,603,-3243</points>
<connection>
<GID>1105</GID>
<name>OUT</name></connection>
<connection>
<GID>1110</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,-3249,584.5,-3229</points>
<intersection>-3249 3</intersection>
<intersection>-3242 1</intersection>
<intersection>-3229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584.5,-3242,588,-3242</points>
<connection>
<GID>1105</GID>
<name>IN_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583.5,-3229,584.5,-3229</points>
<connection>
<GID>1109</GID>
<name>OUT_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>584.5,-3249,605,-3249</points>
<intersection>584.5 0</intersection>
<intersection>605 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>605,-3249,605,-3246</points>
<connection>
<GID>1110</GID>
<name>IN_0</name></connection>
<intersection>-3249 3</intersection></vsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-3232,577.5,-3232</points>
<connection>
<GID>1111</GID>
<name>OUT</name></connection>
<connection>
<GID>1109</GID>
<name>clock</name></connection>
<connection>
<GID>1106</GID>
<name>clock</name></connection>
<connection>
<GID>1103</GID>
<name>clock</name></connection>
<connection>
<GID>1100</GID>
<name>clock</name></connection>
<connection>
<GID>1097</GID>
<name>clock</name></connection>
<connection>
<GID>1094</GID>
<name>clock</name></connection>
<connection>
<GID>1091</GID>
<name>clock</name></connection>
<connection>
<GID>1088</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-3473,-111,-3141</points>
<intersection>-3473 2</intersection>
<intersection>-3159 3</intersection>
<intersection>-3141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-3141,-11.5,-3141</points>
<connection>
<GID>1137</GID>
<name>IN_0</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3473,-111,-3473</points>
<connection>
<GID>1295</GID>
<name>OUT_7</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111,-3159,-30,-3159</points>
<connection>
<GID>1138</GID>
<name>ENABLE_0</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-27.5,-3161,585,-3161</points>
<connection>
<GID>1138</GID>
<name>OUT_0</name></connection>
<intersection>30 38</intersection>
<intersection>104 43</intersection>
<intersection>188 42</intersection>
<intersection>262 45</intersection>
<intersection>353 47</intersection>
<intersection>427 49</intersection>
<intersection>511 51</intersection>
<intersection>585 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>30,-3161,30,-3148.5</points>
<connection>
<GID>1116</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>188,-3161,188,-3150.5</points>
<connection>
<GID>1122</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>104,-3161,104,-3148.5</points>
<connection>
<GID>1113</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>262,-3161,262,-3150.5</points>
<connection>
<GID>1119</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>353,-3161,353,-3152</points>
<connection>
<GID>1128</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>427,-3161,427,-3152</points>
<connection>
<GID>1125</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>511,-3161,511,-3154</points>
<connection>
<GID>1134</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>585,-3161,585,-3154</points>
<connection>
<GID>1131</GID>
<name>IN_1</name></connection>
<intersection>-3161 33</intersection></vsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-3147.5,45.5,-3147.5</points>
<connection>
<GID>1116</GID>
<name>OUT</name></connection>
<connection>
<GID>1115</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-3156,27,-3139</points>
<intersection>-3156 3</intersection>
<intersection>-3146.5 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-3146.5,30,-3146.5</points>
<connection>
<GID>1116</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-3139,27,-3139</points>
<connection>
<GID>1114</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-3156,47.5,-3156</points>
<intersection>27 0</intersection>
<intersection>47.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-3156,47.5,-3150.5</points>
<connection>
<GID>1115</GID>
<name>IN_0</name></connection>
<intersection>-3156 3</intersection></vsegment></shape></wire>
<wire>
<ID>800</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>110,-3147.5,119,-3147.5</points>
<connection>
<GID>1113</GID>
<name>OUT</name></connection>
<connection>
<GID>1118</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-3157.5,100.5,-3139</points>
<intersection>-3157.5 3</intersection>
<intersection>-3146.5 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-3146.5,104,-3146.5</points>
<connection>
<GID>1113</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-3139,100.5,-3139</points>
<connection>
<GID>1117</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100.5,-3157.5,121,-3157.5</points>
<intersection>100.5 0</intersection>
<intersection>121 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>121,-3157.5,121,-3150.5</points>
<connection>
<GID>1118</GID>
<name>IN_0</name></connection>
<intersection>-3157.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,-3149.5,203.5,-3149.5</points>
<connection>
<GID>1122</GID>
<name>OUT</name></connection>
<connection>
<GID>1121</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-3158,185,-3139</points>
<intersection>-3158 3</intersection>
<intersection>-3148.5 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-3148.5,188,-3148.5</points>
<connection>
<GID>1122</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-3139,185,-3139</points>
<connection>
<GID>1120</GID>
<name>OUT_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185,-3158,205.5,-3158</points>
<intersection>185 0</intersection>
<intersection>205.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>205.5,-3158,205.5,-3152.5</points>
<connection>
<GID>1121</GID>
<name>IN_0</name></connection>
<intersection>-3158 3</intersection></vsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>268,-3149.5,277,-3149.5</points>
<connection>
<GID>1119</GID>
<name>OUT</name></connection>
<connection>
<GID>1124</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>805</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-3159.5,258.5,-3139</points>
<connection>
<GID>1123</GID>
<name>OUT_0</name></connection>
<intersection>-3159.5 3</intersection>
<intersection>-3148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,-3148.5,262,-3148.5</points>
<connection>
<GID>1119</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,-3159.5,279,-3159.5</points>
<intersection>258.5 0</intersection>
<intersection>279 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>279,-3159.5,279,-3152.5</points>
<connection>
<GID>1124</GID>
<name>IN_0</name></connection>
<intersection>-3159.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-3151,368.5,-3151</points>
<connection>
<GID>1128</GID>
<name>OUT</name></connection>
<connection>
<GID>1127</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-3159.5,350,-3139</points>
<intersection>-3159.5 3</intersection>
<intersection>-3150 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-3150,353,-3150</points>
<connection>
<GID>1128</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-3139,350,-3139</points>
<connection>
<GID>1126</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>350,-3159.5,370.5,-3159.5</points>
<intersection>350 0</intersection>
<intersection>370.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>370.5,-3159.5,370.5,-3154</points>
<connection>
<GID>1127</GID>
<name>IN_0</name></connection>
<intersection>-3159.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>808</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>433,-3151,442,-3151</points>
<connection>
<GID>1125</GID>
<name>OUT</name></connection>
<connection>
<GID>1130</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-3159.5,423.5,-3139</points>
<intersection>-3159.5 3</intersection>
<intersection>-3150 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423.5,-3150,427,-3150</points>
<connection>
<GID>1125</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422.5,-3139,423.5,-3139</points>
<connection>
<GID>1129</GID>
<name>OUT_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>423.5,-3159.5,444,-3159.5</points>
<intersection>423.5 0</intersection>
<intersection>444 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>444,-3159.5,444,-3154</points>
<connection>
<GID>1130</GID>
<name>IN_0</name></connection>
<intersection>-3159.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>517,-3153,526.5,-3153</points>
<connection>
<GID>1134</GID>
<name>OUT</name></connection>
<connection>
<GID>1133</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508,-3159,508,-3139</points>
<intersection>-3159 3</intersection>
<intersection>-3152 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,-3152,511,-3152</points>
<connection>
<GID>1134</GID>
<name>IN_0</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507,-3139,508,-3139</points>
<connection>
<GID>1132</GID>
<name>OUT_0</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>508,-3159,528.5,-3159</points>
<intersection>508 0</intersection>
<intersection>528.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>528.5,-3159,528.5,-3156</points>
<connection>
<GID>1133</GID>
<name>IN_0</name></connection>
<intersection>-3159 3</intersection></vsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>591,-3153,600,-3153</points>
<connection>
<GID>1131</GID>
<name>OUT</name></connection>
<connection>
<GID>1136</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581.5,-3159,581.5,-3139</points>
<intersection>-3159 3</intersection>
<intersection>-3152 1</intersection>
<intersection>-3139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581.5,-3152,585,-3152</points>
<connection>
<GID>1131</GID>
<name>IN_0</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>580.5,-3139,581.5,-3139</points>
<connection>
<GID>1135</GID>
<name>OUT_0</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>581.5,-3159,602,-3159</points>
<intersection>581.5 0</intersection>
<intersection>602 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>602,-3159,602,-3156</points>
<connection>
<GID>1136</GID>
<name>IN_0</name></connection>
<intersection>-3159 3</intersection></vsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-3142,574.5,-3142</points>
<connection>
<GID>1137</GID>
<name>OUT</name></connection>
<connection>
<GID>1135</GID>
<name>clock</name></connection>
<connection>
<GID>1132</GID>
<name>clock</name></connection>
<connection>
<GID>1129</GID>
<name>clock</name></connection>
<connection>
<GID>1126</GID>
<name>clock</name></connection>
<connection>
<GID>1123</GID>
<name>clock</name></connection>
<connection>
<GID>1120</GID>
<name>clock</name></connection>
<connection>
<GID>1117</GID>
<name>clock</name></connection>
<connection>
<GID>1114</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-3476,-108,-3399</points>
<intersection>-3476 2</intersection>
<intersection>-3417 3</intersection>
<intersection>-3399 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-3399,-4.5,-3399</points>
<connection>
<GID>1163</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3476,-108,-3476</points>
<connection>
<GID>1295</GID>
<name>OUT_4</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-3417,-23,-3417</points>
<connection>
<GID>1164</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>816</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-20.5,-3419,592,-3419</points>
<connection>
<GID>1164</GID>
<name>OUT_0</name></connection>
<intersection>37 38</intersection>
<intersection>111 43</intersection>
<intersection>195 42</intersection>
<intersection>269 45</intersection>
<intersection>360 47</intersection>
<intersection>434 49</intersection>
<intersection>518 51</intersection>
<intersection>592 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>37,-3419,37,-3406.5</points>
<connection>
<GID>1142</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>195,-3419,195,-3408.5</points>
<connection>
<GID>1148</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>111,-3419,111,-3406.5</points>
<connection>
<GID>1139</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>269,-3419,269,-3408.5</points>
<connection>
<GID>1145</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>360,-3419,360,-3410</points>
<connection>
<GID>1154</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>434,-3419,434,-3410</points>
<connection>
<GID>1151</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>518,-3419,518,-3412</points>
<connection>
<GID>1160</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>592,-3419,592,-3412</points>
<connection>
<GID>1157</GID>
<name>IN_1</name></connection>
<intersection>-3419 33</intersection></vsegment></shape></wire>
<wire>
<ID>817</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-3405.5,52.5,-3405.5</points>
<connection>
<GID>1142</GID>
<name>OUT</name></connection>
<connection>
<GID>1141</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-3414,34,-3397</points>
<intersection>-3414 3</intersection>
<intersection>-3404.5 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-3404.5,37,-3404.5</points>
<connection>
<GID>1142</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-3397,34,-3397</points>
<connection>
<GID>1140</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-3414,54.5,-3414</points>
<intersection>34 0</intersection>
<intersection>54.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54.5,-3414,54.5,-3408.5</points>
<connection>
<GID>1141</GID>
<name>IN_0</name></connection>
<intersection>-3414 3</intersection></vsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>117,-3405.5,126,-3405.5</points>
<connection>
<GID>1139</GID>
<name>OUT</name></connection>
<connection>
<GID>1144</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-3415.5,107.5,-3397</points>
<intersection>-3415.5 3</intersection>
<intersection>-3404.5 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-3404.5,111,-3404.5</points>
<connection>
<GID>1139</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-3397,107.5,-3397</points>
<connection>
<GID>1143</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-3415.5,128,-3415.5</points>
<intersection>107.5 0</intersection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-3415.5,128,-3408.5</points>
<connection>
<GID>1144</GID>
<name>IN_0</name></connection>
<intersection>-3415.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201,-3407.5,210.5,-3407.5</points>
<connection>
<GID>1148</GID>
<name>OUT</name></connection>
<connection>
<GID>1147</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-3416,192,-3397</points>
<intersection>-3416 3</intersection>
<intersection>-3406.5 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-3406.5,195,-3406.5</points>
<connection>
<GID>1148</GID>
<name>IN_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-3397,192,-3397</points>
<connection>
<GID>1146</GID>
<name>OUT_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>192,-3416,212.5,-3416</points>
<intersection>192 0</intersection>
<intersection>212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>212.5,-3416,212.5,-3410.5</points>
<connection>
<GID>1147</GID>
<name>IN_0</name></connection>
<intersection>-3416 3</intersection></vsegment></shape></wire>
<wire>
<ID>823</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>275,-3407.5,284,-3407.5</points>
<connection>
<GID>1145</GID>
<name>OUT</name></connection>
<connection>
<GID>1150</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-3417.5,265.5,-3397</points>
<connection>
<GID>1149</GID>
<name>OUT_0</name></connection>
<intersection>-3417.5 3</intersection>
<intersection>-3406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,-3406.5,269,-3406.5</points>
<connection>
<GID>1145</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>265.5,-3417.5,286,-3417.5</points>
<intersection>265.5 0</intersection>
<intersection>286 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>286,-3417.5,286,-3410.5</points>
<connection>
<GID>1150</GID>
<name>IN_0</name></connection>
<intersection>-3417.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366,-3409,375.5,-3409</points>
<connection>
<GID>1154</GID>
<name>OUT</name></connection>
<connection>
<GID>1153</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-3417.5,357,-3397</points>
<intersection>-3417.5 3</intersection>
<intersection>-3408 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-3408,360,-3408</points>
<connection>
<GID>1154</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356,-3397,357,-3397</points>
<connection>
<GID>1152</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-3417.5,377.5,-3417.5</points>
<intersection>357 0</intersection>
<intersection>377.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>377.5,-3417.5,377.5,-3412</points>
<connection>
<GID>1153</GID>
<name>IN_0</name></connection>
<intersection>-3417.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>440,-3409,449,-3409</points>
<connection>
<GID>1151</GID>
<name>OUT</name></connection>
<connection>
<GID>1156</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,-3417.5,430.5,-3397</points>
<intersection>-3417.5 3</intersection>
<intersection>-3408 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430.5,-3408,434,-3408</points>
<connection>
<GID>1151</GID>
<name>IN_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>429.5,-3397,430.5,-3397</points>
<connection>
<GID>1155</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>430.5,-3417.5,451,-3417.5</points>
<intersection>430.5 0</intersection>
<intersection>451 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>451,-3417.5,451,-3412</points>
<connection>
<GID>1156</GID>
<name>IN_0</name></connection>
<intersection>-3417.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524,-3411,533.5,-3411</points>
<connection>
<GID>1160</GID>
<name>OUT</name></connection>
<connection>
<GID>1159</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-3417,515,-3397</points>
<intersection>-3417 3</intersection>
<intersection>-3410 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515,-3410,518,-3410</points>
<connection>
<GID>1160</GID>
<name>IN_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,-3397,515,-3397</points>
<connection>
<GID>1158</GID>
<name>OUT_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>515,-3417,535.5,-3417</points>
<intersection>515 0</intersection>
<intersection>535.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535.5,-3417,535.5,-3414</points>
<connection>
<GID>1159</GID>
<name>IN_0</name></connection>
<intersection>-3417 3</intersection></vsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>598,-3411,607,-3411</points>
<connection>
<GID>1157</GID>
<name>OUT</name></connection>
<connection>
<GID>1162</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588.5,-3417,588.5,-3397</points>
<intersection>-3417 3</intersection>
<intersection>-3410 1</intersection>
<intersection>-3397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588.5,-3410,592,-3410</points>
<connection>
<GID>1157</GID>
<name>IN_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-3397,588.5,-3397</points>
<connection>
<GID>1161</GID>
<name>OUT_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>588.5,-3417,609,-3417</points>
<intersection>588.5 0</intersection>
<intersection>609 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>609,-3417,609,-3414</points>
<connection>
<GID>1162</GID>
<name>IN_0</name></connection>
<intersection>-3417 3</intersection></vsegment></shape></wire>
<wire>
<ID>833</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-3400,581.5,-3400</points>
<connection>
<GID>1163</GID>
<name>OUT</name></connection>
<connection>
<GID>1161</GID>
<name>clock</name></connection>
<connection>
<GID>1158</GID>
<name>clock</name></connection>
<connection>
<GID>1155</GID>
<name>clock</name></connection>
<connection>
<GID>1152</GID>
<name>clock</name></connection>
<connection>
<GID>1149</GID>
<name>clock</name></connection>
<connection>
<GID>1146</GID>
<name>clock</name></connection>
<connection>
<GID>1143</GID>
<name>clock</name></connection>
<connection>
<GID>1140</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>834</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-3475,-109,-3309</points>
<intersection>-3475 2</intersection>
<intersection>-3327 3</intersection>
<intersection>-3309 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-3309,-7.5,-3309</points>
<connection>
<GID>1189</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3475,-109,-3475</points>
<connection>
<GID>1295</GID>
<name>OUT_5</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-3327,-26,-3327</points>
<connection>
<GID>1190</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-3329,589,-3329</points>
<connection>
<GID>1190</GID>
<name>OUT_0</name></connection>
<intersection>34 38</intersection>
<intersection>108 43</intersection>
<intersection>192 42</intersection>
<intersection>266 45</intersection>
<intersection>357 47</intersection>
<intersection>431 49</intersection>
<intersection>515 51</intersection>
<intersection>589 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34,-3329,34,-3316.5</points>
<connection>
<GID>1168</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192,-3329,192,-3318.5</points>
<connection>
<GID>1174</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108,-3329,108,-3316.5</points>
<connection>
<GID>1165</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266,-3329,266,-3318.5</points>
<connection>
<GID>1171</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357,-3329,357,-3320</points>
<connection>
<GID>1180</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431,-3329,431,-3320</points>
<connection>
<GID>1177</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515,-3329,515,-3322</points>
<connection>
<GID>1186</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589,-3329,589,-3322</points>
<connection>
<GID>1183</GID>
<name>IN_1</name></connection>
<intersection>-3329 33</intersection></vsegment></shape></wire>
<wire>
<ID>836</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-3315.5,49.5,-3315.5</points>
<connection>
<GID>1168</GID>
<name>OUT</name></connection>
<connection>
<GID>1167</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-3324,31,-3307</points>
<intersection>-3324 3</intersection>
<intersection>-3314.5 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-3314.5,34,-3314.5</points>
<connection>
<GID>1168</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-3307,31,-3307</points>
<connection>
<GID>1166</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-3324,51.5,-3324</points>
<intersection>31 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-3324,51.5,-3318.5</points>
<connection>
<GID>1167</GID>
<name>IN_0</name></connection>
<intersection>-3324 3</intersection></vsegment></shape></wire>
<wire>
<ID>838</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114,-3315.5,123,-3315.5</points>
<connection>
<GID>1165</GID>
<name>OUT</name></connection>
<connection>
<GID>1170</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-3325.5,104.5,-3307</points>
<intersection>-3325.5 3</intersection>
<intersection>-3314.5 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-3314.5,108,-3314.5</points>
<connection>
<GID>1165</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-3307,104.5,-3307</points>
<connection>
<GID>1169</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-3325.5,125,-3325.5</points>
<intersection>104.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-3325.5,125,-3318.5</points>
<connection>
<GID>1170</GID>
<name>IN_0</name></connection>
<intersection>-3325.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>840</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-3317.5,207.5,-3317.5</points>
<connection>
<GID>1174</GID>
<name>OUT</name></connection>
<connection>
<GID>1173</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-3326,189,-3307</points>
<intersection>-3326 3</intersection>
<intersection>-3316.5 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-3316.5,192,-3316.5</points>
<connection>
<GID>1174</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188,-3307,189,-3307</points>
<connection>
<GID>1172</GID>
<name>OUT_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189,-3326,209.5,-3326</points>
<intersection>189 0</intersection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,-3326,209.5,-3320.5</points>
<connection>
<GID>1173</GID>
<name>IN_0</name></connection>
<intersection>-3326 3</intersection></vsegment></shape></wire>
<wire>
<ID>842</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272,-3317.5,281,-3317.5</points>
<connection>
<GID>1171</GID>
<name>OUT</name></connection>
<connection>
<GID>1176</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>843</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-3327.5,262.5,-3307</points>
<connection>
<GID>1175</GID>
<name>OUT_0</name></connection>
<intersection>-3327.5 3</intersection>
<intersection>-3316.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-3316.5,266,-3316.5</points>
<connection>
<GID>1171</GID>
<name>IN_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262.5,-3327.5,283,-3327.5</points>
<intersection>262.5 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-3327.5,283,-3320.5</points>
<connection>
<GID>1176</GID>
<name>IN_0</name></connection>
<intersection>-3327.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>844</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363,-3319,372.5,-3319</points>
<connection>
<GID>1180</GID>
<name>OUT</name></connection>
<connection>
<GID>1179</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-3327.5,354,-3307</points>
<intersection>-3327.5 3</intersection>
<intersection>-3318 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-3318,357,-3318</points>
<connection>
<GID>1180</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-3307,354,-3307</points>
<connection>
<GID>1178</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354,-3327.5,374.5,-3327.5</points>
<intersection>354 0</intersection>
<intersection>374.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374.5,-3327.5,374.5,-3322</points>
<connection>
<GID>1179</GID>
<name>IN_0</name></connection>
<intersection>-3327.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>846</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437,-3319,446,-3319</points>
<connection>
<GID>1177</GID>
<name>OUT</name></connection>
<connection>
<GID>1182</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-3327.5,427.5,-3307</points>
<intersection>-3327.5 3</intersection>
<intersection>-3318 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-3318,431,-3318</points>
<connection>
<GID>1177</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426.5,-3307,427.5,-3307</points>
<connection>
<GID>1181</GID>
<name>OUT_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-3327.5,448,-3327.5</points>
<intersection>427.5 0</intersection>
<intersection>448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448,-3327.5,448,-3322</points>
<connection>
<GID>1182</GID>
<name>IN_0</name></connection>
<intersection>-3327.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521,-3321,530.5,-3321</points>
<connection>
<GID>1186</GID>
<name>OUT</name></connection>
<connection>
<GID>1185</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,-3327,512,-3307</points>
<intersection>-3327 3</intersection>
<intersection>-3320 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-3320,515,-3320</points>
<connection>
<GID>1186</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,-3307,512,-3307</points>
<connection>
<GID>1184</GID>
<name>OUT_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512,-3327,532.5,-3327</points>
<intersection>512 0</intersection>
<intersection>532.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532.5,-3327,532.5,-3324</points>
<connection>
<GID>1185</GID>
<name>IN_0</name></connection>
<intersection>-3327 3</intersection></vsegment></shape></wire>
<wire>
<ID>850</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595,-3321,604,-3321</points>
<connection>
<GID>1183</GID>
<name>OUT</name></connection>
<connection>
<GID>1188</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-3327,585.5,-3307</points>
<intersection>-3327 3</intersection>
<intersection>-3320 1</intersection>
<intersection>-3307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-3320,589,-3320</points>
<connection>
<GID>1183</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,-3307,585.5,-3307</points>
<connection>
<GID>1187</GID>
<name>OUT_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-3327,606,-3327</points>
<intersection>585.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-3327,606,-3324</points>
<connection>
<GID>1188</GID>
<name>IN_0</name></connection>
<intersection>-3327 3</intersection></vsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-3310,578.5,-3310</points>
<connection>
<GID>1189</GID>
<name>OUT</name></connection>
<connection>
<GID>1187</GID>
<name>clock</name></connection>
<connection>
<GID>1184</GID>
<name>clock</name></connection>
<connection>
<GID>1181</GID>
<name>clock</name></connection>
<connection>
<GID>1178</GID>
<name>clock</name></connection>
<connection>
<GID>1175</GID>
<name>clock</name></connection>
<connection>
<GID>1172</GID>
<name>clock</name></connection>
<connection>
<GID>1169</GID>
<name>clock</name></connection>
<connection>
<GID>1166</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>853</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-3625,-109,-3478</points>
<intersection>-3625 3</intersection>
<intersection>-3607 1</intersection>
<intersection>-3478 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-3607,-6.5,-3607</points>
<connection>
<GID>1215</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3478,-109,-3478</points>
<connection>
<GID>1295</GID>
<name>OUT_2</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-3625,-25,-3625</points>
<connection>
<GID>1216</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-22.5,-3627,590,-3627</points>
<connection>
<GID>1216</GID>
<name>OUT_0</name></connection>
<intersection>35 38</intersection>
<intersection>109 43</intersection>
<intersection>193 42</intersection>
<intersection>267 45</intersection>
<intersection>358 47</intersection>
<intersection>432 49</intersection>
<intersection>516 51</intersection>
<intersection>590 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>35,-3627,35,-3614.5</points>
<connection>
<GID>1194</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>193,-3627,193,-3616.5</points>
<connection>
<GID>1200</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>109,-3627,109,-3614.5</points>
<connection>
<GID>1191</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>267,-3627,267,-3616.5</points>
<connection>
<GID>1197</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>358,-3627,358,-3618</points>
<connection>
<GID>1206</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>432,-3627,432,-3618</points>
<connection>
<GID>1203</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>516,-3627,516,-3620</points>
<connection>
<GID>1212</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>590,-3627,590,-3620</points>
<connection>
<GID>1209</GID>
<name>IN_1</name></connection>
<intersection>-3627 33</intersection></vsegment></shape></wire>
<wire>
<ID>855</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-3613.5,50.5,-3613.5</points>
<connection>
<GID>1194</GID>
<name>OUT</name></connection>
<connection>
<GID>1193</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-3622,32,-3605</points>
<intersection>-3622 3</intersection>
<intersection>-3612.5 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-3612.5,35,-3612.5</points>
<connection>
<GID>1194</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-3605,32,-3605</points>
<connection>
<GID>1192</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-3622,52.5,-3622</points>
<intersection>32 0</intersection>
<intersection>52.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52.5,-3622,52.5,-3616.5</points>
<connection>
<GID>1193</GID>
<name>IN_0</name></connection>
<intersection>-3622 3</intersection></vsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115,-3613.5,124,-3613.5</points>
<connection>
<GID>1191</GID>
<name>OUT</name></connection>
<connection>
<GID>1196</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-3623.5,105.5,-3605</points>
<intersection>-3623.5 3</intersection>
<intersection>-3612.5 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-3612.5,109,-3612.5</points>
<connection>
<GID>1191</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-3605,105.5,-3605</points>
<connection>
<GID>1195</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105.5,-3623.5,126,-3623.5</points>
<intersection>105.5 0</intersection>
<intersection>126 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,-3623.5,126,-3616.5</points>
<connection>
<GID>1196</GID>
<name>IN_0</name></connection>
<intersection>-3623.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-3615.5,208.5,-3615.5</points>
<connection>
<GID>1200</GID>
<name>OUT</name></connection>
<connection>
<GID>1199</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-3624,190,-3605</points>
<intersection>-3624 3</intersection>
<intersection>-3614.5 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-3614.5,193,-3614.5</points>
<connection>
<GID>1200</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,-3605,190,-3605</points>
<connection>
<GID>1198</GID>
<name>OUT_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>190,-3624,210.5,-3624</points>
<intersection>190 0</intersection>
<intersection>210.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210.5,-3624,210.5,-3618.5</points>
<connection>
<GID>1199</GID>
<name>IN_0</name></connection>
<intersection>-3624 3</intersection></vsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>273,-3615.5,282,-3615.5</points>
<connection>
<GID>1197</GID>
<name>OUT</name></connection>
<connection>
<GID>1202</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,-3625.5,263.5,-3605</points>
<connection>
<GID>1201</GID>
<name>OUT_0</name></connection>
<intersection>-3625.5 3</intersection>
<intersection>-3614.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,-3614.5,267,-3614.5</points>
<connection>
<GID>1197</GID>
<name>IN_0</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263.5,-3625.5,284,-3625.5</points>
<intersection>263.5 0</intersection>
<intersection>284 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>284,-3625.5,284,-3618.5</points>
<connection>
<GID>1202</GID>
<name>IN_0</name></connection>
<intersection>-3625.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>863</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364,-3617,373.5,-3617</points>
<connection>
<GID>1206</GID>
<name>OUT</name></connection>
<connection>
<GID>1205</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>864</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-3625.5,355,-3605</points>
<intersection>-3625.5 3</intersection>
<intersection>-3616 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-3616,358,-3616</points>
<connection>
<GID>1206</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-3605,355,-3605</points>
<connection>
<GID>1204</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>355,-3625.5,375.5,-3625.5</points>
<intersection>355 0</intersection>
<intersection>375.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375.5,-3625.5,375.5,-3620</points>
<connection>
<GID>1205</GID>
<name>IN_0</name></connection>
<intersection>-3625.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>865</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>438,-3617,447,-3617</points>
<connection>
<GID>1203</GID>
<name>OUT</name></connection>
<connection>
<GID>1208</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>866</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,-3625.5,428.5,-3605</points>
<intersection>-3625.5 3</intersection>
<intersection>-3616 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,-3616,432,-3616</points>
<connection>
<GID>1203</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,-3605,428.5,-3605</points>
<connection>
<GID>1207</GID>
<name>OUT_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428.5,-3625.5,449,-3625.5</points>
<intersection>428.5 0</intersection>
<intersection>449 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>449,-3625.5,449,-3620</points>
<connection>
<GID>1208</GID>
<name>IN_0</name></connection>
<intersection>-3625.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>867</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,-3619,531.5,-3619</points>
<connection>
<GID>1212</GID>
<name>OUT</name></connection>
<connection>
<GID>1211</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,-3625,513,-3605</points>
<intersection>-3625 3</intersection>
<intersection>-3618 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513,-3618,516,-3618</points>
<connection>
<GID>1212</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>512,-3605,513,-3605</points>
<connection>
<GID>1210</GID>
<name>OUT_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>513,-3625,533.5,-3625</points>
<intersection>513 0</intersection>
<intersection>533.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533.5,-3625,533.5,-3622</points>
<connection>
<GID>1211</GID>
<name>IN_0</name></connection>
<intersection>-3625 3</intersection></vsegment></shape></wire>
<wire>
<ID>869</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>596,-3619,605,-3619</points>
<connection>
<GID>1209</GID>
<name>OUT</name></connection>
<connection>
<GID>1214</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,-3625,586.5,-3605</points>
<intersection>-3625 3</intersection>
<intersection>-3618 1</intersection>
<intersection>-3605 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586.5,-3618,590,-3618</points>
<connection>
<GID>1209</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585.5,-3605,586.5,-3605</points>
<connection>
<GID>1213</GID>
<name>OUT_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586.5,-3625,607,-3625</points>
<intersection>586.5 0</intersection>
<intersection>607 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>607,-3625,607,-3622</points>
<connection>
<GID>1214</GID>
<name>IN_0</name></connection>
<intersection>-3625 3</intersection></vsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-3608,579.5,-3608</points>
<connection>
<GID>1215</GID>
<name>OUT</name></connection>
<connection>
<GID>1213</GID>
<name>clock</name></connection>
<connection>
<GID>1210</GID>
<name>clock</name></connection>
<connection>
<GID>1207</GID>
<name>clock</name></connection>
<connection>
<GID>1204</GID>
<name>clock</name></connection>
<connection>
<GID>1201</GID>
<name>clock</name></connection>
<connection>
<GID>1198</GID>
<name>clock</name></connection>
<connection>
<GID>1195</GID>
<name>clock</name></connection>
<connection>
<GID>1192</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-3535,-108,-3477</points>
<intersection>-3535 3</intersection>
<intersection>-3517 1</intersection>
<intersection>-3477 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-3517,-9.5,-3517</points>
<connection>
<GID>1241</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3477,-108,-3477</points>
<connection>
<GID>1295</GID>
<name>OUT_3</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-3535,-28,-3535</points>
<connection>
<GID>1242</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25.5,-3537,587,-3537</points>
<connection>
<GID>1242</GID>
<name>OUT_0</name></connection>
<intersection>32 38</intersection>
<intersection>106 43</intersection>
<intersection>190 42</intersection>
<intersection>264 45</intersection>
<intersection>355 47</intersection>
<intersection>429 49</intersection>
<intersection>513 51</intersection>
<intersection>587 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32,-3537,32,-3524.5</points>
<connection>
<GID>1220</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190,-3537,190,-3526.5</points>
<connection>
<GID>1226</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106,-3537,106,-3524.5</points>
<connection>
<GID>1217</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264,-3537,264,-3526.5</points>
<connection>
<GID>1223</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355,-3537,355,-3528</points>
<connection>
<GID>1232</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429,-3537,429,-3528</points>
<connection>
<GID>1229</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513,-3537,513,-3530</points>
<connection>
<GID>1238</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587,-3537,587,-3530</points>
<connection>
<GID>1235</GID>
<name>IN_1</name></connection>
<intersection>-3537 33</intersection></vsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-3523.5,47.5,-3523.5</points>
<connection>
<GID>1220</GID>
<name>OUT</name></connection>
<connection>
<GID>1219</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-3532,29,-3515</points>
<intersection>-3532 3</intersection>
<intersection>-3522.5 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-3522.5,32,-3522.5</points>
<connection>
<GID>1220</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-3515,29,-3515</points>
<connection>
<GID>1218</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-3532,49.5,-3532</points>
<intersection>29 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-3532,49.5,-3526.5</points>
<connection>
<GID>1219</GID>
<name>IN_0</name></connection>
<intersection>-3532 3</intersection></vsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112,-3523.5,121,-3523.5</points>
<connection>
<GID>1217</GID>
<name>OUT</name></connection>
<connection>
<GID>1222</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-3533.5,102.5,-3515</points>
<intersection>-3533.5 3</intersection>
<intersection>-3522.5 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-3522.5,106,-3522.5</points>
<connection>
<GID>1217</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-3515,102.5,-3515</points>
<connection>
<GID>1221</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-3533.5,123,-3533.5</points>
<intersection>102.5 0</intersection>
<intersection>123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123,-3533.5,123,-3526.5</points>
<connection>
<GID>1222</GID>
<name>IN_0</name></connection>
<intersection>-3533.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>878</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,-3525.5,205.5,-3525.5</points>
<connection>
<GID>1226</GID>
<name>OUT</name></connection>
<connection>
<GID>1225</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-3534,187,-3515</points>
<intersection>-3534 3</intersection>
<intersection>-3524.5 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-3524.5,190,-3524.5</points>
<connection>
<GID>1226</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-3515,187,-3515</points>
<connection>
<GID>1224</GID>
<name>OUT_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,-3534,207.5,-3534</points>
<intersection>187 0</intersection>
<intersection>207.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207.5,-3534,207.5,-3528.5</points>
<connection>
<GID>1225</GID>
<name>IN_0</name></connection>
<intersection>-3534 3</intersection></vsegment></shape></wire>
<wire>
<ID>880</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270,-3525.5,279,-3525.5</points>
<connection>
<GID>1223</GID>
<name>OUT</name></connection>
<connection>
<GID>1228</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>881</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-3535.5,260.5,-3515</points>
<connection>
<GID>1227</GID>
<name>OUT_0</name></connection>
<intersection>-3535.5 3</intersection>
<intersection>-3524.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-3524.5,264,-3524.5</points>
<connection>
<GID>1223</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-3535.5,281,-3535.5</points>
<intersection>260.5 0</intersection>
<intersection>281 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281,-3535.5,281,-3528.5</points>
<connection>
<GID>1228</GID>
<name>IN_0</name></connection>
<intersection>-3535.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>882</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-3527,370.5,-3527</points>
<connection>
<GID>1232</GID>
<name>OUT</name></connection>
<connection>
<GID>1231</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>883</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-3535.5,352,-3515</points>
<intersection>-3535.5 3</intersection>
<intersection>-3526 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-3526,355,-3526</points>
<connection>
<GID>1232</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-3515,352,-3515</points>
<connection>
<GID>1230</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352,-3535.5,372.5,-3535.5</points>
<intersection>352 0</intersection>
<intersection>372.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372.5,-3535.5,372.5,-3530</points>
<connection>
<GID>1231</GID>
<name>IN_0</name></connection>
<intersection>-3535.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>884</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435,-3527,444,-3527</points>
<connection>
<GID>1229</GID>
<name>OUT</name></connection>
<connection>
<GID>1234</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>885</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-3535.5,425.5,-3515</points>
<intersection>-3535.5 3</intersection>
<intersection>-3526 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,-3526,429,-3526</points>
<connection>
<GID>1229</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,-3515,425.5,-3515</points>
<connection>
<GID>1233</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,-3535.5,446,-3535.5</points>
<intersection>425.5 0</intersection>
<intersection>446 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446,-3535.5,446,-3530</points>
<connection>
<GID>1234</GID>
<name>IN_0</name></connection>
<intersection>-3535.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>886</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-3529,528.5,-3529</points>
<connection>
<GID>1238</GID>
<name>OUT</name></connection>
<connection>
<GID>1237</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>887</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,-3535,510,-3515</points>
<intersection>-3535 3</intersection>
<intersection>-3528 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,-3528,513,-3528</points>
<connection>
<GID>1238</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509,-3515,510,-3515</points>
<connection>
<GID>1236</GID>
<name>OUT_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510,-3535,530.5,-3535</points>
<intersection>510 0</intersection>
<intersection>530.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530.5,-3535,530.5,-3532</points>
<connection>
<GID>1237</GID>
<name>IN_0</name></connection>
<intersection>-3535 3</intersection></vsegment></shape></wire>
<wire>
<ID>888</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593,-3529,602,-3529</points>
<connection>
<GID>1235</GID>
<name>OUT</name></connection>
<connection>
<GID>1240</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>889</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-3535,583.5,-3515</points>
<intersection>-3535 3</intersection>
<intersection>-3528 1</intersection>
<intersection>-3515 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,-3528,587,-3528</points>
<connection>
<GID>1235</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,-3515,583.5,-3515</points>
<connection>
<GID>1239</GID>
<name>OUT_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583.5,-3535,604,-3535</points>
<intersection>583.5 0</intersection>
<intersection>604 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604,-3535,604,-3532</points>
<connection>
<GID>1240</GID>
<name>IN_0</name></connection>
<intersection>-3535 3</intersection></vsegment></shape></wire>
<wire>
<ID>890</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,-3518,576.5,-3518</points>
<connection>
<GID>1241</GID>
<name>OUT</name></connection>
<connection>
<GID>1239</GID>
<name>clock</name></connection>
<connection>
<GID>1236</GID>
<name>clock</name></connection>
<connection>
<GID>1233</GID>
<name>clock</name></connection>
<connection>
<GID>1230</GID>
<name>clock</name></connection>
<connection>
<GID>1227</GID>
<name>clock</name></connection>
<connection>
<GID>1224</GID>
<name>clock</name></connection>
<connection>
<GID>1221</GID>
<name>clock</name></connection>
<connection>
<GID>1218</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-3793,-112,-3480</points>
<intersection>-3793 3</intersection>
<intersection>-3775 1</intersection>
<intersection>-3480 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112,-3775,-2.5,-3775</points>
<connection>
<GID>1267</GID>
<name>IN_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3480,-112,-3480</points>
<connection>
<GID>1295</GID>
<name>OUT_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112,-3793,-21,-3793</points>
<connection>
<GID>1268</GID>
<name>ENABLE_0</name></connection>
<intersection>-112 0</intersection></hsegment></shape></wire>
<wire>
<ID>892</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-18.5,-3795,594,-3795</points>
<connection>
<GID>1268</GID>
<name>OUT_0</name></connection>
<intersection>39 38</intersection>
<intersection>113 43</intersection>
<intersection>197 42</intersection>
<intersection>271 45</intersection>
<intersection>362 47</intersection>
<intersection>436 49</intersection>
<intersection>520 51</intersection>
<intersection>594 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>39,-3795,39,-3782.5</points>
<connection>
<GID>1246</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>197,-3795,197,-3784.5</points>
<connection>
<GID>1252</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>113,-3795,113,-3782.5</points>
<connection>
<GID>1243</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>271,-3795,271,-3784.5</points>
<connection>
<GID>1249</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>362,-3795,362,-3786</points>
<connection>
<GID>1258</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>436,-3795,436,-3786</points>
<connection>
<GID>1255</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>520,-3795,520,-3788</points>
<connection>
<GID>1264</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>594,-3795,594,-3788</points>
<connection>
<GID>1261</GID>
<name>IN_1</name></connection>
<intersection>-3795 33</intersection></vsegment></shape></wire>
<wire>
<ID>893</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-3781.5,54.5,-3781.5</points>
<connection>
<GID>1246</GID>
<name>OUT</name></connection>
<connection>
<GID>1245</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>894</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-3790,36,-3773</points>
<intersection>-3790 3</intersection>
<intersection>-3780.5 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-3780.5,39,-3780.5</points>
<connection>
<GID>1246</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-3773,36,-3773</points>
<connection>
<GID>1244</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-3790,56.5,-3790</points>
<intersection>36 0</intersection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56.5,-3790,56.5,-3784.5</points>
<connection>
<GID>1245</GID>
<name>IN_0</name></connection>
<intersection>-3790 3</intersection></vsegment></shape></wire>
<wire>
<ID>895</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,-3781.5,128,-3781.5</points>
<connection>
<GID>1243</GID>
<name>OUT</name></connection>
<connection>
<GID>1248</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>896</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-3791.5,109.5,-3773</points>
<intersection>-3791.5 3</intersection>
<intersection>-3780.5 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-3780.5,113,-3780.5</points>
<connection>
<GID>1243</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-3773,109.5,-3773</points>
<connection>
<GID>1247</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-3791.5,130,-3791.5</points>
<intersection>109.5 0</intersection>
<intersection>130 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130,-3791.5,130,-3784.5</points>
<connection>
<GID>1248</GID>
<name>IN_0</name></connection>
<intersection>-3791.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>897</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,-3783.5,212.5,-3783.5</points>
<connection>
<GID>1252</GID>
<name>OUT</name></connection>
<connection>
<GID>1251</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>898</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-3792,194,-3773</points>
<intersection>-3792 3</intersection>
<intersection>-3782.5 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,-3782.5,197,-3782.5</points>
<connection>
<GID>1252</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>193,-3773,194,-3773</points>
<connection>
<GID>1250</GID>
<name>OUT_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>194,-3792,214.5,-3792</points>
<intersection>194 0</intersection>
<intersection>214.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>214.5,-3792,214.5,-3786.5</points>
<connection>
<GID>1251</GID>
<name>IN_0</name></connection>
<intersection>-3792 3</intersection></vsegment></shape></wire>
<wire>
<ID>899</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>277,-3783.5,286,-3783.5</points>
<connection>
<GID>1249</GID>
<name>OUT</name></connection>
<connection>
<GID>1254</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>900</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-3793.5,267.5,-3773</points>
<connection>
<GID>1253</GID>
<name>OUT_0</name></connection>
<intersection>-3793.5 3</intersection>
<intersection>-3782.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-3782.5,271,-3782.5</points>
<connection>
<GID>1249</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>267.5,-3793.5,288,-3793.5</points>
<intersection>267.5 0</intersection>
<intersection>288 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>288,-3793.5,288,-3786.5</points>
<connection>
<GID>1254</GID>
<name>IN_0</name></connection>
<intersection>-3793.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>901</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-3785,377.5,-3785</points>
<connection>
<GID>1258</GID>
<name>OUT</name></connection>
<connection>
<GID>1257</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>902</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-3793.5,359,-3773</points>
<intersection>-3793.5 3</intersection>
<intersection>-3784 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-3784,362,-3784</points>
<connection>
<GID>1258</GID>
<name>IN_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>358,-3773,359,-3773</points>
<connection>
<GID>1256</GID>
<name>OUT_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>359,-3793.5,379.5,-3793.5</points>
<intersection>359 0</intersection>
<intersection>379.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>379.5,-3793.5,379.5,-3788</points>
<connection>
<GID>1257</GID>
<name>IN_0</name></connection>
<intersection>-3793.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>903</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>442,-3785,451,-3785</points>
<connection>
<GID>1255</GID>
<name>OUT</name></connection>
<connection>
<GID>1260</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>904</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,-3793.5,432.5,-3773</points>
<intersection>-3793.5 3</intersection>
<intersection>-3784 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,-3784,436,-3784</points>
<connection>
<GID>1255</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-3773,432.5,-3773</points>
<connection>
<GID>1259</GID>
<name>OUT_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432.5,-3793.5,453,-3793.5</points>
<intersection>432.5 0</intersection>
<intersection>453 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>453,-3793.5,453,-3788</points>
<connection>
<GID>1260</GID>
<name>IN_0</name></connection>
<intersection>-3793.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>905</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>526,-3787,535.5,-3787</points>
<connection>
<GID>1264</GID>
<name>OUT</name></connection>
<connection>
<GID>1263</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>906</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,-3793,517,-3773</points>
<intersection>-3793 3</intersection>
<intersection>-3786 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,-3786,520,-3786</points>
<connection>
<GID>1264</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>516,-3773,517,-3773</points>
<connection>
<GID>1262</GID>
<name>OUT_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>517,-3793,537.5,-3793</points>
<intersection>517 0</intersection>
<intersection>537.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>537.5,-3793,537.5,-3790</points>
<connection>
<GID>1263</GID>
<name>IN_0</name></connection>
<intersection>-3793 3</intersection></vsegment></shape></wire>
<wire>
<ID>907</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>600,-3787,609,-3787</points>
<connection>
<GID>1261</GID>
<name>OUT</name></connection>
<connection>
<GID>1266</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,-3793,590.5,-3773</points>
<intersection>-3793 3</intersection>
<intersection>-3786 1</intersection>
<intersection>-3773 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,-3786,594,-3786</points>
<connection>
<GID>1261</GID>
<name>IN_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,-3773,590.5,-3773</points>
<connection>
<GID>1265</GID>
<name>OUT_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>590.5,-3793,611,-3793</points>
<intersection>590.5 0</intersection>
<intersection>611 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>611,-3793,611,-3790</points>
<connection>
<GID>1266</GID>
<name>IN_0</name></connection>
<intersection>-3793 3</intersection></vsegment></shape></wire>
<wire>
<ID>909</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-3776,583.5,-3776</points>
<connection>
<GID>1267</GID>
<name>OUT</name></connection>
<connection>
<GID>1265</GID>
<name>clock</name></connection>
<connection>
<GID>1262</GID>
<name>clock</name></connection>
<connection>
<GID>1259</GID>
<name>clock</name></connection>
<connection>
<GID>1256</GID>
<name>clock</name></connection>
<connection>
<GID>1253</GID>
<name>clock</name></connection>
<connection>
<GID>1250</GID>
<name>clock</name></connection>
<connection>
<GID>1247</GID>
<name>clock</name></connection>
<connection>
<GID>1244</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-3703,-110,-3479</points>
<intersection>-3703 3</intersection>
<intersection>-3685 1</intersection>
<intersection>-3479 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-3685,-5.5,-3685</points>
<connection>
<GID>1293</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-3479,-110,-3479</points>
<connection>
<GID>1295</GID>
<name>OUT_1</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-3703,-24,-3703</points>
<connection>
<GID>1294</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>911</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21.5,-3705,591,-3705</points>
<connection>
<GID>1294</GID>
<name>OUT_0</name></connection>
<intersection>36 38</intersection>
<intersection>110 43</intersection>
<intersection>194 42</intersection>
<intersection>268 45</intersection>
<intersection>359 47</intersection>
<intersection>433 49</intersection>
<intersection>517 51</intersection>
<intersection>591 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36,-3705,36,-3692.5</points>
<connection>
<GID>1272</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194,-3705,194,-3694.5</points>
<connection>
<GID>1278</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110,-3705,110,-3692.5</points>
<connection>
<GID>1269</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268,-3705,268,-3694.5</points>
<connection>
<GID>1275</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359,-3705,359,-3696</points>
<connection>
<GID>1284</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433,-3705,433,-3696</points>
<connection>
<GID>1281</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517,-3705,517,-3698</points>
<connection>
<GID>1290</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591,-3705,591,-3698</points>
<connection>
<GID>1287</GID>
<name>IN_1</name></connection>
<intersection>-3705 33</intersection></vsegment></shape></wire>
<wire>
<ID>912</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-3691.5,51.5,-3691.5</points>
<connection>
<GID>1272</GID>
<name>OUT</name></connection>
<connection>
<GID>1271</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>913</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-3700,33,-3683</points>
<intersection>-3700 3</intersection>
<intersection>-3690.5 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-3690.5,36,-3690.5</points>
<connection>
<GID>1272</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-3683,33,-3683</points>
<connection>
<GID>1270</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-3700,53.5,-3700</points>
<intersection>33 0</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-3700,53.5,-3694.5</points>
<connection>
<GID>1271</GID>
<name>IN_0</name></connection>
<intersection>-3700 3</intersection></vsegment></shape></wire>
<wire>
<ID>914</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116,-3691.5,125,-3691.5</points>
<connection>
<GID>1269</GID>
<name>OUT</name></connection>
<connection>
<GID>1274</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-3701.5,106.5,-3683</points>
<intersection>-3701.5 3</intersection>
<intersection>-3690.5 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-3690.5,110,-3690.5</points>
<connection>
<GID>1269</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-3683,106.5,-3683</points>
<connection>
<GID>1273</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,-3701.5,127,-3701.5</points>
<intersection>106.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-3701.5,127,-3694.5</points>
<connection>
<GID>1274</GID>
<name>IN_0</name></connection>
<intersection>-3701.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-3693.5,209.5,-3693.5</points>
<connection>
<GID>1278</GID>
<name>OUT</name></connection>
<connection>
<GID>1277</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-3702,191,-3683</points>
<intersection>-3702 3</intersection>
<intersection>-3692.5 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-3692.5,194,-3692.5</points>
<connection>
<GID>1278</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,-3683,191,-3683</points>
<connection>
<GID>1276</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191,-3702,211.5,-3702</points>
<intersection>191 0</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211.5,-3702,211.5,-3696.5</points>
<connection>
<GID>1277</GID>
<name>IN_0</name></connection>
<intersection>-3702 3</intersection></vsegment></shape></wire>
<wire>
<ID>918</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274,-3693.5,283,-3693.5</points>
<connection>
<GID>1275</GID>
<name>OUT</name></connection>
<connection>
<GID>1280</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-3703.5,264.5,-3683</points>
<connection>
<GID>1279</GID>
<name>OUT_0</name></connection>
<intersection>-3703.5 3</intersection>
<intersection>-3692.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-3692.5,268,-3692.5</points>
<connection>
<GID>1275</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264.5,-3703.5,285,-3703.5</points>
<intersection>264.5 0</intersection>
<intersection>285 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285,-3703.5,285,-3696.5</points>
<connection>
<GID>1280</GID>
<name>IN_0</name></connection>
<intersection>-3703.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>920</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365,-3695,374.5,-3695</points>
<connection>
<GID>1284</GID>
<name>OUT</name></connection>
<connection>
<GID>1283</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-3703.5,356,-3683</points>
<intersection>-3703.5 3</intersection>
<intersection>-3694 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-3694,359,-3694</points>
<connection>
<GID>1284</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355,-3683,356,-3683</points>
<connection>
<GID>1282</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356,-3703.5,376.5,-3703.5</points>
<intersection>356 0</intersection>
<intersection>376.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376.5,-3703.5,376.5,-3698</points>
<connection>
<GID>1283</GID>
<name>IN_0</name></connection>
<intersection>-3703.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>922</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439,-3695,448,-3695</points>
<connection>
<GID>1281</GID>
<name>OUT</name></connection>
<connection>
<GID>1286</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>923</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-3703.5,429.5,-3683</points>
<intersection>-3703.5 3</intersection>
<intersection>-3694 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,-3694,433,-3694</points>
<connection>
<GID>1281</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,-3683,429.5,-3683</points>
<connection>
<GID>1285</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,-3703.5,450,-3703.5</points>
<intersection>429.5 0</intersection>
<intersection>450 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450,-3703.5,450,-3698</points>
<connection>
<GID>1286</GID>
<name>IN_0</name></connection>
<intersection>-3703.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>924</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523,-3697,532.5,-3697</points>
<connection>
<GID>1290</GID>
<name>OUT</name></connection>
<connection>
<GID>1289</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>925</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-3703,514,-3683</points>
<intersection>-3703 3</intersection>
<intersection>-3696 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-3696,517,-3696</points>
<connection>
<GID>1290</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,-3683,514,-3683</points>
<connection>
<GID>1288</GID>
<name>OUT_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514,-3703,534.5,-3703</points>
<intersection>514 0</intersection>
<intersection>534.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534.5,-3703,534.5,-3700</points>
<connection>
<GID>1289</GID>
<name>IN_0</name></connection>
<intersection>-3703 3</intersection></vsegment></shape></wire>
<wire>
<ID>926</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597,-3697,606,-3697</points>
<connection>
<GID>1287</GID>
<name>OUT</name></connection>
<connection>
<GID>1292</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>927</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,-3703,587.5,-3683</points>
<intersection>-3703 3</intersection>
<intersection>-3696 1</intersection>
<intersection>-3683 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,-3696,591,-3696</points>
<connection>
<GID>1287</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586.5,-3683,587.5,-3683</points>
<connection>
<GID>1291</GID>
<name>OUT_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587.5,-3703,608,-3703</points>
<intersection>587.5 0</intersection>
<intersection>608 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608,-3703,608,-3700</points>
<connection>
<GID>1292</GID>
<name>IN_0</name></connection>
<intersection>-3703 3</intersection></vsegment></shape></wire>
<wire>
<ID>928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-3686,580.5,-3686</points>
<connection>
<GID>1270</GID>
<name>clock</name></connection>
<connection>
<GID>1273</GID>
<name>clock</name></connection>
<connection>
<GID>1279</GID>
<name>clock</name></connection>
<connection>
<GID>1282</GID>
<name>clock</name></connection>
<connection>
<GID>1285</GID>
<name>clock</name></connection>
<connection>
<GID>1288</GID>
<name>clock</name></connection>
<connection>
<GID>1291</GID>
<name>clock</name></connection>
<connection>
<GID>1293</GID>
<name>OUT</name></connection>
<connection>
<GID>1276</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>929</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-4299.5,-110,-4056.5</points>
<intersection>-4299.5 2</intersection>
<intersection>-4074.5 3</intersection>
<intersection>-4056.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-4056.5,-8.5,-4056.5</points>
<connection>
<GID>1390</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4299.5,-110,-4299.5</points>
<connection>
<GID>1365</GID>
<name>OUT_6</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-4074.5,-27,-4074.5</points>
<connection>
<GID>1391</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>930</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-24.5,-4076.5,588,-4076.5</points>
<connection>
<GID>1391</GID>
<name>OUT_0</name></connection>
<intersection>33 38</intersection>
<intersection>107 43</intersection>
<intersection>191 42</intersection>
<intersection>265 45</intersection>
<intersection>356 47</intersection>
<intersection>430 49</intersection>
<intersection>514 51</intersection>
<intersection>588 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>33,-4076.5,33,-4064</points>
<connection>
<GID>1369</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>191,-4076.5,191,-4066</points>
<connection>
<GID>1375</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>107,-4076.5,107,-4064</points>
<connection>
<GID>1366</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>265,-4076.5,265,-4066</points>
<connection>
<GID>1372</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>356,-4076.5,356,-4067.5</points>
<connection>
<GID>1381</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>430,-4076.5,430,-4067.5</points>
<connection>
<GID>1378</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>514,-4076.5,514,-4069.5</points>
<connection>
<GID>1387</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>588,-4076.5,588,-4069.5</points>
<connection>
<GID>1384</GID>
<name>IN_1</name></connection>
<intersection>-4076.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>931</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-4063,48.5,-4063</points>
<connection>
<GID>1369</GID>
<name>OUT</name></connection>
<connection>
<GID>1368</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-4071.5,30,-4054.5</points>
<intersection>-4071.5 3</intersection>
<intersection>-4062 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-4062,33,-4062</points>
<connection>
<GID>1369</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-4054.5,30,-4054.5</points>
<connection>
<GID>1367</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30,-4071.5,50.5,-4071.5</points>
<intersection>30 0</intersection>
<intersection>50.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50.5,-4071.5,50.5,-4066</points>
<connection>
<GID>1368</GID>
<name>IN_0</name></connection>
<intersection>-4071.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113,-4063,122,-4063</points>
<connection>
<GID>1366</GID>
<name>OUT</name></connection>
<connection>
<GID>1371</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-4073,103.5,-4054.5</points>
<intersection>-4073 3</intersection>
<intersection>-4062 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-4062,107,-4062</points>
<connection>
<GID>1366</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-4054.5,103.5,-4054.5</points>
<connection>
<GID>1370</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,-4073,124,-4073</points>
<intersection>103.5 0</intersection>
<intersection>124 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124,-4073,124,-4066</points>
<connection>
<GID>1371</GID>
<name>IN_0</name></connection>
<intersection>-4073 3</intersection></vsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-4065,206.5,-4065</points>
<connection>
<GID>1375</GID>
<name>OUT</name></connection>
<connection>
<GID>1374</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-4073.5,188,-4054.5</points>
<intersection>-4073.5 3</intersection>
<intersection>-4064 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188,-4064,191,-4064</points>
<connection>
<GID>1375</GID>
<name>IN_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-4054.5,188,-4054.5</points>
<connection>
<GID>1373</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188,-4073.5,208.5,-4073.5</points>
<intersection>188 0</intersection>
<intersection>208.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208.5,-4073.5,208.5,-4068</points>
<connection>
<GID>1374</GID>
<name>IN_0</name></connection>
<intersection>-4073.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>271,-4065,280,-4065</points>
<connection>
<GID>1372</GID>
<name>OUT</name></connection>
<connection>
<GID>1377</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-4075,261.5,-4054.5</points>
<connection>
<GID>1376</GID>
<name>OUT_0</name></connection>
<intersection>-4075 3</intersection>
<intersection>-4064 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-4064,265,-4064</points>
<connection>
<GID>1372</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-4075,282,-4075</points>
<intersection>261.5 0</intersection>
<intersection>282 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282,-4075,282,-4068</points>
<connection>
<GID>1377</GID>
<name>IN_0</name></connection>
<intersection>-4075 3</intersection></vsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362,-4066.5,371.5,-4066.5</points>
<connection>
<GID>1381</GID>
<name>OUT</name></connection>
<connection>
<GID>1380</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-4075,353,-4054.5</points>
<intersection>-4075 3</intersection>
<intersection>-4065.5 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-4065.5,356,-4065.5</points>
<connection>
<GID>1381</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-4054.5,353,-4054.5</points>
<connection>
<GID>1379</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353,-4075,373.5,-4075</points>
<intersection>353 0</intersection>
<intersection>373.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>373.5,-4075,373.5,-4069.5</points>
<connection>
<GID>1380</GID>
<name>IN_0</name></connection>
<intersection>-4075 3</intersection></vsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>436,-4066.5,445,-4066.5</points>
<connection>
<GID>1378</GID>
<name>OUT</name></connection>
<connection>
<GID>1383</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-4075,426.5,-4054.5</points>
<intersection>-4075 3</intersection>
<intersection>-4065.5 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426.5,-4065.5,430,-4065.5</points>
<connection>
<GID>1378</GID>
<name>IN_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425.5,-4054.5,426.5,-4054.5</points>
<connection>
<GID>1382</GID>
<name>OUT_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426.5,-4075,447,-4075</points>
<intersection>426.5 0</intersection>
<intersection>447 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447,-4075,447,-4069.5</points>
<connection>
<GID>1383</GID>
<name>IN_0</name></connection>
<intersection>-4075 3</intersection></vsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520,-4068.5,529.5,-4068.5</points>
<connection>
<GID>1387</GID>
<name>OUT</name></connection>
<connection>
<GID>1386</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,-4074.5,511,-4054.5</points>
<intersection>-4074.5 3</intersection>
<intersection>-4067.5 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,-4067.5,514,-4067.5</points>
<connection>
<GID>1387</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>510,-4054.5,511,-4054.5</points>
<connection>
<GID>1385</GID>
<name>OUT_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511,-4074.5,531.5,-4074.5</points>
<intersection>511 0</intersection>
<intersection>531.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531.5,-4074.5,531.5,-4071.5</points>
<connection>
<GID>1386</GID>
<name>IN_0</name></connection>
<intersection>-4074.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>594,-4068.5,603,-4068.5</points>
<connection>
<GID>1384</GID>
<name>OUT</name></connection>
<connection>
<GID>1389</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,-4074.5,584.5,-4054.5</points>
<intersection>-4074.5 3</intersection>
<intersection>-4067.5 1</intersection>
<intersection>-4054.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584.5,-4067.5,588,-4067.5</points>
<connection>
<GID>1384</GID>
<name>IN_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583.5,-4054.5,584.5,-4054.5</points>
<connection>
<GID>1388</GID>
<name>OUT_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>584.5,-4074.5,605,-4074.5</points>
<intersection>584.5 0</intersection>
<intersection>605 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>605,-4074.5,605,-4071.5</points>
<connection>
<GID>1389</GID>
<name>IN_0</name></connection>
<intersection>-4074.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>947</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-4057.5,577.5,-4057.5</points>
<connection>
<GID>1390</GID>
<name>OUT</name></connection>
<connection>
<GID>1388</GID>
<name>clock</name></connection>
<connection>
<GID>1385</GID>
<name>clock</name></connection>
<connection>
<GID>1382</GID>
<name>clock</name></connection>
<connection>
<GID>1379</GID>
<name>clock</name></connection>
<connection>
<GID>1376</GID>
<name>clock</name></connection>
<connection>
<GID>1373</GID>
<name>clock</name></connection>
<connection>
<GID>1370</GID>
<name>clock</name></connection>
<connection>
<GID>1367</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-4298.5,-111,-3966.5</points>
<intersection>-4298.5 2</intersection>
<intersection>-3984.5 3</intersection>
<intersection>-3966.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-3966.5,-11.5,-3966.5</points>
<connection>
<GID>1416</GID>
<name>IN_0</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4298.5,-111,-4298.5</points>
<connection>
<GID>1365</GID>
<name>OUT_7</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111,-3984.5,-30,-3984.5</points>
<connection>
<GID>1417</GID>
<name>ENABLE_0</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-27.5,-3986.5,585,-3986.5</points>
<connection>
<GID>1417</GID>
<name>OUT_0</name></connection>
<intersection>30 38</intersection>
<intersection>104 43</intersection>
<intersection>188 42</intersection>
<intersection>262 45</intersection>
<intersection>353 47</intersection>
<intersection>427 49</intersection>
<intersection>511 51</intersection>
<intersection>585 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>30,-3986.5,30,-3974</points>
<connection>
<GID>1395</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>188,-3986.5,188,-3976</points>
<connection>
<GID>1401</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>104,-3986.5,104,-3974</points>
<connection>
<GID>1392</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>262,-3986.5,262,-3976</points>
<connection>
<GID>1398</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>353,-3986.5,353,-3977.5</points>
<connection>
<GID>1407</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>427,-3986.5,427,-3977.5</points>
<connection>
<GID>1404</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>511,-3986.5,511,-3979.5</points>
<connection>
<GID>1413</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>585,-3986.5,585,-3979.5</points>
<connection>
<GID>1410</GID>
<name>IN_1</name></connection>
<intersection>-3986.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-3973,45.5,-3973</points>
<connection>
<GID>1395</GID>
<name>OUT</name></connection>
<connection>
<GID>1394</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-3981.5,27,-3964.5</points>
<intersection>-3981.5 3</intersection>
<intersection>-3972 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-3972,30,-3972</points>
<connection>
<GID>1395</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-3964.5,27,-3964.5</points>
<connection>
<GID>1393</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-3981.5,47.5,-3981.5</points>
<intersection>27 0</intersection>
<intersection>47.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-3981.5,47.5,-3976</points>
<connection>
<GID>1394</GID>
<name>IN_0</name></connection>
<intersection>-3981.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>110,-3973,119,-3973</points>
<connection>
<GID>1392</GID>
<name>OUT</name></connection>
<connection>
<GID>1397</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-3983,100.5,-3964.5</points>
<intersection>-3983 3</intersection>
<intersection>-3972 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-3972,104,-3972</points>
<connection>
<GID>1392</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-3964.5,100.5,-3964.5</points>
<connection>
<GID>1396</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100.5,-3983,121,-3983</points>
<intersection>100.5 0</intersection>
<intersection>121 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>121,-3983,121,-3976</points>
<connection>
<GID>1397</GID>
<name>IN_0</name></connection>
<intersection>-3983 3</intersection></vsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,-3975,203.5,-3975</points>
<connection>
<GID>1401</GID>
<name>OUT</name></connection>
<connection>
<GID>1400</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-3983.5,185,-3964.5</points>
<intersection>-3983.5 3</intersection>
<intersection>-3974 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-3974,188,-3974</points>
<connection>
<GID>1401</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-3964.5,185,-3964.5</points>
<connection>
<GID>1399</GID>
<name>OUT_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185,-3983.5,205.5,-3983.5</points>
<intersection>185 0</intersection>
<intersection>205.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>205.5,-3983.5,205.5,-3978</points>
<connection>
<GID>1400</GID>
<name>IN_0</name></connection>
<intersection>-3983.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>268,-3975,277,-3975</points>
<connection>
<GID>1398</GID>
<name>OUT</name></connection>
<connection>
<GID>1403</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-3985,258.5,-3964.5</points>
<connection>
<GID>1402</GID>
<name>OUT_0</name></connection>
<intersection>-3985 3</intersection>
<intersection>-3974 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,-3974,262,-3974</points>
<connection>
<GID>1398</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,-3985,279,-3985</points>
<intersection>258.5 0</intersection>
<intersection>279 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>279,-3985,279,-3978</points>
<connection>
<GID>1403</GID>
<name>IN_0</name></connection>
<intersection>-3985 3</intersection></vsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-3976.5,368.5,-3976.5</points>
<connection>
<GID>1407</GID>
<name>OUT</name></connection>
<connection>
<GID>1406</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-3985,350,-3964.5</points>
<intersection>-3985 3</intersection>
<intersection>-3975.5 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-3975.5,353,-3975.5</points>
<connection>
<GID>1407</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-3964.5,350,-3964.5</points>
<connection>
<GID>1405</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>350,-3985,370.5,-3985</points>
<intersection>350 0</intersection>
<intersection>370.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>370.5,-3985,370.5,-3979.5</points>
<connection>
<GID>1406</GID>
<name>IN_0</name></connection>
<intersection>-3985 3</intersection></vsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>433,-3976.5,442,-3976.5</points>
<connection>
<GID>1404</GID>
<name>OUT</name></connection>
<connection>
<GID>1409</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-3985,423.5,-3964.5</points>
<intersection>-3985 3</intersection>
<intersection>-3975.5 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423.5,-3975.5,427,-3975.5</points>
<connection>
<GID>1404</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422.5,-3964.5,423.5,-3964.5</points>
<connection>
<GID>1408</GID>
<name>OUT_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>423.5,-3985,444,-3985</points>
<intersection>423.5 0</intersection>
<intersection>444 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>444,-3985,444,-3979.5</points>
<connection>
<GID>1409</GID>
<name>IN_0</name></connection>
<intersection>-3985 3</intersection></vsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>517,-3978.5,526.5,-3978.5</points>
<connection>
<GID>1413</GID>
<name>OUT</name></connection>
<connection>
<GID>1412</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508,-3984.5,508,-3964.5</points>
<intersection>-3984.5 3</intersection>
<intersection>-3977.5 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,-3977.5,511,-3977.5</points>
<connection>
<GID>1413</GID>
<name>IN_0</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507,-3964.5,508,-3964.5</points>
<connection>
<GID>1411</GID>
<name>OUT_0</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>508,-3984.5,528.5,-3984.5</points>
<intersection>508 0</intersection>
<intersection>528.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>528.5,-3984.5,528.5,-3981.5</points>
<connection>
<GID>1412</GID>
<name>IN_0</name></connection>
<intersection>-3984.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>591,-3978.5,600,-3978.5</points>
<connection>
<GID>1410</GID>
<name>OUT</name></connection>
<connection>
<GID>1415</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>965</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581.5,-3984.5,581.5,-3964.5</points>
<intersection>-3984.5 3</intersection>
<intersection>-3977.5 1</intersection>
<intersection>-3964.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581.5,-3977.5,585,-3977.5</points>
<connection>
<GID>1410</GID>
<name>IN_0</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>580.5,-3964.5,581.5,-3964.5</points>
<connection>
<GID>1414</GID>
<name>OUT_0</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>581.5,-3984.5,602,-3984.5</points>
<intersection>581.5 0</intersection>
<intersection>602 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>602,-3984.5,602,-3981.5</points>
<connection>
<GID>1415</GID>
<name>IN_0</name></connection>
<intersection>-3984.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-3967.5,574.5,-3967.5</points>
<connection>
<GID>1416</GID>
<name>OUT</name></connection>
<connection>
<GID>1414</GID>
<name>clock</name></connection>
<connection>
<GID>1411</GID>
<name>clock</name></connection>
<connection>
<GID>1408</GID>
<name>clock</name></connection>
<connection>
<GID>1405</GID>
<name>clock</name></connection>
<connection>
<GID>1402</GID>
<name>clock</name></connection>
<connection>
<GID>1399</GID>
<name>clock</name></connection>
<connection>
<GID>1396</GID>
<name>clock</name></connection>
<connection>
<GID>1393</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-4301.5,-108,-4224.5</points>
<intersection>-4301.5 2</intersection>
<intersection>-4242.5 3</intersection>
<intersection>-4224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-4224.5,-4.5,-4224.5</points>
<connection>
<GID>1442</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4301.5,-108,-4301.5</points>
<connection>
<GID>1365</GID>
<name>OUT_4</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-4242.5,-23,-4242.5</points>
<connection>
<GID>1443</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-20.5,-4244.5,592,-4244.5</points>
<connection>
<GID>1443</GID>
<name>OUT_0</name></connection>
<intersection>37 38</intersection>
<intersection>111 43</intersection>
<intersection>195 42</intersection>
<intersection>269 45</intersection>
<intersection>360 47</intersection>
<intersection>434 49</intersection>
<intersection>518 51</intersection>
<intersection>592 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>37,-4244.5,37,-4232</points>
<connection>
<GID>1421</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>195,-4244.5,195,-4234</points>
<connection>
<GID>1427</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>111,-4244.5,111,-4232</points>
<connection>
<GID>1418</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>269,-4244.5,269,-4234</points>
<connection>
<GID>1424</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>360,-4244.5,360,-4235.5</points>
<connection>
<GID>1433</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>434,-4244.5,434,-4235.5</points>
<connection>
<GID>1430</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>518,-4244.5,518,-4237.5</points>
<connection>
<GID>1439</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>592,-4244.5,592,-4237.5</points>
<connection>
<GID>1436</GID>
<name>IN_1</name></connection>
<intersection>-4244.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-4231,52.5,-4231</points>
<connection>
<GID>1421</GID>
<name>OUT</name></connection>
<connection>
<GID>1420</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-4239.5,34,-4222.5</points>
<intersection>-4239.5 3</intersection>
<intersection>-4230 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-4230,37,-4230</points>
<connection>
<GID>1421</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-4222.5,34,-4222.5</points>
<connection>
<GID>1419</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-4239.5,54.5,-4239.5</points>
<intersection>34 0</intersection>
<intersection>54.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54.5,-4239.5,54.5,-4234</points>
<connection>
<GID>1420</GID>
<name>IN_0</name></connection>
<intersection>-4239.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>117,-4231,126,-4231</points>
<connection>
<GID>1418</GID>
<name>OUT</name></connection>
<connection>
<GID>1423</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-4241,107.5,-4222.5</points>
<intersection>-4241 3</intersection>
<intersection>-4230 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-4230,111,-4230</points>
<connection>
<GID>1418</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-4222.5,107.5,-4222.5</points>
<connection>
<GID>1422</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-4241,128,-4241</points>
<intersection>107.5 0</intersection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-4241,128,-4234</points>
<connection>
<GID>1423</GID>
<name>IN_0</name></connection>
<intersection>-4241 3</intersection></vsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201,-4233,210.5,-4233</points>
<connection>
<GID>1427</GID>
<name>OUT</name></connection>
<connection>
<GID>1426</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-4241.5,192,-4222.5</points>
<intersection>-4241.5 3</intersection>
<intersection>-4232 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-4232,195,-4232</points>
<connection>
<GID>1427</GID>
<name>IN_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-4222.5,192,-4222.5</points>
<connection>
<GID>1425</GID>
<name>OUT_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>192,-4241.5,212.5,-4241.5</points>
<intersection>192 0</intersection>
<intersection>212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>212.5,-4241.5,212.5,-4236</points>
<connection>
<GID>1426</GID>
<name>IN_0</name></connection>
<intersection>-4241.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>275,-4233,284,-4233</points>
<connection>
<GID>1424</GID>
<name>OUT</name></connection>
<connection>
<GID>1429</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-4243,265.5,-4222.5</points>
<connection>
<GID>1428</GID>
<name>OUT_0</name></connection>
<intersection>-4243 3</intersection>
<intersection>-4232 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265.5,-4232,269,-4232</points>
<connection>
<GID>1424</GID>
<name>IN_0</name></connection>
<intersection>265.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>265.5,-4243,286,-4243</points>
<intersection>265.5 0</intersection>
<intersection>286 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>286,-4243,286,-4236</points>
<connection>
<GID>1429</GID>
<name>IN_0</name></connection>
<intersection>-4243 3</intersection></vsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366,-4234.5,375.5,-4234.5</points>
<connection>
<GID>1433</GID>
<name>OUT</name></connection>
<connection>
<GID>1432</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-4243,357,-4222.5</points>
<intersection>-4243 3</intersection>
<intersection>-4233.5 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-4233.5,360,-4233.5</points>
<connection>
<GID>1433</GID>
<name>IN_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356,-4222.5,357,-4222.5</points>
<connection>
<GID>1431</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-4243,377.5,-4243</points>
<intersection>357 0</intersection>
<intersection>377.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>377.5,-4243,377.5,-4237.5</points>
<connection>
<GID>1432</GID>
<name>IN_0</name></connection>
<intersection>-4243 3</intersection></vsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>440,-4234.5,449,-4234.5</points>
<connection>
<GID>1430</GID>
<name>OUT</name></connection>
<connection>
<GID>1435</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,-4243,430.5,-4222.5</points>
<intersection>-4243 3</intersection>
<intersection>-4233.5 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430.5,-4233.5,434,-4233.5</points>
<connection>
<GID>1430</GID>
<name>IN_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>429.5,-4222.5,430.5,-4222.5</points>
<connection>
<GID>1434</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>430.5,-4243,451,-4243</points>
<intersection>430.5 0</intersection>
<intersection>451 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>451,-4243,451,-4237.5</points>
<connection>
<GID>1435</GID>
<name>IN_0</name></connection>
<intersection>-4243 3</intersection></vsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>524,-4236.5,533.5,-4236.5</points>
<connection>
<GID>1439</GID>
<name>OUT</name></connection>
<connection>
<GID>1438</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-4242.5,515,-4222.5</points>
<intersection>-4242.5 3</intersection>
<intersection>-4235.5 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515,-4235.5,518,-4235.5</points>
<connection>
<GID>1439</GID>
<name>IN_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,-4222.5,515,-4222.5</points>
<connection>
<GID>1437</GID>
<name>OUT_0</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>515,-4242.5,535.5,-4242.5</points>
<intersection>515 0</intersection>
<intersection>535.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535.5,-4242.5,535.5,-4239.5</points>
<connection>
<GID>1438</GID>
<name>IN_0</name></connection>
<intersection>-4242.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>598,-4236.5,607,-4236.5</points>
<connection>
<GID>1436</GID>
<name>OUT</name></connection>
<connection>
<GID>1441</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588.5,-4242.5,588.5,-4222.5</points>
<intersection>-4242.5 3</intersection>
<intersection>-4235.5 1</intersection>
<intersection>-4222.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588.5,-4235.5,592,-4235.5</points>
<connection>
<GID>1436</GID>
<name>IN_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-4222.5,588.5,-4222.5</points>
<connection>
<GID>1440</GID>
<name>OUT_0</name></connection>
<intersection>588.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>588.5,-4242.5,609,-4242.5</points>
<intersection>588.5 0</intersection>
<intersection>609 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>609,-4242.5,609,-4239.5</points>
<connection>
<GID>1441</GID>
<name>IN_0</name></connection>
<intersection>-4242.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-4225.5,581.5,-4225.5</points>
<connection>
<GID>1442</GID>
<name>OUT</name></connection>
<connection>
<GID>1440</GID>
<name>clock</name></connection>
<connection>
<GID>1437</GID>
<name>clock</name></connection>
<connection>
<GID>1434</GID>
<name>clock</name></connection>
<connection>
<GID>1431</GID>
<name>clock</name></connection>
<connection>
<GID>1428</GID>
<name>clock</name></connection>
<connection>
<GID>1425</GID>
<name>clock</name></connection>
<connection>
<GID>1422</GID>
<name>clock</name></connection>
<connection>
<GID>1419</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-4300.5,-109,-4134.5</points>
<intersection>-4300.5 2</intersection>
<intersection>-4152.5 3</intersection>
<intersection>-4134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-4134.5,-7.5,-4134.5</points>
<connection>
<GID>1468</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4300.5,-109,-4300.5</points>
<connection>
<GID>1365</GID>
<name>OUT_5</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-4152.5,-26,-4152.5</points>
<connection>
<GID>1469</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-4154.5,589,-4154.5</points>
<connection>
<GID>1469</GID>
<name>OUT_0</name></connection>
<intersection>34 38</intersection>
<intersection>108 43</intersection>
<intersection>192 42</intersection>
<intersection>266 45</intersection>
<intersection>357 47</intersection>
<intersection>431 49</intersection>
<intersection>515 51</intersection>
<intersection>589 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34,-4154.5,34,-4142</points>
<connection>
<GID>1447</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192,-4154.5,192,-4144</points>
<connection>
<GID>1453</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108,-4154.5,108,-4142</points>
<connection>
<GID>1444</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266,-4154.5,266,-4144</points>
<connection>
<GID>1450</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357,-4154.5,357,-4145.5</points>
<connection>
<GID>1459</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431,-4154.5,431,-4145.5</points>
<connection>
<GID>1456</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515,-4154.5,515,-4147.5</points>
<connection>
<GID>1465</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589,-4154.5,589,-4147.5</points>
<connection>
<GID>1462</GID>
<name>IN_1</name></connection>
<intersection>-4154.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-4141,49.5,-4141</points>
<connection>
<GID>1447</GID>
<name>OUT</name></connection>
<connection>
<GID>1446</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-4149.5,31,-4132.5</points>
<intersection>-4149.5 3</intersection>
<intersection>-4140 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-4140,34,-4140</points>
<connection>
<GID>1447</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-4132.5,31,-4132.5</points>
<connection>
<GID>1445</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-4149.5,51.5,-4149.5</points>
<intersection>31 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-4149.5,51.5,-4144</points>
<connection>
<GID>1446</GID>
<name>IN_0</name></connection>
<intersection>-4149.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114,-4141,123,-4141</points>
<connection>
<GID>1444</GID>
<name>OUT</name></connection>
<connection>
<GID>1449</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-4151,104.5,-4132.5</points>
<intersection>-4151 3</intersection>
<intersection>-4140 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-4140,108,-4140</points>
<connection>
<GID>1444</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-4132.5,104.5,-4132.5</points>
<connection>
<GID>1448</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-4151,125,-4151</points>
<intersection>104.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-4151,125,-4144</points>
<connection>
<GID>1449</GID>
<name>IN_0</name></connection>
<intersection>-4151 3</intersection></vsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-4143,207.5,-4143</points>
<connection>
<GID>1453</GID>
<name>OUT</name></connection>
<connection>
<GID>1452</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-4151.5,189,-4132.5</points>
<intersection>-4151.5 3</intersection>
<intersection>-4142 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-4142,192,-4142</points>
<connection>
<GID>1453</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188,-4132.5,189,-4132.5</points>
<connection>
<GID>1451</GID>
<name>OUT_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189,-4151.5,209.5,-4151.5</points>
<intersection>189 0</intersection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,-4151.5,209.5,-4146</points>
<connection>
<GID>1452</GID>
<name>IN_0</name></connection>
<intersection>-4151.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272,-4143,281,-4143</points>
<connection>
<GID>1450</GID>
<name>OUT</name></connection>
<connection>
<GID>1455</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-4153,262.5,-4132.5</points>
<connection>
<GID>1454</GID>
<name>OUT_0</name></connection>
<intersection>-4153 3</intersection>
<intersection>-4142 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-4142,266,-4142</points>
<connection>
<GID>1450</GID>
<name>IN_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262.5,-4153,283,-4153</points>
<intersection>262.5 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-4153,283,-4146</points>
<connection>
<GID>1455</GID>
<name>IN_0</name></connection>
<intersection>-4153 3</intersection></vsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363,-4144.5,372.5,-4144.5</points>
<connection>
<GID>1459</GID>
<name>OUT</name></connection>
<connection>
<GID>1458</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-4153,354,-4132.5</points>
<intersection>-4153 3</intersection>
<intersection>-4143.5 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-4143.5,357,-4143.5</points>
<connection>
<GID>1459</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-4132.5,354,-4132.5</points>
<connection>
<GID>1457</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354,-4153,374.5,-4153</points>
<intersection>354 0</intersection>
<intersection>374.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374.5,-4153,374.5,-4147.5</points>
<connection>
<GID>1458</GID>
<name>IN_0</name></connection>
<intersection>-4153 3</intersection></vsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437,-4144.5,446,-4144.5</points>
<connection>
<GID>1456</GID>
<name>OUT</name></connection>
<connection>
<GID>1461</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-4153,427.5,-4132.5</points>
<intersection>-4153 3</intersection>
<intersection>-4143.5 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-4143.5,431,-4143.5</points>
<connection>
<GID>1456</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426.5,-4132.5,427.5,-4132.5</points>
<connection>
<GID>1460</GID>
<name>OUT_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-4153,448,-4153</points>
<intersection>427.5 0</intersection>
<intersection>448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448,-4153,448,-4147.5</points>
<connection>
<GID>1461</GID>
<name>IN_0</name></connection>
<intersection>-4153 3</intersection></vsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521,-4146.5,530.5,-4146.5</points>
<connection>
<GID>1465</GID>
<name>OUT</name></connection>
<connection>
<GID>1464</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1001</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,-4152.5,512,-4132.5</points>
<intersection>-4152.5 3</intersection>
<intersection>-4145.5 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-4145.5,515,-4145.5</points>
<connection>
<GID>1465</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,-4132.5,512,-4132.5</points>
<connection>
<GID>1463</GID>
<name>OUT_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512,-4152.5,532.5,-4152.5</points>
<intersection>512 0</intersection>
<intersection>532.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532.5,-4152.5,532.5,-4149.5</points>
<connection>
<GID>1464</GID>
<name>IN_0</name></connection>
<intersection>-4152.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595,-4146.5,604,-4146.5</points>
<connection>
<GID>1462</GID>
<name>OUT</name></connection>
<connection>
<GID>1467</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1003</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-4152.5,585.5,-4132.5</points>
<intersection>-4152.5 3</intersection>
<intersection>-4145.5 1</intersection>
<intersection>-4132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-4145.5,589,-4145.5</points>
<connection>
<GID>1462</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,-4132.5,585.5,-4132.5</points>
<connection>
<GID>1466</GID>
<name>OUT_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-4152.5,606,-4152.5</points>
<intersection>585.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-4152.5,606,-4149.5</points>
<connection>
<GID>1467</GID>
<name>IN_0</name></connection>
<intersection>-4152.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-4135.5,578.5,-4135.5</points>
<connection>
<GID>1468</GID>
<name>OUT</name></connection>
<connection>
<GID>1466</GID>
<name>clock</name></connection>
<connection>
<GID>1463</GID>
<name>clock</name></connection>
<connection>
<GID>1460</GID>
<name>clock</name></connection>
<connection>
<GID>1457</GID>
<name>clock</name></connection>
<connection>
<GID>1454</GID>
<name>clock</name></connection>
<connection>
<GID>1451</GID>
<name>clock</name></connection>
<connection>
<GID>1448</GID>
<name>clock</name></connection>
<connection>
<GID>1445</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-4450.5,-109,-4303.5</points>
<intersection>-4450.5 3</intersection>
<intersection>-4432.5 1</intersection>
<intersection>-4303.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-4432.5,-6.5,-4432.5</points>
<connection>
<GID>1494</GID>
<name>IN_0</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4303.5,-109,-4303.5</points>
<connection>
<GID>1365</GID>
<name>OUT_2</name></connection>
<intersection>-109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-109,-4450.5,-25,-4450.5</points>
<connection>
<GID>1495</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-22.5,-4452.5,590,-4452.5</points>
<connection>
<GID>1495</GID>
<name>OUT_0</name></connection>
<intersection>35 38</intersection>
<intersection>109 43</intersection>
<intersection>193 42</intersection>
<intersection>267 45</intersection>
<intersection>358 47</intersection>
<intersection>432 49</intersection>
<intersection>516 51</intersection>
<intersection>590 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>35,-4452.5,35,-4440</points>
<connection>
<GID>1473</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>193,-4452.5,193,-4442</points>
<connection>
<GID>1479</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>109,-4452.5,109,-4440</points>
<connection>
<GID>1470</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>267,-4452.5,267,-4442</points>
<connection>
<GID>1476</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>358,-4452.5,358,-4443.5</points>
<connection>
<GID>1485</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>432,-4452.5,432,-4443.5</points>
<connection>
<GID>1482</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>516,-4452.5,516,-4445.5</points>
<connection>
<GID>1491</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>590,-4452.5,590,-4445.5</points>
<connection>
<GID>1488</GID>
<name>IN_1</name></connection>
<intersection>-4452.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-4439,50.5,-4439</points>
<connection>
<GID>1473</GID>
<name>OUT</name></connection>
<connection>
<GID>1472</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-4447.5,32,-4430.5</points>
<intersection>-4447.5 3</intersection>
<intersection>-4438 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-4438,35,-4438</points>
<connection>
<GID>1473</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-4430.5,32,-4430.5</points>
<connection>
<GID>1471</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-4447.5,52.5,-4447.5</points>
<intersection>32 0</intersection>
<intersection>52.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52.5,-4447.5,52.5,-4442</points>
<connection>
<GID>1472</GID>
<name>IN_0</name></connection>
<intersection>-4447.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115,-4439,124,-4439</points>
<connection>
<GID>1470</GID>
<name>OUT</name></connection>
<connection>
<GID>1475</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-4449,105.5,-4430.5</points>
<intersection>-4449 3</intersection>
<intersection>-4438 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-4438,109,-4438</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-4430.5,105.5,-4430.5</points>
<connection>
<GID>1474</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105.5,-4449,126,-4449</points>
<intersection>105.5 0</intersection>
<intersection>126 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>126,-4449,126,-4442</points>
<connection>
<GID>1475</GID>
<name>IN_0</name></connection>
<intersection>-4449 3</intersection></vsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199,-4441,208.5,-4441</points>
<connection>
<GID>1479</GID>
<name>OUT</name></connection>
<connection>
<GID>1478</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-4449.5,190,-4430.5</points>
<intersection>-4449.5 3</intersection>
<intersection>-4440 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-4440,193,-4440</points>
<connection>
<GID>1479</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,-4430.5,190,-4430.5</points>
<connection>
<GID>1477</GID>
<name>OUT_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>190,-4449.5,210.5,-4449.5</points>
<intersection>190 0</intersection>
<intersection>210.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210.5,-4449.5,210.5,-4444</points>
<connection>
<GID>1478</GID>
<name>IN_0</name></connection>
<intersection>-4449.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>273,-4441,282,-4441</points>
<connection>
<GID>1476</GID>
<name>OUT</name></connection>
<connection>
<GID>1481</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,-4451,263.5,-4430.5</points>
<intersection>-4451 3</intersection>
<intersection>-4440 1</intersection>
<intersection>-4430.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263.5,-4440,267,-4440</points>
<connection>
<GID>1476</GID>
<name>IN_0</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263.5,-4451,284,-4451</points>
<intersection>263.5 0</intersection>
<intersection>284 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>284,-4451,284,-4444</points>
<connection>
<GID>1481</GID>
<name>IN_0</name></connection>
<intersection>-4451 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>262.5,-4430.5,263.5,-4430.5</points>
<connection>
<GID>1480</GID>
<name>OUT_0</name></connection>
<intersection>263.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364,-4442.5,373.5,-4442.5</points>
<connection>
<GID>1485</GID>
<name>OUT</name></connection>
<connection>
<GID>1484</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,-4451,355,-4430.5</points>
<intersection>-4451 3</intersection>
<intersection>-4441.5 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-4441.5,358,-4441.5</points>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>354,-4430.5,355,-4430.5</points>
<connection>
<GID>1483</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>355,-4451,375.5,-4451</points>
<intersection>355 0</intersection>
<intersection>375.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375.5,-4451,375.5,-4445.5</points>
<connection>
<GID>1484</GID>
<name>IN_0</name></connection>
<intersection>-4451 3</intersection></vsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>438,-4442.5,447,-4442.5</points>
<connection>
<GID>1482</GID>
<name>OUT</name></connection>
<connection>
<GID>1487</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,-4451,428.5,-4430.5</points>
<intersection>-4451 3</intersection>
<intersection>-4441.5 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,-4441.5,432,-4441.5</points>
<connection>
<GID>1482</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,-4430.5,428.5,-4430.5</points>
<connection>
<GID>1486</GID>
<name>OUT_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428.5,-4451,449,-4451</points>
<intersection>428.5 0</intersection>
<intersection>449 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>449,-4451,449,-4445.5</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<intersection>-4451 3</intersection></vsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,-4444.5,531.5,-4444.5</points>
<connection>
<GID>1491</GID>
<name>OUT</name></connection>
<connection>
<GID>1490</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,-4450.5,513,-4430.5</points>
<intersection>-4450.5 3</intersection>
<intersection>-4443.5 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513,-4443.5,516,-4443.5</points>
<connection>
<GID>1491</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>512,-4430.5,513,-4430.5</points>
<connection>
<GID>1489</GID>
<name>OUT_0</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>513,-4450.5,533.5,-4450.5</points>
<intersection>513 0</intersection>
<intersection>533.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533.5,-4450.5,533.5,-4447.5</points>
<connection>
<GID>1490</GID>
<name>IN_0</name></connection>
<intersection>-4450.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>596,-4444.5,605,-4444.5</points>
<connection>
<GID>1488</GID>
<name>OUT</name></connection>
<connection>
<GID>1493</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,-4450.5,586.5,-4430.5</points>
<intersection>-4450.5 3</intersection>
<intersection>-4443.5 1</intersection>
<intersection>-4430.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586.5,-4443.5,590,-4443.5</points>
<connection>
<GID>1488</GID>
<name>IN_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585.5,-4430.5,586.5,-4430.5</points>
<connection>
<GID>1492</GID>
<name>OUT_0</name></connection>
<intersection>586.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586.5,-4450.5,607,-4450.5</points>
<intersection>586.5 0</intersection>
<intersection>607 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>607,-4450.5,607,-4447.5</points>
<connection>
<GID>1493</GID>
<name>IN_0</name></connection>
<intersection>-4450.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-4433.5,579.5,-4433.5</points>
<connection>
<GID>1480</GID>
<name>clock</name></connection>
<connection>
<GID>1494</GID>
<name>OUT</name></connection>
<connection>
<GID>1492</GID>
<name>clock</name></connection>
<connection>
<GID>1486</GID>
<name>clock</name></connection>
<connection>
<GID>1483</GID>
<name>clock</name></connection>
<connection>
<GID>1477</GID>
<name>clock</name></connection>
<connection>
<GID>1474</GID>
<name>clock</name></connection>
<connection>
<GID>1471</GID>
<name>clock</name></connection>
<connection>
<GID>1489</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-4360.5,-108,-4302.5</points>
<intersection>-4360.5 3</intersection>
<intersection>-4342.5 1</intersection>
<intersection>-4302.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-4342.5,-9.5,-4342.5</points>
<connection>
<GID>1311</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4302.5,-108,-4302.5</points>
<connection>
<GID>1365</GID>
<name>OUT_3</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-4360.5,-28,-4360.5</points>
<connection>
<GID>1312</GID>
<name>ENABLE_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25.5,-4362.5,587,-4362.5</points>
<connection>
<GID>1312</GID>
<name>OUT_0</name></connection>
<intersection>32 38</intersection>
<intersection>106 43</intersection>
<intersection>190 42</intersection>
<intersection>264 45</intersection>
<intersection>355 47</intersection>
<intersection>429 49</intersection>
<intersection>513 51</intersection>
<intersection>587 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32,-4362.5,32,-4350</points>
<connection>
<GID>1499</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190,-4362.5,190,-4352</points>
<connection>
<GID>1296</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106,-4362.5,106,-4350</points>
<connection>
<GID>1496</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264,-4362.5,264,-4352</points>
<connection>
<GID>1502</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355,-4362.5,355,-4353.5</points>
<connection>
<GID>1302</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429,-4362.5,429,-4353.5</points>
<connection>
<GID>1299</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513,-4362.5,513,-4355.5</points>
<connection>
<GID>1308</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587,-4362.5,587,-4355.5</points>
<connection>
<GID>1305</GID>
<name>IN_1</name></connection>
<intersection>-4362.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-4349,47.5,-4349</points>
<connection>
<GID>1499</GID>
<name>OUT</name></connection>
<connection>
<GID>1498</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-4357.5,29,-4340.5</points>
<intersection>-4357.5 3</intersection>
<intersection>-4348 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-4348,32,-4348</points>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-4340.5,29,-4340.5</points>
<connection>
<GID>1497</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-4357.5,49.5,-4357.5</points>
<intersection>29 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-4357.5,49.5,-4352</points>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection>
<intersection>-4357.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112,-4349,121,-4349</points>
<connection>
<GID>1496</GID>
<name>OUT</name></connection>
<connection>
<GID>1501</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-4359,102.5,-4340.5</points>
<intersection>-4359 3</intersection>
<intersection>-4348 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-4348,106,-4348</points>
<connection>
<GID>1496</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-4340.5,102.5,-4340.5</points>
<connection>
<GID>1500</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-4359,123,-4359</points>
<intersection>102.5 0</intersection>
<intersection>123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123,-4359,123,-4352</points>
<connection>
<GID>1501</GID>
<name>IN_0</name></connection>
<intersection>-4359 3</intersection></vsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,-4351,205.5,-4351</points>
<connection>
<GID>1296</GID>
<name>OUT</name></connection>
<connection>
<GID>1504</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-4359.5,187,-4340.5</points>
<intersection>-4359.5 3</intersection>
<intersection>-4350 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-4350,190,-4350</points>
<connection>
<GID>1296</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-4340.5,187,-4340.5</points>
<connection>
<GID>1503</GID>
<name>OUT_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,-4359.5,207.5,-4359.5</points>
<intersection>187 0</intersection>
<intersection>207.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207.5,-4359.5,207.5,-4354</points>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>-4359.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270,-4351,279,-4351</points>
<connection>
<GID>1502</GID>
<name>OUT</name></connection>
<connection>
<GID>1298</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-4361,260.5,-4340.5</points>
<connection>
<GID>1297</GID>
<name>OUT_0</name></connection>
<intersection>-4361 3</intersection>
<intersection>-4350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-4350,264,-4350</points>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-4361,281,-4361</points>
<intersection>260.5 0</intersection>
<intersection>281 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281,-4361,281,-4354</points>
<connection>
<GID>1298</GID>
<name>IN_0</name></connection>
<intersection>-4361 3</intersection></vsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-4352.5,370.5,-4352.5</points>
<connection>
<GID>1302</GID>
<name>OUT</name></connection>
<connection>
<GID>1301</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-4361,352,-4340.5</points>
<intersection>-4361 3</intersection>
<intersection>-4351.5 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-4351.5,355,-4351.5</points>
<connection>
<GID>1302</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-4340.5,352,-4340.5</points>
<connection>
<GID>1300</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352,-4361,372.5,-4361</points>
<intersection>352 0</intersection>
<intersection>372.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372.5,-4361,372.5,-4355.5</points>
<connection>
<GID>1301</GID>
<name>IN_0</name></connection>
<intersection>-4361 3</intersection></vsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435,-4352.5,444,-4352.5</points>
<connection>
<GID>1299</GID>
<name>OUT</name></connection>
<connection>
<GID>1304</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-4361,425.5,-4340.5</points>
<intersection>-4361 3</intersection>
<intersection>-4351.5 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,-4351.5,429,-4351.5</points>
<connection>
<GID>1299</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,-4340.5,425.5,-4340.5</points>
<connection>
<GID>1303</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,-4361,446,-4361</points>
<intersection>425.5 0</intersection>
<intersection>446 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446,-4361,446,-4355.5</points>
<connection>
<GID>1304</GID>
<name>IN_0</name></connection>
<intersection>-4361 3</intersection></vsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-4354.5,528.5,-4354.5</points>
<connection>
<GID>1308</GID>
<name>OUT</name></connection>
<connection>
<GID>1307</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,-4360.5,510,-4340.5</points>
<intersection>-4360.5 3</intersection>
<intersection>-4353.5 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,-4353.5,513,-4353.5</points>
<connection>
<GID>1308</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509,-4340.5,510,-4340.5</points>
<connection>
<GID>1306</GID>
<name>OUT_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510,-4360.5,530.5,-4360.5</points>
<intersection>510 0</intersection>
<intersection>530.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530.5,-4360.5,530.5,-4357.5</points>
<connection>
<GID>1307</GID>
<name>IN_0</name></connection>
<intersection>-4360.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593,-4354.5,602,-4354.5</points>
<connection>
<GID>1305</GID>
<name>OUT</name></connection>
<connection>
<GID>1310</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-4360.5,583.5,-4340.5</points>
<intersection>-4360.5 3</intersection>
<intersection>-4353.5 1</intersection>
<intersection>-4340.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,-4353.5,587,-4353.5</points>
<connection>
<GID>1305</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,-4340.5,583.5,-4340.5</points>
<connection>
<GID>1309</GID>
<name>OUT_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583.5,-4360.5,604,-4360.5</points>
<intersection>583.5 0</intersection>
<intersection>604 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604,-4360.5,604,-4357.5</points>
<connection>
<GID>1310</GID>
<name>IN_0</name></connection>
<intersection>-4360.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,-4343.5,576.5,-4343.5</points>
<connection>
<GID>1503</GID>
<name>clock</name></connection>
<connection>
<GID>1500</GID>
<name>clock</name></connection>
<connection>
<GID>1497</GID>
<name>clock</name></connection>
<connection>
<GID>1311</GID>
<name>OUT</name></connection>
<connection>
<GID>1309</GID>
<name>clock</name></connection>
<connection>
<GID>1306</GID>
<name>clock</name></connection>
<connection>
<GID>1303</GID>
<name>clock</name></connection>
<connection>
<GID>1300</GID>
<name>clock</name></connection>
<connection>
<GID>1297</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-4618.5,-112,-4305.5</points>
<intersection>-4618.5 3</intersection>
<intersection>-4600.5 1</intersection>
<intersection>-4305.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112,-4600.5,-2.5,-4600.5</points>
<connection>
<GID>1337</GID>
<name>IN_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4305.5,-112,-4305.5</points>
<connection>
<GID>1365</GID>
<name>OUT_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112,-4618.5,-21,-4618.5</points>
<connection>
<GID>1338</GID>
<name>ENABLE_0</name></connection>
<intersection>-112 0</intersection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-18.5,-4620.5,594,-4620.5</points>
<connection>
<GID>1338</GID>
<name>OUT_0</name></connection>
<intersection>39 38</intersection>
<intersection>113 43</intersection>
<intersection>197 42</intersection>
<intersection>271 45</intersection>
<intersection>362 47</intersection>
<intersection>436 49</intersection>
<intersection>520 51</intersection>
<intersection>594 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>39,-4620.5,39,-4608</points>
<connection>
<GID>1316</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>197,-4620.5,197,-4610</points>
<connection>
<GID>1322</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>113,-4620.5,113,-4608</points>
<connection>
<GID>1313</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>271,-4620.5,271,-4610</points>
<connection>
<GID>1319</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>362,-4620.5,362,-4611.5</points>
<connection>
<GID>1328</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>436,-4620.5,436,-4611.5</points>
<connection>
<GID>1325</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>520,-4620.5,520,-4613.5</points>
<connection>
<GID>1334</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>594,-4620.5,594,-4613.5</points>
<connection>
<GID>1331</GID>
<name>IN_1</name></connection>
<intersection>-4620.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-4607,54.5,-4607</points>
<connection>
<GID>1316</GID>
<name>OUT</name></connection>
<connection>
<GID>1315</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-4615.5,36,-4598.5</points>
<intersection>-4615.5 3</intersection>
<intersection>-4606 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-4606,39,-4606</points>
<connection>
<GID>1316</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-4598.5,36,-4598.5</points>
<connection>
<GID>1314</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-4615.5,56.5,-4615.5</points>
<intersection>36 0</intersection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56.5,-4615.5,56.5,-4610</points>
<connection>
<GID>1315</GID>
<name>IN_0</name></connection>
<intersection>-4615.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119,-4607,128,-4607</points>
<connection>
<GID>1313</GID>
<name>OUT</name></connection>
<connection>
<GID>1318</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-4617,109.5,-4598.5</points>
<intersection>-4617 3</intersection>
<intersection>-4606 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-4606,113,-4606</points>
<connection>
<GID>1313</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-4598.5,109.5,-4598.5</points>
<connection>
<GID>1317</GID>
<name>OUT_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-4617,130,-4617</points>
<intersection>109.5 0</intersection>
<intersection>130 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130,-4617,130,-4610</points>
<connection>
<GID>1318</GID>
<name>IN_0</name></connection>
<intersection>-4617 3</intersection></vsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,-4609,212.5,-4609</points>
<connection>
<GID>1322</GID>
<name>OUT</name></connection>
<connection>
<GID>1321</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-4617.5,194,-4598.5</points>
<intersection>-4617.5 3</intersection>
<intersection>-4608 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,-4608,197,-4608</points>
<connection>
<GID>1322</GID>
<name>IN_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>193,-4598.5,194,-4598.5</points>
<connection>
<GID>1320</GID>
<name>OUT_0</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>194,-4617.5,214.5,-4617.5</points>
<intersection>194 0</intersection>
<intersection>214.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>214.5,-4617.5,214.5,-4612</points>
<connection>
<GID>1321</GID>
<name>IN_0</name></connection>
<intersection>-4617.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>277,-4609,286,-4609</points>
<connection>
<GID>1319</GID>
<name>OUT</name></connection>
<connection>
<GID>1324</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-4619,267.5,-4598.5</points>
<connection>
<GID>1323</GID>
<name>OUT_0</name></connection>
<intersection>-4619 3</intersection>
<intersection>-4608 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-4608,271,-4608</points>
<connection>
<GID>1319</GID>
<name>IN_0</name></connection>
<intersection>267.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>267.5,-4619,288,-4619</points>
<intersection>267.5 0</intersection>
<intersection>288 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>288,-4619,288,-4612</points>
<connection>
<GID>1324</GID>
<name>IN_0</name></connection>
<intersection>-4619 3</intersection></vsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368,-4610.5,377.5,-4610.5</points>
<connection>
<GID>1328</GID>
<name>OUT</name></connection>
<connection>
<GID>1327</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-4619,359,-4598.5</points>
<intersection>-4619 3</intersection>
<intersection>-4609.5 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-4609.5,362,-4609.5</points>
<connection>
<GID>1328</GID>
<name>IN_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>358,-4598.5,359,-4598.5</points>
<connection>
<GID>1326</GID>
<name>OUT_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>359,-4619,379.5,-4619</points>
<intersection>359 0</intersection>
<intersection>379.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>379.5,-4619,379.5,-4613.5</points>
<connection>
<GID>1327</GID>
<name>IN_0</name></connection>
<intersection>-4619 3</intersection></vsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>442,-4610.5,451,-4610.5</points>
<connection>
<GID>1325</GID>
<name>OUT</name></connection>
<connection>
<GID>1330</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,-4619,432.5,-4598.5</points>
<intersection>-4619 3</intersection>
<intersection>-4609.5 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,-4609.5,436,-4609.5</points>
<connection>
<GID>1325</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-4598.5,432.5,-4598.5</points>
<connection>
<GID>1329</GID>
<name>OUT_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432.5,-4619,453,-4619</points>
<intersection>432.5 0</intersection>
<intersection>453 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>453,-4619,453,-4613.5</points>
<connection>
<GID>1330</GID>
<name>IN_0</name></connection>
<intersection>-4619 3</intersection></vsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>526,-4612.5,535.5,-4612.5</points>
<connection>
<GID>1334</GID>
<name>OUT</name></connection>
<connection>
<GID>1333</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,-4618.5,517,-4598.5</points>
<intersection>-4618.5 3</intersection>
<intersection>-4611.5 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,-4611.5,520,-4611.5</points>
<connection>
<GID>1334</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>516,-4598.5,517,-4598.5</points>
<connection>
<GID>1332</GID>
<name>OUT_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>517,-4618.5,537.5,-4618.5</points>
<intersection>517 0</intersection>
<intersection>537.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>537.5,-4618.5,537.5,-4615.5</points>
<connection>
<GID>1333</GID>
<name>IN_0</name></connection>
<intersection>-4618.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>600,-4612.5,609,-4612.5</points>
<connection>
<GID>1331</GID>
<name>OUT</name></connection>
<connection>
<GID>1336</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,-4618.5,590.5,-4598.5</points>
<intersection>-4618.5 3</intersection>
<intersection>-4611.5 1</intersection>
<intersection>-4598.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,-4611.5,594,-4611.5</points>
<connection>
<GID>1331</GID>
<name>IN_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,-4598.5,590.5,-4598.5</points>
<connection>
<GID>1335</GID>
<name>OUT_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>590.5,-4618.5,611,-4618.5</points>
<intersection>590.5 0</intersection>
<intersection>611 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>611,-4618.5,611,-4615.5</points>
<connection>
<GID>1336</GID>
<name>IN_0</name></connection>
<intersection>-4618.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-4601.5,583.5,-4601.5</points>
<connection>
<GID>1337</GID>
<name>OUT</name></connection>
<connection>
<GID>1335</GID>
<name>clock</name></connection>
<connection>
<GID>1332</GID>
<name>clock</name></connection>
<connection>
<GID>1329</GID>
<name>clock</name></connection>
<connection>
<GID>1326</GID>
<name>clock</name></connection>
<connection>
<GID>1323</GID>
<name>clock</name></connection>
<connection>
<GID>1320</GID>
<name>clock</name></connection>
<connection>
<GID>1317</GID>
<name>clock</name></connection>
<connection>
<GID>1314</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-4528.5,-110,-4304.5</points>
<intersection>-4528.5 3</intersection>
<intersection>-4510.5 1</intersection>
<intersection>-4304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110,-4510.5,-5.5,-4510.5</points>
<connection>
<GID>1363</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-118.5,-4304.5,-110,-4304.5</points>
<connection>
<GID>1365</GID>
<name>OUT_1</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110,-4528.5,-24,-4528.5</points>
<connection>
<GID>1364</GID>
<name>ENABLE_0</name></connection>
<intersection>-110 0</intersection></hsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21.5,-4530.5,591,-4530.5</points>
<connection>
<GID>1364</GID>
<name>OUT_0</name></connection>
<intersection>36 38</intersection>
<intersection>110 43</intersection>
<intersection>194 42</intersection>
<intersection>268 45</intersection>
<intersection>359 47</intersection>
<intersection>433 49</intersection>
<intersection>517 51</intersection>
<intersection>591 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36,-4530.5,36,-4518</points>
<connection>
<GID>1342</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194,-4530.5,194,-4520</points>
<connection>
<GID>1348</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110,-4530.5,110,-4518</points>
<connection>
<GID>1339</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268,-4530.5,268,-4520</points>
<connection>
<GID>1345</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359,-4530.5,359,-4521.5</points>
<connection>
<GID>1354</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433,-4530.5,433,-4521.5</points>
<connection>
<GID>1351</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517,-4530.5,517,-4523.5</points>
<connection>
<GID>1360</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591,-4530.5,591,-4523.5</points>
<connection>
<GID>1357</GID>
<name>IN_1</name></connection>
<intersection>-4530.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-4517,51.5,-4517</points>
<connection>
<GID>1342</GID>
<name>OUT</name></connection>
<connection>
<GID>1341</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-4525.5,33,-4508.5</points>
<intersection>-4525.5 3</intersection>
<intersection>-4516 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-4516,36,-4516</points>
<connection>
<GID>1342</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-4508.5,33,-4508.5</points>
<connection>
<GID>1340</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-4525.5,53.5,-4525.5</points>
<intersection>33 0</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-4525.5,53.5,-4520</points>
<connection>
<GID>1341</GID>
<name>IN_0</name></connection>
<intersection>-4525.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116,-4517,125,-4517</points>
<connection>
<GID>1339</GID>
<name>OUT</name></connection>
<connection>
<GID>1344</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-4527,106.5,-4508.5</points>
<intersection>-4527 3</intersection>
<intersection>-4516 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-4516,110,-4516</points>
<connection>
<GID>1339</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-4508.5,106.5,-4508.5</points>
<connection>
<GID>1343</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,-4527,127,-4527</points>
<intersection>106.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-4527,127,-4520</points>
<connection>
<GID>1344</GID>
<name>IN_0</name></connection>
<intersection>-4527 3</intersection></vsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-4519,209.5,-4519</points>
<connection>
<GID>1348</GID>
<name>OUT</name></connection>
<connection>
<GID>1347</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-4527.5,191,-4508.5</points>
<intersection>-4527.5 3</intersection>
<intersection>-4518 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-4518,194,-4518</points>
<connection>
<GID>1348</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,-4508.5,191,-4508.5</points>
<connection>
<GID>1346</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191,-4527.5,211.5,-4527.5</points>
<intersection>191 0</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211.5,-4527.5,211.5,-4522</points>
<connection>
<GID>1347</GID>
<name>IN_0</name></connection>
<intersection>-4527.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274,-4519,283,-4519</points>
<connection>
<GID>1345</GID>
<name>OUT</name></connection>
<connection>
<GID>1350</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-4529,264.5,-4508.5</points>
<connection>
<GID>1349</GID>
<name>OUT_0</name></connection>
<intersection>-4529 3</intersection>
<intersection>-4518 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-4518,268,-4518</points>
<connection>
<GID>1345</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264.5,-4529,285,-4529</points>
<intersection>264.5 0</intersection>
<intersection>285 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285,-4529,285,-4522</points>
<connection>
<GID>1350</GID>
<name>IN_0</name></connection>
<intersection>-4529 3</intersection></vsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365,-4520.5,374.5,-4520.5</points>
<connection>
<GID>1354</GID>
<name>OUT</name></connection>
<connection>
<GID>1353</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-4529,356,-4508.5</points>
<intersection>-4529 3</intersection>
<intersection>-4519.5 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-4519.5,359,-4519.5</points>
<connection>
<GID>1354</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355,-4508.5,356,-4508.5</points>
<connection>
<GID>1352</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356,-4529,376.5,-4529</points>
<intersection>356 0</intersection>
<intersection>376.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376.5,-4529,376.5,-4523.5</points>
<connection>
<GID>1353</GID>
<name>IN_0</name></connection>
<intersection>-4529 3</intersection></vsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439,-4520.5,448,-4520.5</points>
<connection>
<GID>1351</GID>
<name>OUT</name></connection>
<connection>
<GID>1356</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-4529,429.5,-4508.5</points>
<intersection>-4529 3</intersection>
<intersection>-4519.5 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,-4519.5,433,-4519.5</points>
<connection>
<GID>1351</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,-4508.5,429.5,-4508.5</points>
<connection>
<GID>1355</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,-4529,450,-4529</points>
<intersection>429.5 0</intersection>
<intersection>450 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450,-4529,450,-4523.5</points>
<connection>
<GID>1356</GID>
<name>IN_0</name></connection>
<intersection>-4529 3</intersection></vsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523,-4522.5,532.5,-4522.5</points>
<connection>
<GID>1360</GID>
<name>OUT</name></connection>
<connection>
<GID>1359</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-4528.5,514,-4508.5</points>
<intersection>-4528.5 3</intersection>
<intersection>-4521.5 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-4521.5,517,-4521.5</points>
<connection>
<GID>1360</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,-4508.5,514,-4508.5</points>
<connection>
<GID>1358</GID>
<name>OUT_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514,-4528.5,534.5,-4528.5</points>
<intersection>514 0</intersection>
<intersection>534.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534.5,-4528.5,534.5,-4525.5</points>
<connection>
<GID>1359</GID>
<name>IN_0</name></connection>
<intersection>-4528.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597,-4522.5,606,-4522.5</points>
<connection>
<GID>1357</GID>
<name>OUT</name></connection>
<connection>
<GID>1362</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,-4528.5,587.5,-4508.5</points>
<intersection>-4528.5 3</intersection>
<intersection>-4521.5 1</intersection>
<intersection>-4508.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,-4521.5,591,-4521.5</points>
<connection>
<GID>1357</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586.5,-4508.5,587.5,-4508.5</points>
<connection>
<GID>1361</GID>
<name>OUT_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587.5,-4528.5,608,-4528.5</points>
<intersection>587.5 0</intersection>
<intersection>608 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608,-4528.5,608,-4525.5</points>
<connection>
<GID>1362</GID>
<name>IN_0</name></connection>
<intersection>-4528.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-4511.5,580.5,-4511.5</points>
<connection>
<GID>1363</GID>
<name>OUT</name></connection>
<connection>
<GID>1361</GID>
<name>clock</name></connection>
<connection>
<GID>1358</GID>
<name>clock</name></connection>
<connection>
<GID>1355</GID>
<name>clock</name></connection>
<connection>
<GID>1352</GID>
<name>clock</name></connection>
<connection>
<GID>1349</GID>
<name>clock</name></connection>
<connection>
<GID>1346</GID>
<name>clock</name></connection>
<connection>
<GID>1343</GID>
<name>clock</name></connection>
<connection>
<GID>1340</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112.5,-5224,-112.5,-4981</points>
<intersection>-5224 2</intersection>
<intersection>-4999 3</intersection>
<intersection>-4981 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112.5,-4981,-11,-4981</points>
<connection>
<GID>1599</GID>
<name>IN_0</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5224,-112.5,-5224</points>
<connection>
<GID>1574</GID>
<name>OUT_6</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112.5,-4999,-29.5,-4999</points>
<connection>
<GID>1600</GID>
<name>ENABLE_0</name></connection>
<intersection>-112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-27,-5001,585.5,-5001</points>
<connection>
<GID>1600</GID>
<name>OUT_0</name></connection>
<intersection>30.5 38</intersection>
<intersection>104.5 43</intersection>
<intersection>188.5 42</intersection>
<intersection>262.5 45</intersection>
<intersection>353.5 47</intersection>
<intersection>427.5 49</intersection>
<intersection>511.5 51</intersection>
<intersection>585.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>30.5,-5001,30.5,-4988.5</points>
<connection>
<GID>1578</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>188.5,-5001,188.5,-4990.5</points>
<connection>
<GID>1584</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>104.5,-5001,104.5,-4988.5</points>
<connection>
<GID>1575</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>262.5,-5001,262.5,-4990.5</points>
<connection>
<GID>1581</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>353.5,-5001,353.5,-4992</points>
<connection>
<GID>1590</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>427.5,-5001,427.5,-4992</points>
<connection>
<GID>1587</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>511.5,-5001,511.5,-4994</points>
<connection>
<GID>1596</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>585.5,-5001,585.5,-4994</points>
<connection>
<GID>1593</GID>
<name>IN_1</name></connection>
<intersection>-5001 33</intersection></vsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-4987.5,46,-4987.5</points>
<connection>
<GID>1578</GID>
<name>OUT</name></connection>
<connection>
<GID>1577</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-4996,27.5,-4979</points>
<intersection>-4996 3</intersection>
<intersection>-4986.5 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-4986.5,30.5,-4986.5</points>
<connection>
<GID>1578</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-4979,27.5,-4979</points>
<connection>
<GID>1576</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-4996,48,-4996</points>
<intersection>27.5 0</intersection>
<intersection>48 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48,-4996,48,-4990.5</points>
<connection>
<GID>1577</GID>
<name>IN_0</name></connection>
<intersection>-4996 3</intersection></vsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>110.5,-4987.5,119.5,-4987.5</points>
<connection>
<GID>1575</GID>
<name>OUT</name></connection>
<connection>
<GID>1580</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-4997.5,101,-4979</points>
<intersection>-4997.5 3</intersection>
<intersection>-4986.5 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-4986.5,104.5,-4986.5</points>
<connection>
<GID>1575</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-4979,101,-4979</points>
<connection>
<GID>1579</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101,-4997.5,121.5,-4997.5</points>
<intersection>101 0</intersection>
<intersection>121.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>121.5,-4997.5,121.5,-4990.5</points>
<connection>
<GID>1580</GID>
<name>IN_0</name></connection>
<intersection>-4997.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-4989.5,204,-4989.5</points>
<connection>
<GID>1584</GID>
<name>OUT</name></connection>
<connection>
<GID>1583</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-4998,185.5,-4979</points>
<intersection>-4998 3</intersection>
<intersection>-4988.5 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,-4988.5,188.5,-4988.5</points>
<connection>
<GID>1584</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-4979,185.5,-4979</points>
<connection>
<GID>1582</GID>
<name>OUT_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185.5,-4998,206,-4998</points>
<intersection>185.5 0</intersection>
<intersection>206 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>206,-4998,206,-4992.5</points>
<connection>
<GID>1583</GID>
<name>IN_0</name></connection>
<intersection>-4998 3</intersection></vsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>268.5,-4989.5,277.5,-4989.5</points>
<connection>
<GID>1581</GID>
<name>OUT</name></connection>
<connection>
<GID>1586</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-4999.5,259,-4979</points>
<connection>
<GID>1585</GID>
<name>OUT_0</name></connection>
<intersection>-4999.5 3</intersection>
<intersection>-4988.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259,-4988.5,262.5,-4988.5</points>
<connection>
<GID>1581</GID>
<name>IN_0</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259,-4999.5,279.5,-4999.5</points>
<intersection>259 0</intersection>
<intersection>279.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>279.5,-4999.5,279.5,-4992.5</points>
<connection>
<GID>1586</GID>
<name>IN_0</name></connection>
<intersection>-4999.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359.5,-4991,369,-4991</points>
<connection>
<GID>1590</GID>
<name>OUT</name></connection>
<connection>
<GID>1589</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350.5,-4999.5,350.5,-4979</points>
<intersection>-4999.5 3</intersection>
<intersection>-4990 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350.5,-4990,353.5,-4990</points>
<connection>
<GID>1590</GID>
<name>IN_0</name></connection>
<intersection>350.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-4979,350.5,-4979</points>
<connection>
<GID>1588</GID>
<name>OUT_0</name></connection>
<intersection>350.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>350.5,-4999.5,371,-4999.5</points>
<intersection>350.5 0</intersection>
<intersection>371 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>371,-4999.5,371,-4994</points>
<connection>
<GID>1589</GID>
<name>IN_0</name></connection>
<intersection>-4999.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>433.5,-4991,442.5,-4991</points>
<connection>
<GID>1587</GID>
<name>OUT</name></connection>
<connection>
<GID>1592</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424,-4999.5,424,-4979</points>
<intersection>-4999.5 3</intersection>
<intersection>-4990 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424,-4990,427.5,-4990</points>
<connection>
<GID>1587</GID>
<name>IN_0</name></connection>
<intersection>424 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423,-4979,424,-4979</points>
<connection>
<GID>1591</GID>
<name>OUT_0</name></connection>
<intersection>424 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>424,-4999.5,444.5,-4999.5</points>
<intersection>424 0</intersection>
<intersection>444.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>444.5,-4999.5,444.5,-4994</points>
<connection>
<GID>1592</GID>
<name>IN_0</name></connection>
<intersection>-4999.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>517.5,-4993,527,-4993</points>
<connection>
<GID>1596</GID>
<name>OUT</name></connection>
<connection>
<GID>1595</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508.5,-4999,508.5,-4979</points>
<intersection>-4999 3</intersection>
<intersection>-4992 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508.5,-4992,511.5,-4992</points>
<connection>
<GID>1596</GID>
<name>IN_0</name></connection>
<intersection>508.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507.5,-4979,508.5,-4979</points>
<connection>
<GID>1594</GID>
<name>OUT_0</name></connection>
<intersection>508.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>508.5,-4999,529,-4999</points>
<intersection>508.5 0</intersection>
<intersection>529 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>529,-4999,529,-4996</points>
<connection>
<GID>1595</GID>
<name>IN_0</name></connection>
<intersection>-4999 3</intersection></vsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>591.5,-4993,600.5,-4993</points>
<connection>
<GID>1593</GID>
<name>OUT</name></connection>
<connection>
<GID>1598</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>582,-4999,582,-4979</points>
<intersection>-4999 3</intersection>
<intersection>-4992 1</intersection>
<intersection>-4979 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>582,-4992,585.5,-4992</points>
<connection>
<GID>1593</GID>
<name>IN_0</name></connection>
<intersection>582 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>581,-4979,582,-4979</points>
<connection>
<GID>1597</GID>
<name>OUT_0</name></connection>
<intersection>582 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>582,-4999,602.5,-4999</points>
<intersection>582 0</intersection>
<intersection>602.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>602.5,-4999,602.5,-4996</points>
<connection>
<GID>1598</GID>
<name>IN_0</name></connection>
<intersection>-4999 3</intersection></vsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-4982,575,-4982</points>
<connection>
<GID>1576</GID>
<name>clock</name></connection>
<connection>
<GID>1579</GID>
<name>clock</name></connection>
<connection>
<GID>1582</GID>
<name>clock</name></connection>
<connection>
<GID>1585</GID>
<name>clock</name></connection>
<connection>
<GID>1591</GID>
<name>clock</name></connection>
<connection>
<GID>1594</GID>
<name>clock</name></connection>
<connection>
<GID>1597</GID>
<name>clock</name></connection>
<connection>
<GID>1599</GID>
<name>OUT</name></connection>
<connection>
<GID>1588</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113.5,-5223,-113.5,-4891</points>
<intersection>-5223 2</intersection>
<intersection>-4909 3</intersection>
<intersection>-4891 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-113.5,-4891,-14,-4891</points>
<connection>
<GID>1625</GID>
<name>IN_0</name></connection>
<intersection>-113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5223,-113.5,-5223</points>
<connection>
<GID>1574</GID>
<name>OUT_7</name></connection>
<intersection>-113.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-113.5,-4909,-32.5,-4909</points>
<connection>
<GID>1626</GID>
<name>ENABLE_0</name></connection>
<intersection>-113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-30,-4911,582.5,-4911</points>
<connection>
<GID>1626</GID>
<name>OUT_0</name></connection>
<intersection>27.5 38</intersection>
<intersection>101.5 43</intersection>
<intersection>185.5 42</intersection>
<intersection>259.5 45</intersection>
<intersection>350.5 47</intersection>
<intersection>424.5 49</intersection>
<intersection>508.5 51</intersection>
<intersection>582.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>27.5,-4911,27.5,-4898.5</points>
<connection>
<GID>1604</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>185.5,-4911,185.5,-4900.5</points>
<connection>
<GID>1610</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>101.5,-4911,101.5,-4898.5</points>
<connection>
<GID>1601</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>259.5,-4911,259.5,-4900.5</points>
<connection>
<GID>1607</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>350.5,-4911,350.5,-4902</points>
<connection>
<GID>1616</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>424.5,-4911,424.5,-4902</points>
<connection>
<GID>1613</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>508.5,-4911,508.5,-4904</points>
<connection>
<GID>1622</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>582.5,-4911,582.5,-4904</points>
<connection>
<GID>1619</GID>
<name>IN_1</name></connection>
<intersection>-4911 33</intersection></vsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-4897.5,43,-4897.5</points>
<connection>
<GID>1604</GID>
<name>OUT</name></connection>
<connection>
<GID>1603</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-4906,24.5,-4889</points>
<intersection>-4906 3</intersection>
<intersection>-4896.5 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-4896.5,27.5,-4896.5</points>
<connection>
<GID>1604</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-4889,24.5,-4889</points>
<connection>
<GID>1602</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-4906,45,-4906</points>
<intersection>24.5 0</intersection>
<intersection>45 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45,-4906,45,-4900.5</points>
<connection>
<GID>1603</GID>
<name>IN_0</name></connection>
<intersection>-4906 3</intersection></vsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>107.5,-4897.5,116.5,-4897.5</points>
<connection>
<GID>1601</GID>
<name>OUT</name></connection>
<connection>
<GID>1606</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-4907.5,98,-4889</points>
<intersection>-4907.5 3</intersection>
<intersection>-4896.5 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-4896.5,101.5,-4896.5</points>
<connection>
<GID>1601</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-4889,98,-4889</points>
<connection>
<GID>1605</GID>
<name>OUT_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>98,-4907.5,118.5,-4907.5</points>
<intersection>98 0</intersection>
<intersection>118.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>118.5,-4907.5,118.5,-4900.5</points>
<connection>
<GID>1606</GID>
<name>IN_0</name></connection>
<intersection>-4907.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191.5,-4899.5,201,-4899.5</points>
<connection>
<GID>1610</GID>
<name>OUT</name></connection>
<connection>
<GID>1609</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-4908,182.5,-4889</points>
<intersection>-4908 3</intersection>
<intersection>-4898.5 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>182.5,-4898.5,185.5,-4898.5</points>
<connection>
<GID>1610</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-4889,182.5,-4889</points>
<connection>
<GID>1608</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>182.5,-4908,203,-4908</points>
<intersection>182.5 0</intersection>
<intersection>203 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>203,-4908,203,-4902.5</points>
<connection>
<GID>1609</GID>
<name>IN_0</name></connection>
<intersection>-4908 3</intersection></vsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>265.5,-4899.5,274.5,-4899.5</points>
<connection>
<GID>1607</GID>
<name>OUT</name></connection>
<connection>
<GID>1612</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,-4909.5,256,-4889</points>
<connection>
<GID>1611</GID>
<name>OUT_0</name></connection>
<intersection>-4909.5 3</intersection>
<intersection>-4898.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,-4898.5,259.5,-4898.5</points>
<connection>
<GID>1607</GID>
<name>IN_0</name></connection>
<intersection>256 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>256,-4909.5,276.5,-4909.5</points>
<intersection>256 0</intersection>
<intersection>276.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>276.5,-4909.5,276.5,-4902.5</points>
<connection>
<GID>1612</GID>
<name>IN_0</name></connection>
<intersection>-4909.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>356.5,-4901,366,-4901</points>
<connection>
<GID>1616</GID>
<name>OUT</name></connection>
<connection>
<GID>1615</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347.5,-4909.5,347.5,-4889</points>
<intersection>-4909.5 3</intersection>
<intersection>-4900 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347.5,-4900,350.5,-4900</points>
<connection>
<GID>1616</GID>
<name>IN_0</name></connection>
<intersection>347.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346.5,-4889,347.5,-4889</points>
<connection>
<GID>1614</GID>
<name>OUT_0</name></connection>
<intersection>347.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>347.5,-4909.5,368,-4909.5</points>
<intersection>347.5 0</intersection>
<intersection>368 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>368,-4909.5,368,-4904</points>
<connection>
<GID>1615</GID>
<name>IN_0</name></connection>
<intersection>-4909.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>430.5,-4901,439.5,-4901</points>
<connection>
<GID>1613</GID>
<name>OUT</name></connection>
<connection>
<GID>1618</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421,-4909.5,421,-4889</points>
<intersection>-4909.5 3</intersection>
<intersection>-4900 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>421,-4900,424.5,-4900</points>
<connection>
<GID>1613</GID>
<name>IN_0</name></connection>
<intersection>421 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>420,-4889,421,-4889</points>
<connection>
<GID>1617</GID>
<name>OUT_0</name></connection>
<intersection>421 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>421,-4909.5,441.5,-4909.5</points>
<intersection>421 0</intersection>
<intersection>441.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>441.5,-4909.5,441.5,-4904</points>
<connection>
<GID>1618</GID>
<name>IN_0</name></connection>
<intersection>-4909.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>514.5,-4903,524,-4903</points>
<connection>
<GID>1622</GID>
<name>OUT</name></connection>
<connection>
<GID>1621</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,-4909,505.5,-4889</points>
<intersection>-4909 3</intersection>
<intersection>-4902 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505.5,-4902,508.5,-4902</points>
<connection>
<GID>1622</GID>
<name>IN_0</name></connection>
<intersection>505.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>504.5,-4889,505.5,-4889</points>
<connection>
<GID>1620</GID>
<name>OUT_0</name></connection>
<intersection>505.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>505.5,-4909,526,-4909</points>
<intersection>505.5 0</intersection>
<intersection>526 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>526,-4909,526,-4906</points>
<connection>
<GID>1621</GID>
<name>IN_0</name></connection>
<intersection>-4909 3</intersection></vsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>588.5,-4903,597.5,-4903</points>
<connection>
<GID>1619</GID>
<name>OUT</name></connection>
<connection>
<GID>1624</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579,-4909,579,-4889</points>
<intersection>-4909 3</intersection>
<intersection>-4902 1</intersection>
<intersection>-4889 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>579,-4902,582.5,-4902</points>
<connection>
<GID>1619</GID>
<name>IN_0</name></connection>
<intersection>579 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>578,-4889,579,-4889</points>
<connection>
<GID>1623</GID>
<name>OUT_0</name></connection>
<intersection>579 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>579,-4909,599.5,-4909</points>
<intersection>579 0</intersection>
<intersection>599.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>599.5,-4909,599.5,-4906</points>
<connection>
<GID>1624</GID>
<name>IN_0</name></connection>
<intersection>-4909 3</intersection></vsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-4892,572,-4892</points>
<connection>
<GID>1625</GID>
<name>OUT</name></connection>
<connection>
<GID>1623</GID>
<name>clock</name></connection>
<connection>
<GID>1620</GID>
<name>clock</name></connection>
<connection>
<GID>1617</GID>
<name>clock</name></connection>
<connection>
<GID>1614</GID>
<name>clock</name></connection>
<connection>
<GID>1611</GID>
<name>clock</name></connection>
<connection>
<GID>1608</GID>
<name>clock</name></connection>
<connection>
<GID>1605</GID>
<name>clock</name></connection>
<connection>
<GID>1602</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110.5,-5226,-110.5,-5149</points>
<intersection>-5226 2</intersection>
<intersection>-5167 3</intersection>
<intersection>-5149 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-5149,-7,-5149</points>
<connection>
<GID>1651</GID>
<name>IN_0</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5226,-110.5,-5226</points>
<connection>
<GID>1574</GID>
<name>OUT_4</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110.5,-5167,-25.5,-5167</points>
<connection>
<GID>1652</GID>
<name>ENABLE_0</name></connection>
<intersection>-110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23,-5169,589.5,-5169</points>
<connection>
<GID>1652</GID>
<name>OUT_0</name></connection>
<intersection>34.5 38</intersection>
<intersection>108.5 43</intersection>
<intersection>192.5 42</intersection>
<intersection>266.5 45</intersection>
<intersection>357.5 47</intersection>
<intersection>431.5 49</intersection>
<intersection>515.5 51</intersection>
<intersection>589.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34.5,-5169,34.5,-5156.5</points>
<connection>
<GID>1630</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192.5,-5169,192.5,-5158.5</points>
<connection>
<GID>1636</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108.5,-5169,108.5,-5156.5</points>
<connection>
<GID>1627</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266.5,-5169,266.5,-5158.5</points>
<connection>
<GID>1633</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357.5,-5169,357.5,-5160</points>
<connection>
<GID>1642</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431.5,-5169,431.5,-5160</points>
<connection>
<GID>1639</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515.5,-5169,515.5,-5162</points>
<connection>
<GID>1648</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589.5,-5169,589.5,-5162</points>
<connection>
<GID>1645</GID>
<name>IN_1</name></connection>
<intersection>-5169 33</intersection></vsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-5155.5,50,-5155.5</points>
<connection>
<GID>1630</GID>
<name>OUT</name></connection>
<connection>
<GID>1629</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-5164,31.5,-5147</points>
<intersection>-5164 3</intersection>
<intersection>-5154.5 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-5154.5,34.5,-5154.5</points>
<connection>
<GID>1630</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-5147,31.5,-5147</points>
<connection>
<GID>1628</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-5164,52,-5164</points>
<intersection>31.5 0</intersection>
<intersection>52 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52,-5164,52,-5158.5</points>
<connection>
<GID>1629</GID>
<name>IN_0</name></connection>
<intersection>-5164 3</intersection></vsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114.5,-5155.5,123.5,-5155.5</points>
<connection>
<GID>1627</GID>
<name>OUT</name></connection>
<connection>
<GID>1632</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-5165.5,105,-5147</points>
<intersection>-5165.5 3</intersection>
<intersection>-5154.5 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-5154.5,108.5,-5154.5</points>
<connection>
<GID>1627</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-5147,105,-5147</points>
<connection>
<GID>1631</GID>
<name>OUT_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105,-5165.5,125.5,-5165.5</points>
<intersection>105 0</intersection>
<intersection>125.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125.5,-5165.5,125.5,-5158.5</points>
<connection>
<GID>1632</GID>
<name>IN_0</name></connection>
<intersection>-5165.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198.5,-5157.5,208,-5157.5</points>
<connection>
<GID>1636</GID>
<name>OUT</name></connection>
<connection>
<GID>1635</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-5166,189.5,-5147</points>
<intersection>-5166 3</intersection>
<intersection>-5156.5 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,-5156.5,192.5,-5156.5</points>
<connection>
<GID>1636</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,-5147,189.5,-5147</points>
<connection>
<GID>1634</GID>
<name>OUT_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189.5,-5166,210,-5166</points>
<intersection>189.5 0</intersection>
<intersection>210 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>210,-5166,210,-5160.5</points>
<connection>
<GID>1635</GID>
<name>IN_0</name></connection>
<intersection>-5166 3</intersection></vsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272.5,-5157.5,281.5,-5157.5</points>
<connection>
<GID>1633</GID>
<name>OUT</name></connection>
<connection>
<GID>1638</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-5167.5,263,-5147</points>
<connection>
<GID>1637</GID>
<name>OUT_0</name></connection>
<intersection>-5167.5 3</intersection>
<intersection>-5156.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-5156.5,266.5,-5156.5</points>
<connection>
<GID>1633</GID>
<name>IN_0</name></connection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>263,-5167.5,283.5,-5167.5</points>
<intersection>263 0</intersection>
<intersection>283.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283.5,-5167.5,283.5,-5160.5</points>
<connection>
<GID>1638</GID>
<name>IN_0</name></connection>
<intersection>-5167.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363.5,-5159,373,-5159</points>
<connection>
<GID>1642</GID>
<name>OUT</name></connection>
<connection>
<GID>1641</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-5167.5,354.5,-5147</points>
<intersection>-5167.5 3</intersection>
<intersection>-5158 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354.5,-5158,357.5,-5158</points>
<connection>
<GID>1642</GID>
<name>IN_0</name></connection>
<intersection>354.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353.5,-5147,354.5,-5147</points>
<connection>
<GID>1640</GID>
<name>OUT_0</name></connection>
<intersection>354.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354.5,-5167.5,375,-5167.5</points>
<intersection>354.5 0</intersection>
<intersection>375 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>375,-5167.5,375,-5162</points>
<connection>
<GID>1641</GID>
<name>IN_0</name></connection>
<intersection>-5167.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437.5,-5159,446.5,-5159</points>
<connection>
<GID>1639</GID>
<name>OUT</name></connection>
<connection>
<GID>1644</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,-5167.5,428,-5147</points>
<intersection>-5167.5 3</intersection>
<intersection>-5158 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428,-5158,431.5,-5158</points>
<connection>
<GID>1639</GID>
<name>IN_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427,-5147,428,-5147</points>
<connection>
<GID>1643</GID>
<name>OUT_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428,-5167.5,448.5,-5167.5</points>
<intersection>428 0</intersection>
<intersection>448.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448.5,-5167.5,448.5,-5162</points>
<connection>
<GID>1644</GID>
<name>IN_0</name></connection>
<intersection>-5167.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521.5,-5161,531,-5161</points>
<connection>
<GID>1648</GID>
<name>OUT</name></connection>
<connection>
<GID>1647</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512.5,-5167,512.5,-5147</points>
<intersection>-5167 3</intersection>
<intersection>-5160 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512.5,-5160,515.5,-5160</points>
<connection>
<GID>1648</GID>
<name>IN_0</name></connection>
<intersection>512.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511.5,-5147,512.5,-5147</points>
<connection>
<GID>1646</GID>
<name>OUT_0</name></connection>
<intersection>512.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512.5,-5167,533,-5167</points>
<intersection>512.5 0</intersection>
<intersection>533 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>533,-5167,533,-5164</points>
<connection>
<GID>1647</GID>
<name>IN_0</name></connection>
<intersection>-5167 3</intersection></vsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595.5,-5161,604.5,-5161</points>
<connection>
<GID>1645</GID>
<name>OUT</name></connection>
<connection>
<GID>1650</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586,-5167,586,-5147</points>
<intersection>-5167 3</intersection>
<intersection>-5160 1</intersection>
<intersection>-5147 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>586,-5160,589.5,-5160</points>
<connection>
<GID>1645</GID>
<name>IN_0</name></connection>
<intersection>586 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585,-5147,586,-5147</points>
<connection>
<GID>1649</GID>
<name>OUT_0</name></connection>
<intersection>586 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>586,-5167,606.5,-5167</points>
<intersection>586 0</intersection>
<intersection>606.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606.5,-5167,606.5,-5164</points>
<connection>
<GID>1650</GID>
<name>IN_0</name></connection>
<intersection>-5167 3</intersection></vsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-5150,579,-5150</points>
<connection>
<GID>1628</GID>
<name>clock</name></connection>
<connection>
<GID>1631</GID>
<name>clock</name></connection>
<connection>
<GID>1634</GID>
<name>clock</name></connection>
<connection>
<GID>1637</GID>
<name>clock</name></connection>
<connection>
<GID>1640</GID>
<name>clock</name></connection>
<connection>
<GID>1643</GID>
<name>clock</name></connection>
<connection>
<GID>1646</GID>
<name>clock</name></connection>
<connection>
<GID>1651</GID>
<name>OUT</name></connection>
<connection>
<GID>1649</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111.5,-5225,-111.5,-5059</points>
<intersection>-5225 2</intersection>
<intersection>-5077 3</intersection>
<intersection>-5059 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111.5,-5059,-10,-5059</points>
<connection>
<GID>1677</GID>
<name>IN_0</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5225,-111.5,-5225</points>
<connection>
<GID>1574</GID>
<name>OUT_5</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111.5,-5077,-28.5,-5077</points>
<connection>
<GID>1678</GID>
<name>ENABLE_0</name></connection>
<intersection>-111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-26,-5079,586.5,-5079</points>
<connection>
<GID>1678</GID>
<name>OUT_0</name></connection>
<intersection>29 54</intersection>
<intersection>105.5 43</intersection>
<intersection>189.5 42</intersection>
<intersection>263.5 45</intersection>
<intersection>354.5 47</intersection>
<intersection>428.5 49</intersection>
<intersection>512.5 51</intersection>
<intersection>586.5 53</intersection></hsegment>
<vsegment>
<ID>42</ID>
<points>189.5,-5079,189.5,-5068.5</points>
<connection>
<GID>1662</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>105.5,-5079,105.5,-5066.5</points>
<connection>
<GID>1653</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>263.5,-5079,263.5,-5068.5</points>
<connection>
<GID>1659</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>354.5,-5079,354.5,-5070</points>
<connection>
<GID>1668</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>428.5,-5079,428.5,-5070</points>
<connection>
<GID>1665</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>512.5,-5079,512.5,-5072</points>
<connection>
<GID>1674</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>586.5,-5079,586.5,-5072</points>
<connection>
<GID>1671</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>29,-5079,29,-5067</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>-5079 33</intersection></vsegment></shape></wire>
<wire>
<ID>1142</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>111.5,-5065.5,120.5,-5065.5</points>
<connection>
<GID>1653</GID>
<name>OUT</name></connection>
<connection>
<GID>1658</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-5075.5,102,-5057</points>
<intersection>-5075.5 3</intersection>
<intersection>-5064.5 1</intersection>
<intersection>-5057 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-5064.5,105.5,-5064.5</points>
<connection>
<GID>1653</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-5057,102,-5057</points>
<connection>
<GID>1657</GID>
<name>OUT_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,-5075.5,122.5,-5075.5</points>
<intersection>102 0</intersection>
<intersection>122.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122.5,-5075.5,122.5,-5068.5</points>
<connection>
<GID>1658</GID>
<name>IN_0</name></connection>
<intersection>-5075.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195.5,-5067.5,205,-5067.5</points>
<connection>
<GID>1662</GID>
<name>OUT</name></connection>
<connection>
<GID>1661</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-5076,186.5,-5057</points>
<intersection>-5076 3</intersection>
<intersection>-5066.5 1</intersection>
<intersection>-5057 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,-5066.5,189.5,-5066.5</points>
<connection>
<GID>1662</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185.5,-5057,186.5,-5057</points>
<connection>
<GID>1660</GID>
<name>OUT_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>186.5,-5076,207,-5076</points>
<intersection>186.5 0</intersection>
<intersection>207 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207,-5076,207,-5070.5</points>
<connection>
<GID>1661</GID>
<name>IN_0</name></connection>
<intersection>-5076 3</intersection></vsegment></shape></wire>
<wire>
<ID>1146</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>269.5,-5067.5,278.5,-5067.5</points>
<connection>
<GID>1659</GID>
<name>OUT</name></connection>
<connection>
<GID>1664</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-5077.5,260,-5057</points>
<connection>
<GID>1663</GID>
<name>OUT_0</name></connection>
<intersection>-5077.5 3</intersection>
<intersection>-5066.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-5066.5,263.5,-5066.5</points>
<connection>
<GID>1659</GID>
<name>IN_0</name></connection>
<intersection>260 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260,-5077.5,280.5,-5077.5</points>
<intersection>260 0</intersection>
<intersection>280.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>280.5,-5077.5,280.5,-5070.5</points>
<connection>
<GID>1664</GID>
<name>IN_0</name></connection>
<intersection>-5077.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360.5,-5069,370,-5069</points>
<connection>
<GID>1668</GID>
<name>OUT</name></connection>
<connection>
<GID>1667</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,-5077.5,351.5,-5057</points>
<intersection>-5077.5 3</intersection>
<intersection>-5068 1</intersection>
<intersection>-5057 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,-5068,354.5,-5068</points>
<connection>
<GID>1668</GID>
<name>IN_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350.5,-5057,351.5,-5057</points>
<connection>
<GID>1666</GID>
<name>OUT_0</name></connection>
<intersection>351.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>351.5,-5077.5,372,-5077.5</points>
<intersection>351.5 0</intersection>
<intersection>372 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372,-5077.5,372,-5072</points>
<connection>
<GID>1667</GID>
<name>IN_0</name></connection>
<intersection>-5077.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1150</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>434.5,-5069,443.5,-5069</points>
<connection>
<GID>1665</GID>
<name>OUT</name></connection>
<connection>
<GID>1670</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425,-5077.5,425,-5057</points>
<intersection>-5077.5 3</intersection>
<intersection>-5068 1</intersection>
<intersection>-5057 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425,-5068,428.5,-5068</points>
<connection>
<GID>1665</GID>
<name>IN_0</name></connection>
<intersection>425 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424,-5057,425,-5057</points>
<connection>
<GID>1669</GID>
<name>OUT_0</name></connection>
<intersection>425 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425,-5077.5,445.5,-5077.5</points>
<intersection>425 0</intersection>
<intersection>445.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>445.5,-5077.5,445.5,-5072</points>
<connection>
<GID>1670</GID>
<name>IN_0</name></connection>
<intersection>-5077.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509.5,-5077,509.5,-5057</points>
<intersection>-5077 3</intersection>
<intersection>-5070 1</intersection>
<intersection>-5057 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,-5070,512.5,-5070</points>
<connection>
<GID>1674</GID>
<name>IN_0</name></connection>
<intersection>509.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>508.5,-5057,509.5,-5057</points>
<connection>
<GID>1672</GID>
<name>OUT_0</name></connection>
<intersection>509.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>509.5,-5077,530,-5077</points>
<intersection>509.5 0</intersection>
<intersection>530 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530,-5077,530,-5074</points>
<connection>
<GID>1673</GID>
<name>IN_0</name></connection>
<intersection>-5077 3</intersection></vsegment></shape></wire>
<wire>
<ID>1154</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>592.5,-5071,601.5,-5071</points>
<connection>
<GID>1671</GID>
<name>OUT</name></connection>
<connection>
<GID>1676</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583,-5077,583,-5057</points>
<intersection>-5077 3</intersection>
<intersection>-5070 1</intersection>
<intersection>-5057 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583,-5070,586.5,-5070</points>
<connection>
<GID>1671</GID>
<name>IN_0</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582,-5057,583,-5057</points>
<connection>
<GID>1675</GID>
<name>OUT_0</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583,-5077,603.5,-5077</points>
<intersection>583 0</intersection>
<intersection>603.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>603.5,-5077,603.5,-5074</points>
<connection>
<GID>1676</GID>
<name>IN_0</name></connection>
<intersection>-5077 3</intersection></vsegment></shape></wire>
<wire>
<ID>1156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-5060,576,-5060</points>
<connection>
<GID>1677</GID>
<name>OUT</name></connection>
<connection>
<GID>1675</GID>
<name>clock</name></connection>
<connection>
<GID>1672</GID>
<name>clock</name></connection>
<connection>
<GID>1669</GID>
<name>clock</name></connection>
<connection>
<GID>1666</GID>
<name>clock</name></connection>
<connection>
<GID>1663</GID>
<name>clock</name></connection>
<connection>
<GID>1660</GID>
<name>clock</name></connection>
<connection>
<GID>1657</GID>
<name>clock</name></connection>
<connection>
<GID>1654</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111.5,-5375,-111.5,-5228</points>
<intersection>-5375 3</intersection>
<intersection>-5357 1</intersection>
<intersection>-5228 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111.5,-5357,-9,-5357</points>
<connection>
<GID>1703</GID>
<name>IN_0</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5228,-111.5,-5228</points>
<connection>
<GID>1574</GID>
<name>OUT_2</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111.5,-5375,-27.5,-5375</points>
<connection>
<GID>1704</GID>
<name>ENABLE_0</name></connection>
<intersection>-111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1158</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25,-5377,587.5,-5377</points>
<connection>
<GID>1704</GID>
<name>OUT_0</name></connection>
<intersection>32.5 38</intersection>
<intersection>106.5 43</intersection>
<intersection>190.5 42</intersection>
<intersection>264.5 45</intersection>
<intersection>355.5 47</intersection>
<intersection>429.5 49</intersection>
<intersection>513.5 51</intersection>
<intersection>587.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32.5,-5377,32.5,-5364.5</points>
<connection>
<GID>1682</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190.5,-5377,190.5,-5366.5</points>
<connection>
<GID>1688</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106.5,-5377,106.5,-5364.5</points>
<connection>
<GID>1679</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264.5,-5377,264.5,-5366.5</points>
<connection>
<GID>1685</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355.5,-5377,355.5,-5368</points>
<connection>
<GID>1694</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429.5,-5377,429.5,-5368</points>
<connection>
<GID>1691</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513.5,-5377,513.5,-5370</points>
<connection>
<GID>1700</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587.5,-5377,587.5,-5370</points>
<connection>
<GID>1697</GID>
<name>IN_1</name></connection>
<intersection>-5377 33</intersection></vsegment></shape></wire>
<wire>
<ID>1159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-5363.5,48,-5363.5</points>
<connection>
<GID>1682</GID>
<name>OUT</name></connection>
<connection>
<GID>1681</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-5372,29.5,-5355</points>
<intersection>-5372 3</intersection>
<intersection>-5362.5 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-5362.5,32.5,-5362.5</points>
<connection>
<GID>1682</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-5355,29.5,-5355</points>
<connection>
<GID>1680</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-5372,50,-5372</points>
<intersection>29.5 0</intersection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,-5372,50,-5366.5</points>
<connection>
<GID>1681</GID>
<name>IN_0</name></connection>
<intersection>-5372 3</intersection></vsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112.5,-5363.5,121.5,-5363.5</points>
<connection>
<GID>1679</GID>
<name>OUT</name></connection>
<connection>
<GID>1684</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-5373.5,103,-5355</points>
<intersection>-5373.5 3</intersection>
<intersection>-5362.5 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-5362.5,106.5,-5362.5</points>
<connection>
<GID>1679</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-5355,103,-5355</points>
<connection>
<GID>1683</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,-5373.5,123.5,-5373.5</points>
<intersection>103 0</intersection>
<intersection>123.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123.5,-5373.5,123.5,-5366.5</points>
<connection>
<GID>1684</GID>
<name>IN_0</name></connection>
<intersection>-5373.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,-5365.5,206,-5365.5</points>
<connection>
<GID>1688</GID>
<name>OUT</name></connection>
<connection>
<GID>1687</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-5374,187.5,-5355</points>
<intersection>-5374 3</intersection>
<intersection>-5364.5 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,-5364.5,190.5,-5364.5</points>
<connection>
<GID>1688</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186.5,-5355,187.5,-5355</points>
<connection>
<GID>1686</GID>
<name>OUT_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-5374,208,-5374</points>
<intersection>187.5 0</intersection>
<intersection>208 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208,-5374,208,-5368.5</points>
<connection>
<GID>1687</GID>
<name>IN_0</name></connection>
<intersection>-5374 3</intersection></vsegment></shape></wire>
<wire>
<ID>1165</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270.5,-5365.5,279.5,-5365.5</points>
<connection>
<GID>1685</GID>
<name>OUT</name></connection>
<connection>
<GID>1690</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-5375.5,261,-5355</points>
<connection>
<GID>1689</GID>
<name>OUT_0</name></connection>
<intersection>-5375.5 3</intersection>
<intersection>-5364.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-5364.5,264.5,-5364.5</points>
<connection>
<GID>1685</GID>
<name>IN_0</name></connection>
<intersection>261 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>261,-5375.5,281.5,-5375.5</points>
<intersection>261 0</intersection>
<intersection>281.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281.5,-5375.5,281.5,-5368.5</points>
<connection>
<GID>1690</GID>
<name>IN_0</name></connection>
<intersection>-5375.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361.5,-5367,371,-5367</points>
<connection>
<GID>1694</GID>
<name>OUT</name></connection>
<connection>
<GID>1693</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352.5,-5375.5,352.5,-5355</points>
<intersection>-5375.5 3</intersection>
<intersection>-5366 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352.5,-5366,355.5,-5366</points>
<connection>
<GID>1694</GID>
<name>IN_0</name></connection>
<intersection>352.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351.5,-5355,352.5,-5355</points>
<connection>
<GID>1692</GID>
<name>OUT_0</name></connection>
<intersection>352.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352.5,-5375.5,373,-5375.5</points>
<intersection>352.5 0</intersection>
<intersection>373 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>373,-5375.5,373,-5370</points>
<connection>
<GID>1693</GID>
<name>IN_0</name></connection>
<intersection>-5375.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1169</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435.5,-5367,444.5,-5367</points>
<connection>
<GID>1691</GID>
<name>OUT</name></connection>
<connection>
<GID>1696</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,-5375.5,426,-5355</points>
<intersection>-5375.5 3</intersection>
<intersection>-5366 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426,-5366,429.5,-5366</points>
<connection>
<GID>1691</GID>
<name>IN_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425,-5355,426,-5355</points>
<connection>
<GID>1695</GID>
<name>OUT_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426,-5375.5,446.5,-5375.5</points>
<intersection>426 0</intersection>
<intersection>446.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446.5,-5375.5,446.5,-5370</points>
<connection>
<GID>1696</GID>
<name>IN_0</name></connection>
<intersection>-5375.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519.5,-5369,529,-5369</points>
<connection>
<GID>1700</GID>
<name>OUT</name></connection>
<connection>
<GID>1699</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510.5,-5375,510.5,-5355</points>
<intersection>-5375 3</intersection>
<intersection>-5368 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,-5368,513.5,-5368</points>
<connection>
<GID>1700</GID>
<name>IN_0</name></connection>
<intersection>510.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509.5,-5355,510.5,-5355</points>
<connection>
<GID>1698</GID>
<name>OUT_0</name></connection>
<intersection>510.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510.5,-5375,531,-5375</points>
<intersection>510.5 0</intersection>
<intersection>531 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531,-5375,531,-5372</points>
<connection>
<GID>1699</GID>
<name>IN_0</name></connection>
<intersection>-5375 3</intersection></vsegment></shape></wire>
<wire>
<ID>1173</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593.5,-5369,602.5,-5369</points>
<connection>
<GID>1697</GID>
<name>OUT</name></connection>
<connection>
<GID>1702</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584,-5375,584,-5355</points>
<intersection>-5375 3</intersection>
<intersection>-5368 1</intersection>
<intersection>-5355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584,-5368,587.5,-5368</points>
<connection>
<GID>1697</GID>
<name>IN_0</name></connection>
<intersection>584 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583,-5355,584,-5355</points>
<connection>
<GID>1701</GID>
<name>OUT_0</name></connection>
<intersection>584 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>584,-5375,604.5,-5375</points>
<intersection>584 0</intersection>
<intersection>604.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604.5,-5375,604.5,-5372</points>
<connection>
<GID>1702</GID>
<name>IN_0</name></connection>
<intersection>-5375 3</intersection></vsegment></shape></wire>
<wire>
<ID>1175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3,-5358,577,-5358</points>
<connection>
<GID>1703</GID>
<name>OUT</name></connection>
<connection>
<GID>1701</GID>
<name>clock</name></connection>
<connection>
<GID>1698</GID>
<name>clock</name></connection>
<connection>
<GID>1695</GID>
<name>clock</name></connection>
<connection>
<GID>1692</GID>
<name>clock</name></connection>
<connection>
<GID>1689</GID>
<name>clock</name></connection>
<connection>
<GID>1686</GID>
<name>clock</name></connection>
<connection>
<GID>1683</GID>
<name>clock</name></connection>
<connection>
<GID>1680</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110.5,-5285,-110.5,-5227</points>
<intersection>-5285 3</intersection>
<intersection>-5267 1</intersection>
<intersection>-5227 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-110.5,-5267,-12,-5267</points>
<connection>
<GID>1520</GID>
<name>IN_0</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5227,-110.5,-5227</points>
<connection>
<GID>1574</GID>
<name>OUT_3</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110.5,-5285,-30.5,-5285</points>
<connection>
<GID>1521</GID>
<name>ENABLE_0</name></connection>
<intersection>-110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1177</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-28,-5287,584.5,-5287</points>
<connection>
<GID>1521</GID>
<name>OUT_0</name></connection>
<intersection>29.5 38</intersection>
<intersection>103.5 43</intersection>
<intersection>187.5 42</intersection>
<intersection>261.5 45</intersection>
<intersection>352.5 47</intersection>
<intersection>426.5 49</intersection>
<intersection>510.5 51</intersection>
<intersection>584.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>29.5,-5287,29.5,-5274.5</points>
<connection>
<GID>1708</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>187.5,-5287,187.5,-5276.5</points>
<connection>
<GID>1505</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>103.5,-5287,103.5,-5274.5</points>
<connection>
<GID>1705</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>261.5,-5287,261.5,-5276.5</points>
<connection>
<GID>1711</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>352.5,-5287,352.5,-5278</points>
<connection>
<GID>1511</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>426.5,-5287,426.5,-5278</points>
<connection>
<GID>1508</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>510.5,-5287,510.5,-5280</points>
<connection>
<GID>1517</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>584.5,-5287,584.5,-5280</points>
<connection>
<GID>1514</GID>
<name>IN_1</name></connection>
<intersection>-5287 33</intersection></vsegment></shape></wire>
<wire>
<ID>1178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-5273.5,45,-5273.5</points>
<connection>
<GID>1708</GID>
<name>OUT</name></connection>
<connection>
<GID>1707</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-5282,26.5,-5265</points>
<intersection>-5282 3</intersection>
<intersection>-5272.5 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-5272.5,29.5,-5272.5</points>
<connection>
<GID>1708</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-5265,26.5,-5265</points>
<connection>
<GID>1706</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-5282,47,-5282</points>
<intersection>26.5 0</intersection>
<intersection>47 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>47,-5282,47,-5276.5</points>
<connection>
<GID>1707</GID>
<name>IN_0</name></connection>
<intersection>-5282 3</intersection></vsegment></shape></wire>
<wire>
<ID>1180</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>109.5,-5273.5,118.5,-5273.5</points>
<connection>
<GID>1705</GID>
<name>OUT</name></connection>
<connection>
<GID>1710</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-5283.5,100,-5265</points>
<intersection>-5283.5 3</intersection>
<intersection>-5272.5 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-5272.5,103.5,-5272.5</points>
<connection>
<GID>1705</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-5265,100,-5265</points>
<connection>
<GID>1709</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100,-5283.5,120.5,-5283.5</points>
<intersection>100 0</intersection>
<intersection>120.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>120.5,-5283.5,120.5,-5276.5</points>
<connection>
<GID>1710</GID>
<name>IN_0</name></connection>
<intersection>-5283.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>193.5,-5275.5,203,-5275.5</points>
<connection>
<GID>1505</GID>
<name>OUT</name></connection>
<connection>
<GID>1713</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-5284,184.5,-5265</points>
<intersection>-5284 3</intersection>
<intersection>-5274.5 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-5274.5,187.5,-5274.5</points>
<connection>
<GID>1505</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-5265,184.5,-5265</points>
<connection>
<GID>1712</GID>
<name>OUT_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184.5,-5284,205,-5284</points>
<intersection>184.5 0</intersection>
<intersection>205 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>205,-5284,205,-5278.5</points>
<connection>
<GID>1713</GID>
<name>IN_0</name></connection>
<intersection>-5284 3</intersection></vsegment></shape></wire>
<wire>
<ID>1184</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>267.5,-5275.5,276.5,-5275.5</points>
<connection>
<GID>1711</GID>
<name>OUT</name></connection>
<connection>
<GID>1507</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-5285.5,258,-5265</points>
<connection>
<GID>1506</GID>
<name>OUT_0</name></connection>
<intersection>-5285.5 3</intersection>
<intersection>-5274.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-5274.5,261.5,-5274.5</points>
<connection>
<GID>1711</GID>
<name>IN_0</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258,-5285.5,278.5,-5285.5</points>
<intersection>258 0</intersection>
<intersection>278.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>278.5,-5285.5,278.5,-5278.5</points>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection>
<intersection>-5285.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358.5,-5277,368,-5277</points>
<connection>
<GID>1511</GID>
<name>OUT</name></connection>
<connection>
<GID>1510</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-5285.5,349.5,-5265</points>
<intersection>-5285.5 3</intersection>
<intersection>-5276 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349.5,-5276,352.5,-5276</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,-5265,349.5,-5265</points>
<connection>
<GID>1509</GID>
<name>OUT_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>349.5,-5285.5,370,-5285.5</points>
<intersection>349.5 0</intersection>
<intersection>370 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>370,-5285.5,370,-5280</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<intersection>-5285.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1188</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>432.5,-5277,441.5,-5277</points>
<connection>
<GID>1508</GID>
<name>OUT</name></connection>
<connection>
<GID>1513</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423,-5285.5,423,-5265</points>
<intersection>-5285.5 3</intersection>
<intersection>-5276 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,-5276,426.5,-5276</points>
<connection>
<GID>1508</GID>
<name>IN_0</name></connection>
<intersection>423 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422,-5265,423,-5265</points>
<connection>
<GID>1512</GID>
<name>OUT_0</name></connection>
<intersection>423 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>423,-5285.5,443.5,-5285.5</points>
<intersection>423 0</intersection>
<intersection>443.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>443.5,-5285.5,443.5,-5280</points>
<connection>
<GID>1513</GID>
<name>IN_0</name></connection>
<intersection>-5285.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>516.5,-5279,526,-5279</points>
<connection>
<GID>1517</GID>
<name>OUT</name></connection>
<connection>
<GID>1516</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507.5,-5285,507.5,-5265</points>
<intersection>-5285 3</intersection>
<intersection>-5278 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507.5,-5278,510.5,-5278</points>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>507.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>506.5,-5265,507.5,-5265</points>
<connection>
<GID>1515</GID>
<name>OUT_0</name></connection>
<intersection>507.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>507.5,-5285,528,-5285</points>
<intersection>507.5 0</intersection>
<intersection>528 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>528,-5285,528,-5282</points>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>-5285 3</intersection></vsegment></shape></wire>
<wire>
<ID>1192</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>590.5,-5279,599.5,-5279</points>
<connection>
<GID>1514</GID>
<name>OUT</name></connection>
<connection>
<GID>1519</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,-5285,581,-5265</points>
<intersection>-5285 3</intersection>
<intersection>-5278 1</intersection>
<intersection>-5265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581,-5278,584.5,-5278</points>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>581 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>580,-5265,581,-5265</points>
<connection>
<GID>1518</GID>
<name>OUT_0</name></connection>
<intersection>581 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>581,-5285,601.5,-5285</points>
<intersection>581 0</intersection>
<intersection>601.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>601.5,-5285,601.5,-5282</points>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>-5285 3</intersection></vsegment></shape></wire>
<wire>
<ID>1194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-5268,574,-5268</points>
<connection>
<GID>1712</GID>
<name>clock</name></connection>
<connection>
<GID>1709</GID>
<name>clock</name></connection>
<connection>
<GID>1706</GID>
<name>clock</name></connection>
<connection>
<GID>1520</GID>
<name>OUT</name></connection>
<connection>
<GID>1518</GID>
<name>clock</name></connection>
<connection>
<GID>1515</GID>
<name>clock</name></connection>
<connection>
<GID>1512</GID>
<name>clock</name></connection>
<connection>
<GID>1509</GID>
<name>clock</name></connection>
<connection>
<GID>1506</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114.5,-5543,-114.5,-5230</points>
<intersection>-5543 3</intersection>
<intersection>-5525 1</intersection>
<intersection>-5230 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-114.5,-5525,-5,-5525</points>
<connection>
<GID>1546</GID>
<name>IN_0</name></connection>
<intersection>-114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5230,-114.5,-5230</points>
<connection>
<GID>1574</GID>
<name>OUT_0</name></connection>
<intersection>-114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-114.5,-5543,-23.5,-5543</points>
<connection>
<GID>1547</GID>
<name>ENABLE_0</name></connection>
<intersection>-114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1196</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21,-5545,591.5,-5545</points>
<connection>
<GID>1547</GID>
<name>OUT_0</name></connection>
<intersection>36.5 38</intersection>
<intersection>110.5 43</intersection>
<intersection>194.5 42</intersection>
<intersection>268.5 45</intersection>
<intersection>359.5 47</intersection>
<intersection>433.5 49</intersection>
<intersection>517.5 51</intersection>
<intersection>591.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36.5,-5545,36.5,-5532.5</points>
<connection>
<GID>1525</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194.5,-5545,194.5,-5534.5</points>
<connection>
<GID>1531</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110.5,-5545,110.5,-5532.5</points>
<connection>
<GID>1522</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268.5,-5545,268.5,-5534.5</points>
<connection>
<GID>1528</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359.5,-5545,359.5,-5536</points>
<connection>
<GID>1537</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433.5,-5545,433.5,-5536</points>
<connection>
<GID>1534</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517.5,-5545,517.5,-5538</points>
<connection>
<GID>1543</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591.5,-5545,591.5,-5538</points>
<connection>
<GID>1540</GID>
<name>IN_1</name></connection>
<intersection>-5545 33</intersection></vsegment></shape></wire>
<wire>
<ID>1197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-5531.5,52,-5531.5</points>
<connection>
<GID>1525</GID>
<name>OUT</name></connection>
<connection>
<GID>1524</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-5540,33.5,-5523</points>
<intersection>-5540 3</intersection>
<intersection>-5530.5 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-5530.5,36.5,-5530.5</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-5523,33.5,-5523</points>
<connection>
<GID>1523</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-5540,54,-5540</points>
<intersection>33.5 0</intersection>
<intersection>54 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54,-5540,54,-5534.5</points>
<connection>
<GID>1524</GID>
<name>IN_0</name></connection>
<intersection>-5540 3</intersection></vsegment></shape></wire>
<wire>
<ID>1199</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116.5,-5531.5,125.5,-5531.5</points>
<connection>
<GID>1522</GID>
<name>OUT</name></connection>
<connection>
<GID>1527</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-5541.5,107,-5523</points>
<intersection>-5541.5 3</intersection>
<intersection>-5530.5 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-5530.5,110.5,-5530.5</points>
<connection>
<GID>1522</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,-5523,107,-5523</points>
<connection>
<GID>1526</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107,-5541.5,127.5,-5541.5</points>
<intersection>107 0</intersection>
<intersection>127.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127.5,-5541.5,127.5,-5534.5</points>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection>
<intersection>-5541.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,-5533.5,210,-5533.5</points>
<connection>
<GID>1531</GID>
<name>OUT</name></connection>
<connection>
<GID>1530</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-5542,191.5,-5523</points>
<intersection>-5542 3</intersection>
<intersection>-5532.5 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-5532.5,194.5,-5532.5</points>
<connection>
<GID>1531</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190.5,-5523,191.5,-5523</points>
<connection>
<GID>1529</GID>
<name>OUT_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191.5,-5542,212,-5542</points>
<intersection>191.5 0</intersection>
<intersection>212 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>212,-5542,212,-5536.5</points>
<connection>
<GID>1530</GID>
<name>IN_0</name></connection>
<intersection>-5542 3</intersection></vsegment></shape></wire>
<wire>
<ID>1203</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274.5,-5533.5,283.5,-5533.5</points>
<connection>
<GID>1528</GID>
<name>OUT</name></connection>
<connection>
<GID>1533</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265,-5543.5,265,-5523</points>
<connection>
<GID>1532</GID>
<name>OUT_0</name></connection>
<intersection>-5543.5 3</intersection>
<intersection>-5532.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265,-5532.5,268.5,-5532.5</points>
<connection>
<GID>1528</GID>
<name>IN_0</name></connection>
<intersection>265 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>265,-5543.5,285.5,-5543.5</points>
<intersection>265 0</intersection>
<intersection>285.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285.5,-5543.5,285.5,-5536.5</points>
<connection>
<GID>1533</GID>
<name>IN_0</name></connection>
<intersection>-5543.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365.5,-5535,375,-5535</points>
<connection>
<GID>1537</GID>
<name>OUT</name></connection>
<connection>
<GID>1536</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,-5543.5,356.5,-5523</points>
<intersection>-5543.5 3</intersection>
<intersection>-5534 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356.5,-5534,359.5,-5534</points>
<connection>
<GID>1537</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355.5,-5523,356.5,-5523</points>
<connection>
<GID>1535</GID>
<name>OUT_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356.5,-5543.5,377,-5543.5</points>
<intersection>356.5 0</intersection>
<intersection>377 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>377,-5543.5,377,-5538</points>
<connection>
<GID>1536</GID>
<name>IN_0</name></connection>
<intersection>-5543.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1207</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439.5,-5535,448.5,-5535</points>
<connection>
<GID>1534</GID>
<name>OUT</name></connection>
<connection>
<GID>1539</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,-5543.5,430,-5523</points>
<intersection>-5543.5 3</intersection>
<intersection>-5534 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430,-5534,433.5,-5534</points>
<connection>
<GID>1534</GID>
<name>IN_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>429,-5523,430,-5523</points>
<connection>
<GID>1538</GID>
<name>OUT_0</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>430,-5543.5,450.5,-5543.5</points>
<intersection>430 0</intersection>
<intersection>450.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450.5,-5543.5,450.5,-5538</points>
<connection>
<GID>1539</GID>
<name>IN_0</name></connection>
<intersection>-5543.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523.5,-5537,533,-5537</points>
<connection>
<GID>1543</GID>
<name>OUT</name></connection>
<connection>
<GID>1542</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514.5,-5543,514.5,-5523</points>
<intersection>-5543 3</intersection>
<intersection>-5536 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514.5,-5536,517.5,-5536</points>
<connection>
<GID>1543</GID>
<name>IN_0</name></connection>
<intersection>514.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513.5,-5523,514.5,-5523</points>
<connection>
<GID>1541</GID>
<name>OUT_0</name></connection>
<intersection>514.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514.5,-5543,535,-5543</points>
<intersection>514.5 0</intersection>
<intersection>535 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>535,-5543,535,-5540</points>
<connection>
<GID>1542</GID>
<name>IN_0</name></connection>
<intersection>-5543 3</intersection></vsegment></shape></wire>
<wire>
<ID>1211</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597.5,-5537,606.5,-5537</points>
<connection>
<GID>1540</GID>
<name>OUT</name></connection>
<connection>
<GID>1545</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588,-5543,588,-5523</points>
<intersection>-5543 3</intersection>
<intersection>-5536 1</intersection>
<intersection>-5523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588,-5536,591.5,-5536</points>
<connection>
<GID>1540</GID>
<name>IN_0</name></connection>
<intersection>588 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587,-5523,588,-5523</points>
<connection>
<GID>1544</GID>
<name>OUT_0</name></connection>
<intersection>588 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>588,-5543,608.5,-5543</points>
<intersection>588 0</intersection>
<intersection>608.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608.5,-5543,608.5,-5540</points>
<connection>
<GID>1545</GID>
<name>IN_0</name></connection>
<intersection>-5543 3</intersection></vsegment></shape></wire>
<wire>
<ID>1213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-5526,581,-5526</points>
<connection>
<GID>1523</GID>
<name>clock</name></connection>
<connection>
<GID>1526</GID>
<name>clock</name></connection>
<connection>
<GID>1529</GID>
<name>clock</name></connection>
<connection>
<GID>1535</GID>
<name>clock</name></connection>
<connection>
<GID>1538</GID>
<name>clock</name></connection>
<connection>
<GID>1541</GID>
<name>clock</name></connection>
<connection>
<GID>1544</GID>
<name>clock</name></connection>
<connection>
<GID>1546</GID>
<name>OUT</name></connection>
<connection>
<GID>1532</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112.5,-5453,-112.5,-5229</points>
<intersection>-5453 3</intersection>
<intersection>-5435 1</intersection>
<intersection>-5229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112.5,-5435,-8,-5435</points>
<connection>
<GID>1572</GID>
<name>IN_0</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5229,-112.5,-5229</points>
<connection>
<GID>1574</GID>
<name>OUT_1</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112.5,-5453,-26.5,-5453</points>
<connection>
<GID>1573</GID>
<name>ENABLE_0</name></connection>
<intersection>-112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1215</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-24,-5455,588.5,-5455</points>
<connection>
<GID>1573</GID>
<name>OUT_0</name></connection>
<intersection>33.5 38</intersection>
<intersection>107.5 43</intersection>
<intersection>191.5 42</intersection>
<intersection>265.5 45</intersection>
<intersection>356.5 47</intersection>
<intersection>430.5 49</intersection>
<intersection>514.5 51</intersection>
<intersection>588.5 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>33.5,-5455,33.5,-5442.5</points>
<connection>
<GID>1551</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>191.5,-5455,191.5,-5444.5</points>
<connection>
<GID>1557</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>107.5,-5455,107.5,-5442.5</points>
<connection>
<GID>1548</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>265.5,-5455,265.5,-5444.5</points>
<connection>
<GID>1554</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>356.5,-5455,356.5,-5446</points>
<connection>
<GID>1563</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>430.5,-5455,430.5,-5446</points>
<connection>
<GID>1560</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>514.5,-5455,514.5,-5448</points>
<connection>
<GID>1569</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>588.5,-5455,588.5,-5448</points>
<connection>
<GID>1566</GID>
<name>IN_1</name></connection>
<intersection>-5455 33</intersection></vsegment></shape></wire>
<wire>
<ID>1216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-5441.5,49,-5441.5</points>
<connection>
<GID>1551</GID>
<name>OUT</name></connection>
<connection>
<GID>1550</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-5450,30.5,-5433</points>
<intersection>-5450 3</intersection>
<intersection>-5440.5 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-5440.5,33.5,-5440.5</points>
<connection>
<GID>1551</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-5433,30.5,-5433</points>
<connection>
<GID>1549</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-5450,51,-5450</points>
<intersection>30.5 0</intersection>
<intersection>51 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51,-5450,51,-5444.5</points>
<connection>
<GID>1550</GID>
<name>IN_0</name></connection>
<intersection>-5450 3</intersection></vsegment></shape></wire>
<wire>
<ID>1218</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113.5,-5441.5,122.5,-5441.5</points>
<connection>
<GID>1548</GID>
<name>OUT</name></connection>
<connection>
<GID>1553</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-5451.5,104,-5433</points>
<intersection>-5451.5 3</intersection>
<intersection>-5440.5 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-5440.5,107.5,-5440.5</points>
<connection>
<GID>1548</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-5433,104,-5433</points>
<connection>
<GID>1552</GID>
<name>OUT_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-5451.5,124.5,-5451.5</points>
<intersection>104 0</intersection>
<intersection>124.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124.5,-5451.5,124.5,-5444.5</points>
<connection>
<GID>1553</GID>
<name>IN_0</name></connection>
<intersection>-5451.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197.5,-5443.5,207,-5443.5</points>
<connection>
<GID>1557</GID>
<name>OUT</name></connection>
<connection>
<GID>1556</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-5452,188.5,-5433</points>
<intersection>-5452 3</intersection>
<intersection>-5442.5 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-5442.5,191.5,-5442.5</points>
<connection>
<GID>1557</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-5433,188.5,-5433</points>
<connection>
<GID>1555</GID>
<name>OUT_0</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188.5,-5452,209,-5452</points>
<intersection>188.5 0</intersection>
<intersection>209 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209,-5452,209,-5446.5</points>
<connection>
<GID>1556</GID>
<name>IN_0</name></connection>
<intersection>-5452 3</intersection></vsegment></shape></wire>
<wire>
<ID>1222</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>271.5,-5443.5,280.5,-5443.5</points>
<connection>
<GID>1554</GID>
<name>OUT</name></connection>
<connection>
<GID>1559</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-5453.5,262,-5433</points>
<connection>
<GID>1558</GID>
<name>OUT_0</name></connection>
<intersection>-5453.5 3</intersection>
<intersection>-5442.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-5442.5,265.5,-5442.5</points>
<connection>
<GID>1554</GID>
<name>IN_0</name></connection>
<intersection>262 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262,-5453.5,282.5,-5453.5</points>
<intersection>262 0</intersection>
<intersection>282.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282.5,-5453.5,282.5,-5446.5</points>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection>
<intersection>-5453.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362.5,-5445,372,-5445</points>
<connection>
<GID>1563</GID>
<name>OUT</name></connection>
<connection>
<GID>1562</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353.5,-5453.5,353.5,-5433</points>
<intersection>-5453.5 3</intersection>
<intersection>-5444 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353.5,-5444,356.5,-5444</points>
<connection>
<GID>1563</GID>
<name>IN_0</name></connection>
<intersection>353.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352.5,-5433,353.5,-5433</points>
<connection>
<GID>1561</GID>
<name>OUT_0</name></connection>
<intersection>353.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353.5,-5453.5,374,-5453.5</points>
<intersection>353.5 0</intersection>
<intersection>374 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374,-5453.5,374,-5448</points>
<connection>
<GID>1562</GID>
<name>IN_0</name></connection>
<intersection>-5453.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1226</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>436.5,-5445,445.5,-5445</points>
<connection>
<GID>1560</GID>
<name>OUT</name></connection>
<connection>
<GID>1565</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427,-5453.5,427,-5433</points>
<intersection>-5453.5 3</intersection>
<intersection>-5444 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427,-5444,430.5,-5444</points>
<connection>
<GID>1560</GID>
<name>IN_0</name></connection>
<intersection>427 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426,-5433,427,-5433</points>
<connection>
<GID>1564</GID>
<name>OUT_0</name></connection>
<intersection>427 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427,-5453.5,447.5,-5453.5</points>
<intersection>427 0</intersection>
<intersection>447.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447.5,-5453.5,447.5,-5448</points>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection>
<intersection>-5453.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520.5,-5447,530,-5447</points>
<connection>
<GID>1569</GID>
<name>OUT</name></connection>
<connection>
<GID>1568</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-5453,511.5,-5433</points>
<intersection>-5453 3</intersection>
<intersection>-5446 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511.5,-5446,514.5,-5446</points>
<connection>
<GID>1569</GID>
<name>IN_0</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>510.5,-5433,511.5,-5433</points>
<connection>
<GID>1567</GID>
<name>OUT_0</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511.5,-5453,532,-5453</points>
<intersection>511.5 0</intersection>
<intersection>532 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532,-5453,532,-5450</points>
<connection>
<GID>1568</GID>
<name>IN_0</name></connection>
<intersection>-5453 3</intersection></vsegment></shape></wire>
<wire>
<ID>1230</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>594.5,-5447,603.5,-5447</points>
<connection>
<GID>1566</GID>
<name>OUT</name></connection>
<connection>
<GID>1571</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585,-5453,585,-5433</points>
<intersection>-5453 3</intersection>
<intersection>-5446 1</intersection>
<intersection>-5433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585,-5446,588.5,-5446</points>
<connection>
<GID>1566</GID>
<name>IN_0</name></connection>
<intersection>585 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584,-5433,585,-5433</points>
<connection>
<GID>1570</GID>
<name>OUT_0</name></connection>
<intersection>585 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585,-5453,605.5,-5453</points>
<intersection>585 0</intersection>
<intersection>605.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>605.5,-5453,605.5,-5450</points>
<connection>
<GID>1571</GID>
<name>IN_0</name></connection>
<intersection>-5453 3</intersection></vsegment></shape></wire>
<wire>
<ID>1232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-5436,578,-5436</points>
<connection>
<GID>1572</GID>
<name>OUT</name></connection>
<connection>
<GID>1570</GID>
<name>clock</name></connection>
<connection>
<GID>1567</GID>
<name>clock</name></connection>
<connection>
<GID>1564</GID>
<name>clock</name></connection>
<connection>
<GID>1561</GID>
<name>clock</name></connection>
<connection>
<GID>1558</GID>
<name>clock</name></connection>
<connection>
<GID>1555</GID>
<name>clock</name></connection>
<connection>
<GID>1552</GID>
<name>clock</name></connection>
<connection>
<GID>1549</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113,-6095.5,-113,-5852.5</points>
<intersection>-6095.5 2</intersection>
<intersection>-5870.5 3</intersection>
<intersection>-5852.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-113,-5852.5,-11.5,-5852.5</points>
<connection>
<GID>1808</GID>
<name>IN_0</name></connection>
<intersection>-113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6095.5,-113,-6095.5</points>
<connection>
<GID>1783</GID>
<name>OUT_6</name></connection>
<intersection>-113 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-113,-5870.5,-30,-5870.5</points>
<connection>
<GID>1809</GID>
<name>ENABLE_0</name></connection>
<intersection>-113 0</intersection></hsegment></shape></wire>
<wire>
<ID>1234</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-27.5,-5872.5,585,-5872.5</points>
<connection>
<GID>1809</GID>
<name>OUT_0</name></connection>
<intersection>30 38</intersection>
<intersection>104 43</intersection>
<intersection>188 42</intersection>
<intersection>262 45</intersection>
<intersection>353 47</intersection>
<intersection>427 49</intersection>
<intersection>511 51</intersection>
<intersection>585 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>30,-5872.5,30,-5860</points>
<connection>
<GID>1787</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>188,-5872.5,188,-5862</points>
<connection>
<GID>1793</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>104,-5872.5,104,-5860</points>
<connection>
<GID>1784</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>262,-5872.5,262,-5862</points>
<connection>
<GID>1790</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>353,-5872.5,353,-5863.5</points>
<connection>
<GID>1799</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>427,-5872.5,427,-5863.5</points>
<connection>
<GID>1796</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>511,-5872.5,511,-5865.5</points>
<connection>
<GID>1805</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>585,-5872.5,585,-5865.5</points>
<connection>
<GID>1802</GID>
<name>IN_1</name></connection>
<intersection>-5872.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-5859,45.5,-5859</points>
<connection>
<GID>1787</GID>
<name>OUT</name></connection>
<connection>
<GID>1786</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-5867.5,27,-5850.5</points>
<intersection>-5867.5 3</intersection>
<intersection>-5858 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-5858,30,-5858</points>
<connection>
<GID>1787</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-5850.5,27,-5850.5</points>
<connection>
<GID>1785</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-5867.5,47.5,-5867.5</points>
<intersection>27 0</intersection>
<intersection>47.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-5867.5,47.5,-5862</points>
<connection>
<GID>1786</GID>
<name>IN_0</name></connection>
<intersection>-5867.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1237</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>110,-5859,119,-5859</points>
<connection>
<GID>1784</GID>
<name>OUT</name></connection>
<connection>
<GID>1789</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-5869,100.5,-5850.5</points>
<intersection>-5869 3</intersection>
<intersection>-5858 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-5858,104,-5858</points>
<connection>
<GID>1784</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-5850.5,100.5,-5850.5</points>
<connection>
<GID>1788</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100.5,-5869,121,-5869</points>
<intersection>100.5 0</intersection>
<intersection>121 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>121,-5869,121,-5862</points>
<connection>
<GID>1789</GID>
<name>IN_0</name></connection>
<intersection>-5869 3</intersection></vsegment></shape></wire>
<wire>
<ID>1239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,-5861,203.5,-5861</points>
<connection>
<GID>1793</GID>
<name>OUT</name></connection>
<connection>
<GID>1792</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-5869.5,185,-5850.5</points>
<intersection>-5869.5 3</intersection>
<intersection>-5860 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-5860,188,-5860</points>
<connection>
<GID>1793</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-5850.5,185,-5850.5</points>
<connection>
<GID>1791</GID>
<name>OUT_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185,-5869.5,205.5,-5869.5</points>
<intersection>185 0</intersection>
<intersection>205.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>205.5,-5869.5,205.5,-5864</points>
<connection>
<GID>1792</GID>
<name>IN_0</name></connection>
<intersection>-5869.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1241</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>268,-5861,277,-5861</points>
<connection>
<GID>1790</GID>
<name>OUT</name></connection>
<connection>
<GID>1795</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-5871,258.5,-5850.5</points>
<connection>
<GID>1794</GID>
<name>OUT_0</name></connection>
<intersection>-5871 3</intersection>
<intersection>-5860 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,-5860,262,-5860</points>
<connection>
<GID>1790</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,-5871,279,-5871</points>
<intersection>258.5 0</intersection>
<intersection>279 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>279,-5871,279,-5864</points>
<connection>
<GID>1795</GID>
<name>IN_0</name></connection>
<intersection>-5871 3</intersection></vsegment></shape></wire>
<wire>
<ID>1243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-5862.5,368.5,-5862.5</points>
<connection>
<GID>1799</GID>
<name>OUT</name></connection>
<connection>
<GID>1798</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-5871,350,-5850.5</points>
<intersection>-5871 3</intersection>
<intersection>-5861.5 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-5861.5,353,-5861.5</points>
<connection>
<GID>1799</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-5850.5,350,-5850.5</points>
<connection>
<GID>1797</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>350,-5871,370.5,-5871</points>
<intersection>350 0</intersection>
<intersection>370.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>370.5,-5871,370.5,-5865.5</points>
<connection>
<GID>1798</GID>
<name>IN_0</name></connection>
<intersection>-5871 3</intersection></vsegment></shape></wire>
<wire>
<ID>1245</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>433,-5862.5,442,-5862.5</points>
<connection>
<GID>1796</GID>
<name>OUT</name></connection>
<connection>
<GID>1801</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-5871,423.5,-5850.5</points>
<intersection>-5871 3</intersection>
<intersection>-5861.5 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423.5,-5861.5,427,-5861.5</points>
<connection>
<GID>1796</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422.5,-5850.5,423.5,-5850.5</points>
<connection>
<GID>1800</GID>
<name>OUT_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>423.5,-5871,444,-5871</points>
<intersection>423.5 0</intersection>
<intersection>444 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>444,-5871,444,-5865.5</points>
<connection>
<GID>1801</GID>
<name>IN_0</name></connection>
<intersection>-5871 3</intersection></vsegment></shape></wire>
<wire>
<ID>1247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>517,-5864.5,526.5,-5864.5</points>
<connection>
<GID>1805</GID>
<name>OUT</name></connection>
<connection>
<GID>1804</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508,-5870.5,508,-5850.5</points>
<intersection>-5870.5 3</intersection>
<intersection>-5863.5 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,-5863.5,511,-5863.5</points>
<connection>
<GID>1805</GID>
<name>IN_0</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507,-5850.5,508,-5850.5</points>
<connection>
<GID>1803</GID>
<name>OUT_0</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>508,-5870.5,528.5,-5870.5</points>
<intersection>508 0</intersection>
<intersection>528.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>528.5,-5870.5,528.5,-5867.5</points>
<connection>
<GID>1804</GID>
<name>IN_0</name></connection>
<intersection>-5870.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1249</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>591,-5864.5,600,-5864.5</points>
<connection>
<GID>1802</GID>
<name>OUT</name></connection>
<connection>
<GID>1807</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581.5,-5870.5,581.5,-5850.5</points>
<intersection>-5870.5 3</intersection>
<intersection>-5863.5 1</intersection>
<intersection>-5850.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581.5,-5863.5,585,-5863.5</points>
<connection>
<GID>1802</GID>
<name>IN_0</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>580.5,-5850.5,581.5,-5850.5</points>
<connection>
<GID>1806</GID>
<name>OUT_0</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>581.5,-5870.5,602,-5870.5</points>
<intersection>581.5 0</intersection>
<intersection>602 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>602,-5870.5,602,-5867.5</points>
<connection>
<GID>1807</GID>
<name>IN_0</name></connection>
<intersection>-5870.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-5853.5,574.5,-5853.5</points>
<connection>
<GID>1808</GID>
<name>OUT</name></connection>
<connection>
<GID>1806</GID>
<name>clock</name></connection>
<connection>
<GID>1803</GID>
<name>clock</name></connection>
<connection>
<GID>1800</GID>
<name>clock</name></connection>
<connection>
<GID>1797</GID>
<name>clock</name></connection>
<connection>
<GID>1794</GID>
<name>clock</name></connection>
<connection>
<GID>1791</GID>
<name>clock</name></connection>
<connection>
<GID>1788</GID>
<name>clock</name></connection>
<connection>
<GID>1785</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114,-6094.5,-114,-5762.5</points>
<intersection>-6094.5 2</intersection>
<intersection>-5780.5 3</intersection>
<intersection>-5762.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-114,-5762.5,-14.5,-5762.5</points>
<connection>
<GID>1834</GID>
<name>IN_0</name></connection>
<intersection>-114 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6094.5,-114,-6094.5</points>
<connection>
<GID>1783</GID>
<name>OUT_7</name></connection>
<intersection>-114 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-114,-5780.5,-33,-5780.5</points>
<connection>
<GID>1835</GID>
<name>ENABLE_0</name></connection>
<intersection>-114 0</intersection></hsegment></shape></wire>
<wire>
<ID>1253</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-30.5,-5782.5,582,-5782.5</points>
<connection>
<GID>1835</GID>
<name>OUT_0</name></connection>
<intersection>27 38</intersection>
<intersection>101 43</intersection>
<intersection>185 42</intersection>
<intersection>259 45</intersection>
<intersection>350 47</intersection>
<intersection>424 49</intersection>
<intersection>508 51</intersection>
<intersection>582 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>27,-5782.5,27,-5770</points>
<connection>
<GID>1813</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>185,-5782.5,185,-5772</points>
<connection>
<GID>1819</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>101,-5782.5,101,-5770</points>
<connection>
<GID>1810</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>259,-5782.5,259,-5772</points>
<connection>
<GID>1816</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>350,-5782.5,350,-5773.5</points>
<connection>
<GID>1825</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>424,-5782.5,424,-5773.5</points>
<connection>
<GID>1822</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>508,-5782.5,508,-5775.5</points>
<connection>
<GID>1831</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>582,-5782.5,582,-5775.5</points>
<connection>
<GID>1828</GID>
<name>IN_1</name></connection>
<intersection>-5782.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-5769,42.5,-5769</points>
<connection>
<GID>1813</GID>
<name>OUT</name></connection>
<connection>
<GID>1812</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-5777.5,24,-5760.5</points>
<intersection>-5777.5 3</intersection>
<intersection>-5768 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-5768,27,-5768</points>
<connection>
<GID>1813</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-5760.5,24,-5760.5</points>
<connection>
<GID>1811</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-5777.5,44.5,-5777.5</points>
<intersection>24 0</intersection>
<intersection>44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-5777.5,44.5,-5772</points>
<connection>
<GID>1812</GID>
<name>IN_0</name></connection>
<intersection>-5777.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1256</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>107,-5769,116,-5769</points>
<connection>
<GID>1810</GID>
<name>OUT</name></connection>
<connection>
<GID>1815</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-5779,97.5,-5760.5</points>
<intersection>-5779 3</intersection>
<intersection>-5768 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-5768,101,-5768</points>
<connection>
<GID>1810</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-5760.5,97.5,-5760.5</points>
<connection>
<GID>1814</GID>
<name>OUT_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>97.5,-5779,118,-5779</points>
<intersection>97.5 0</intersection>
<intersection>118 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>118,-5779,118,-5772</points>
<connection>
<GID>1815</GID>
<name>IN_0</name></connection>
<intersection>-5779 3</intersection></vsegment></shape></wire>
<wire>
<ID>1258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191,-5771,200.5,-5771</points>
<connection>
<GID>1819</GID>
<name>OUT</name></connection>
<connection>
<GID>1818</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-5779.5,182,-5760.5</points>
<intersection>-5779.5 3</intersection>
<intersection>-5770 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>182,-5770,185,-5770</points>
<connection>
<GID>1819</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181,-5760.5,182,-5760.5</points>
<connection>
<GID>1817</GID>
<name>OUT_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>182,-5779.5,202.5,-5779.5</points>
<intersection>182 0</intersection>
<intersection>202.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>202.5,-5779.5,202.5,-5774</points>
<connection>
<GID>1818</GID>
<name>IN_0</name></connection>
<intersection>-5779.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1260</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>265,-5771,274,-5771</points>
<connection>
<GID>1816</GID>
<name>OUT</name></connection>
<connection>
<GID>1821</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-5781,255.5,-5760.5</points>
<connection>
<GID>1820</GID>
<name>OUT_0</name></connection>
<intersection>-5781 3</intersection>
<intersection>-5770 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-5770,259,-5770</points>
<connection>
<GID>1816</GID>
<name>IN_0</name></connection>
<intersection>255.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>255.5,-5781,276,-5781</points>
<intersection>255.5 0</intersection>
<intersection>276 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>276,-5781,276,-5774</points>
<connection>
<GID>1821</GID>
<name>IN_0</name></connection>
<intersection>-5781 3</intersection></vsegment></shape></wire>
<wire>
<ID>1262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>356,-5772.5,365.5,-5772.5</points>
<connection>
<GID>1825</GID>
<name>OUT</name></connection>
<connection>
<GID>1824</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,-5781,347,-5760.5</points>
<intersection>-5781 3</intersection>
<intersection>-5771.5 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,-5771.5,350,-5771.5</points>
<connection>
<GID>1825</GID>
<name>IN_0</name></connection>
<intersection>347 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346,-5760.5,347,-5760.5</points>
<connection>
<GID>1823</GID>
<name>OUT_0</name></connection>
<intersection>347 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>347,-5781,367.5,-5781</points>
<intersection>347 0</intersection>
<intersection>367.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>367.5,-5781,367.5,-5775.5</points>
<connection>
<GID>1824</GID>
<name>IN_0</name></connection>
<intersection>-5781 3</intersection></vsegment></shape></wire>
<wire>
<ID>1264</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>430,-5772.5,439,-5772.5</points>
<connection>
<GID>1822</GID>
<name>OUT</name></connection>
<connection>
<GID>1827</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420.5,-5781,420.5,-5760.5</points>
<intersection>-5781 3</intersection>
<intersection>-5771.5 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420.5,-5771.5,424,-5771.5</points>
<connection>
<GID>1822</GID>
<name>IN_0</name></connection>
<intersection>420.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>419.5,-5760.5,420.5,-5760.5</points>
<connection>
<GID>1826</GID>
<name>OUT_0</name></connection>
<intersection>420.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>420.5,-5781,441,-5781</points>
<intersection>420.5 0</intersection>
<intersection>441 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>441,-5781,441,-5775.5</points>
<connection>
<GID>1827</GID>
<name>IN_0</name></connection>
<intersection>-5781 3</intersection></vsegment></shape></wire>
<wire>
<ID>1266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>514,-5774.5,523.5,-5774.5</points>
<connection>
<GID>1831</GID>
<name>OUT</name></connection>
<connection>
<GID>1830</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505,-5780.5,505,-5760.5</points>
<intersection>-5780.5 3</intersection>
<intersection>-5773.5 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505,-5773.5,508,-5773.5</points>
<connection>
<GID>1831</GID>
<name>IN_0</name></connection>
<intersection>505 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>504,-5760.5,505,-5760.5</points>
<connection>
<GID>1829</GID>
<name>OUT_0</name></connection>
<intersection>505 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>505,-5780.5,525.5,-5780.5</points>
<intersection>505 0</intersection>
<intersection>525.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>525.5,-5780.5,525.5,-5777.5</points>
<connection>
<GID>1830</GID>
<name>IN_0</name></connection>
<intersection>-5780.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1268</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>588,-5774.5,597,-5774.5</points>
<connection>
<GID>1828</GID>
<name>OUT</name></connection>
<connection>
<GID>1833</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>578.5,-5780.5,578.5,-5760.5</points>
<intersection>-5780.5 3</intersection>
<intersection>-5773.5 1</intersection>
<intersection>-5760.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>578.5,-5773.5,582,-5773.5</points>
<connection>
<GID>1828</GID>
<name>IN_0</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>577.5,-5760.5,578.5,-5760.5</points>
<connection>
<GID>1832</GID>
<name>OUT_0</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>578.5,-5780.5,599,-5780.5</points>
<intersection>578.5 0</intersection>
<intersection>599 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>599,-5780.5,599,-5777.5</points>
<connection>
<GID>1833</GID>
<name>IN_0</name></connection>
<intersection>-5780.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-5763.5,571.5,-5763.5</points>
<connection>
<GID>1811</GID>
<name>clock</name></connection>
<connection>
<GID>1814</GID>
<name>clock</name></connection>
<connection>
<GID>1817</GID>
<name>clock</name></connection>
<connection>
<GID>1820</GID>
<name>clock</name></connection>
<connection>
<GID>1823</GID>
<name>clock</name></connection>
<connection>
<GID>1826</GID>
<name>clock</name></connection>
<connection>
<GID>1829</GID>
<name>clock</name></connection>
<connection>
<GID>1834</GID>
<name>OUT</name></connection>
<connection>
<GID>1832</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-6097.5,-111,-6020.5</points>
<intersection>-6097.5 2</intersection>
<intersection>-6038.5 3</intersection>
<intersection>-6020.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-6020.5,-7.5,-6020.5</points>
<connection>
<GID>1860</GID>
<name>IN_0</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6097.5,-111,-6097.5</points>
<connection>
<GID>1783</GID>
<name>OUT_4</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111,-6038.5,-26,-6038.5</points>
<connection>
<GID>1861</GID>
<name>ENABLE_0</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>1272</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-23.5,-6040.5,589,-6040.5</points>
<connection>
<GID>1861</GID>
<name>OUT_0</name></connection>
<intersection>34 38</intersection>
<intersection>108 43</intersection>
<intersection>192 42</intersection>
<intersection>266 45</intersection>
<intersection>357 47</intersection>
<intersection>431 49</intersection>
<intersection>515 51</intersection>
<intersection>589 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>34,-6040.5,34,-6028</points>
<connection>
<GID>1839</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>192,-6040.5,192,-6030</points>
<connection>
<GID>1845</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>108,-6040.5,108,-6028</points>
<connection>
<GID>1836</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>266,-6040.5,266,-6030</points>
<connection>
<GID>1842</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>357,-6040.5,357,-6031.5</points>
<connection>
<GID>1851</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>431,-6040.5,431,-6031.5</points>
<connection>
<GID>1848</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>515,-6040.5,515,-6033.5</points>
<connection>
<GID>1857</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>589,-6040.5,589,-6033.5</points>
<connection>
<GID>1854</GID>
<name>IN_1</name></connection>
<intersection>-6040.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-6027,49.5,-6027</points>
<connection>
<GID>1839</GID>
<name>OUT</name></connection>
<connection>
<GID>1838</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-6035.5,31,-6018.5</points>
<intersection>-6035.5 3</intersection>
<intersection>-6026 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-6026,34,-6026</points>
<connection>
<GID>1839</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-6018.5,31,-6018.5</points>
<connection>
<GID>1837</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-6035.5,51.5,-6035.5</points>
<intersection>31 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-6035.5,51.5,-6030</points>
<connection>
<GID>1838</GID>
<name>IN_0</name></connection>
<intersection>-6035.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1275</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114,-6027,123,-6027</points>
<connection>
<GID>1836</GID>
<name>OUT</name></connection>
<connection>
<GID>1841</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-6037,104.5,-6018.5</points>
<intersection>-6037 3</intersection>
<intersection>-6026 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-6026,108,-6026</points>
<connection>
<GID>1836</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-6018.5,104.5,-6018.5</points>
<connection>
<GID>1840</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-6037,125,-6037</points>
<intersection>104.5 0</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-6037,125,-6030</points>
<connection>
<GID>1841</GID>
<name>IN_0</name></connection>
<intersection>-6037 3</intersection></vsegment></shape></wire>
<wire>
<ID>1277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-6029,207.5,-6029</points>
<connection>
<GID>1845</GID>
<name>OUT</name></connection>
<connection>
<GID>1844</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-6037.5,189,-6018.5</points>
<intersection>-6037.5 3</intersection>
<intersection>-6028 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-6028,192,-6028</points>
<connection>
<GID>1845</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188,-6018.5,189,-6018.5</points>
<connection>
<GID>1843</GID>
<name>OUT_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189,-6037.5,209.5,-6037.5</points>
<intersection>189 0</intersection>
<intersection>209.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>209.5,-6037.5,209.5,-6032</points>
<connection>
<GID>1844</GID>
<name>IN_0</name></connection>
<intersection>-6037.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1279</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>272,-6029,281,-6029</points>
<connection>
<GID>1842</GID>
<name>OUT</name></connection>
<connection>
<GID>1847</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-6039,262.5,-6018.5</points>
<connection>
<GID>1846</GID>
<name>OUT_0</name></connection>
<intersection>-6039 3</intersection>
<intersection>-6028 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-6028,266,-6028</points>
<connection>
<GID>1842</GID>
<name>IN_0</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>262.5,-6039,283,-6039</points>
<intersection>262.5 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-6039,283,-6032</points>
<connection>
<GID>1847</GID>
<name>IN_0</name></connection>
<intersection>-6039 3</intersection></vsegment></shape></wire>
<wire>
<ID>1281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363,-6030.5,372.5,-6030.5</points>
<connection>
<GID>1851</GID>
<name>OUT</name></connection>
<connection>
<GID>1850</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-6039,354,-6018.5</points>
<intersection>-6039 3</intersection>
<intersection>-6029.5 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-6029.5,357,-6029.5</points>
<connection>
<GID>1851</GID>
<name>IN_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-6018.5,354,-6018.5</points>
<connection>
<GID>1849</GID>
<name>OUT_0</name></connection>
<intersection>354 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>354,-6039,374.5,-6039</points>
<intersection>354 0</intersection>
<intersection>374.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>374.5,-6039,374.5,-6033.5</points>
<connection>
<GID>1850</GID>
<name>IN_0</name></connection>
<intersection>-6039 3</intersection></vsegment></shape></wire>
<wire>
<ID>1283</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>437,-6030.5,446,-6030.5</points>
<connection>
<GID>1848</GID>
<name>OUT</name></connection>
<connection>
<GID>1853</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-6039,427.5,-6018.5</points>
<intersection>-6039 3</intersection>
<intersection>-6029.5 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-6029.5,431,-6029.5</points>
<connection>
<GID>1848</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426.5,-6018.5,427.5,-6018.5</points>
<connection>
<GID>1852</GID>
<name>OUT_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-6039,448,-6039</points>
<intersection>427.5 0</intersection>
<intersection>448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>448,-6039,448,-6033.5</points>
<connection>
<GID>1853</GID>
<name>IN_0</name></connection>
<intersection>-6039 3</intersection></vsegment></shape></wire>
<wire>
<ID>1285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>521,-6032.5,530.5,-6032.5</points>
<connection>
<GID>1857</GID>
<name>OUT</name></connection>
<connection>
<GID>1856</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512,-6038.5,512,-6018.5</points>
<intersection>-6038.5 3</intersection>
<intersection>-6031.5 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-6031.5,515,-6031.5</points>
<connection>
<GID>1857</GID>
<name>IN_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,-6018.5,512,-6018.5</points>
<connection>
<GID>1855</GID>
<name>OUT_0</name></connection>
<intersection>512 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>512,-6038.5,532.5,-6038.5</points>
<intersection>512 0</intersection>
<intersection>532.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>532.5,-6038.5,532.5,-6035.5</points>
<connection>
<GID>1856</GID>
<name>IN_0</name></connection>
<intersection>-6038.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1287</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>595,-6032.5,604,-6032.5</points>
<connection>
<GID>1854</GID>
<name>OUT</name></connection>
<connection>
<GID>1859</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-6038.5,585.5,-6018.5</points>
<intersection>-6038.5 3</intersection>
<intersection>-6031.5 1</intersection>
<intersection>-6018.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-6031.5,589,-6031.5</points>
<connection>
<GID>1854</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>584.5,-6018.5,585.5,-6018.5</points>
<connection>
<GID>1858</GID>
<name>OUT_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-6038.5,606,-6038.5</points>
<intersection>585.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-6038.5,606,-6035.5</points>
<connection>
<GID>1859</GID>
<name>IN_0</name></connection>
<intersection>-6038.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-6021.5,578.5,-6021.5</points>
<connection>
<GID>1837</GID>
<name>clock</name></connection>
<connection>
<GID>1840</GID>
<name>clock</name></connection>
<connection>
<GID>1843</GID>
<name>clock</name></connection>
<connection>
<GID>1846</GID>
<name>clock</name></connection>
<connection>
<GID>1849</GID>
<name>clock</name></connection>
<connection>
<GID>1852</GID>
<name>clock</name></connection>
<connection>
<GID>1858</GID>
<name>clock</name></connection>
<connection>
<GID>1860</GID>
<name>OUT</name></connection>
<connection>
<GID>1855</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-6096.5,-112,-5930.5</points>
<intersection>-6096.5 2</intersection>
<intersection>-5948.5 3</intersection>
<intersection>-5930.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112,-5930.5,-10.5,-5930.5</points>
<connection>
<GID>1886</GID>
<name>IN_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6096.5,-112,-6096.5</points>
<connection>
<GID>1783</GID>
<name>OUT_5</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112,-5948.5,-29,-5948.5</points>
<connection>
<GID>1887</GID>
<name>ENABLE_0</name></connection>
<intersection>-112 0</intersection></hsegment></shape></wire>
<wire>
<ID>1291</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-26.5,-5950.5,586,-5950.5</points>
<connection>
<GID>1887</GID>
<name>OUT_0</name></connection>
<intersection>31 38</intersection>
<intersection>105 43</intersection>
<intersection>189 42</intersection>
<intersection>263 45</intersection>
<intersection>354 47</intersection>
<intersection>428 49</intersection>
<intersection>512 51</intersection>
<intersection>586 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>31,-5950.5,31,-5938</points>
<connection>
<GID>1865</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>189,-5950.5,189,-5940</points>
<connection>
<GID>1871</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>105,-5950.5,105,-5938</points>
<connection>
<GID>1862</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>263,-5950.5,263,-5940</points>
<connection>
<GID>1868</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>354,-5950.5,354,-5941.5</points>
<connection>
<GID>1877</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>428,-5950.5,428,-5941.5</points>
<connection>
<GID>1874</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>512,-5950.5,512,-5943.5</points>
<connection>
<GID>1883</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>586,-5950.5,586,-5943.5</points>
<connection>
<GID>1880</GID>
<name>IN_1</name></connection>
<intersection>-5950.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-5937,46.5,-5937</points>
<connection>
<GID>1865</GID>
<name>OUT</name></connection>
<connection>
<GID>1864</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-5945.5,28,-5928.5</points>
<intersection>-5945.5 3</intersection>
<intersection>-5936 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-5936,31,-5936</points>
<connection>
<GID>1865</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-5928.5,28,-5928.5</points>
<connection>
<GID>1863</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-5945.5,48.5,-5945.5</points>
<intersection>28 0</intersection>
<intersection>48.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-5945.5,48.5,-5940</points>
<connection>
<GID>1864</GID>
<name>IN_0</name></connection>
<intersection>-5945.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1294</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>111,-5937,120,-5937</points>
<connection>
<GID>1862</GID>
<name>OUT</name></connection>
<connection>
<GID>1867</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-5947,101.5,-5928.5</points>
<intersection>-5947 3</intersection>
<intersection>-5936 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-5936,105,-5936</points>
<connection>
<GID>1862</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-5928.5,101.5,-5928.5</points>
<connection>
<GID>1866</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101.5,-5947,122,-5947</points>
<intersection>101.5 0</intersection>
<intersection>122 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122,-5947,122,-5940</points>
<connection>
<GID>1867</GID>
<name>IN_0</name></connection>
<intersection>-5947 3</intersection></vsegment></shape></wire>
<wire>
<ID>1296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-5939,204.5,-5939</points>
<connection>
<GID>1871</GID>
<name>OUT</name></connection>
<connection>
<GID>1870</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-5947.5,186,-5928.5</points>
<intersection>-5947.5 3</intersection>
<intersection>-5938 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186,-5938,189,-5938</points>
<connection>
<GID>1871</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-5928.5,186,-5928.5</points>
<connection>
<GID>1869</GID>
<name>OUT_0</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>186,-5947.5,206.5,-5947.5</points>
<intersection>186 0</intersection>
<intersection>206.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>206.5,-5947.5,206.5,-5942</points>
<connection>
<GID>1870</GID>
<name>IN_0</name></connection>
<intersection>-5947.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1298</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>269,-5939,278,-5939</points>
<connection>
<GID>1868</GID>
<name>OUT</name></connection>
<connection>
<GID>1873</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259.5,-5949,259.5,-5928.5</points>
<connection>
<GID>1872</GID>
<name>OUT_0</name></connection>
<intersection>-5949 3</intersection>
<intersection>-5938 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-5938,263,-5938</points>
<connection>
<GID>1868</GID>
<name>IN_0</name></connection>
<intersection>259.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>259.5,-5949,280,-5949</points>
<intersection>259.5 0</intersection>
<intersection>280 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>280,-5949,280,-5942</points>
<connection>
<GID>1873</GID>
<name>IN_0</name></connection>
<intersection>-5949 3</intersection></vsegment></shape></wire>
<wire>
<ID>1300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360,-5940.5,369.5,-5940.5</points>
<connection>
<GID>1877</GID>
<name>OUT</name></connection>
<connection>
<GID>1876</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,-5949,351,-5928.5</points>
<intersection>-5949 3</intersection>
<intersection>-5939.5 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,-5939.5,354,-5939.5</points>
<connection>
<GID>1877</GID>
<name>IN_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-5928.5,351,-5928.5</points>
<connection>
<GID>1875</GID>
<name>OUT_0</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>351,-5949,371.5,-5949</points>
<intersection>351 0</intersection>
<intersection>371.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>371.5,-5949,371.5,-5943.5</points>
<connection>
<GID>1876</GID>
<name>IN_0</name></connection>
<intersection>-5949 3</intersection></vsegment></shape></wire>
<wire>
<ID>1302</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>434,-5940.5,443,-5940.5</points>
<connection>
<GID>1874</GID>
<name>OUT</name></connection>
<connection>
<GID>1879</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,-5949,424.5,-5928.5</points>
<intersection>-5949 3</intersection>
<intersection>-5939.5 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424.5,-5939.5,428,-5939.5</points>
<connection>
<GID>1874</GID>
<name>IN_0</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423.5,-5928.5,424.5,-5928.5</points>
<connection>
<GID>1878</GID>
<name>OUT_0</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>424.5,-5949,445,-5949</points>
<intersection>424.5 0</intersection>
<intersection>445 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>445,-5949,445,-5943.5</points>
<connection>
<GID>1879</GID>
<name>IN_0</name></connection>
<intersection>-5949 3</intersection></vsegment></shape></wire>
<wire>
<ID>1304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>518,-5942.5,527.5,-5942.5</points>
<connection>
<GID>1883</GID>
<name>OUT</name></connection>
<connection>
<GID>1882</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,-5948.5,509,-5928.5</points>
<intersection>-5948.5 3</intersection>
<intersection>-5941.5 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509,-5941.5,512,-5941.5</points>
<connection>
<GID>1883</GID>
<name>IN_0</name></connection>
<intersection>509 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>508,-5928.5,509,-5928.5</points>
<connection>
<GID>1881</GID>
<name>OUT_0</name></connection>
<intersection>509 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>509,-5948.5,529.5,-5948.5</points>
<intersection>509 0</intersection>
<intersection>529.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>529.5,-5948.5,529.5,-5945.5</points>
<connection>
<GID>1882</GID>
<name>IN_0</name></connection>
<intersection>-5948.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1306</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>592,-5942.5,601,-5942.5</points>
<connection>
<GID>1880</GID>
<name>OUT</name></connection>
<connection>
<GID>1885</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>582.5,-5948.5,582.5,-5928.5</points>
<intersection>-5948.5 3</intersection>
<intersection>-5941.5 1</intersection>
<intersection>-5928.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>582.5,-5941.5,586,-5941.5</points>
<connection>
<GID>1880</GID>
<name>IN_0</name></connection>
<intersection>582.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>581.5,-5928.5,582.5,-5928.5</points>
<connection>
<GID>1884</GID>
<name>OUT_0</name></connection>
<intersection>582.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>582.5,-5948.5,603,-5948.5</points>
<intersection>582.5 0</intersection>
<intersection>603 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>603,-5948.5,603,-5945.5</points>
<connection>
<GID>1885</GID>
<name>IN_0</name></connection>
<intersection>-5948.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,-5931.5,575.5,-5931.5</points>
<connection>
<GID>1886</GID>
<name>OUT</name></connection>
<connection>
<GID>1884</GID>
<name>clock</name></connection>
<connection>
<GID>1881</GID>
<name>clock</name></connection>
<connection>
<GID>1878</GID>
<name>clock</name></connection>
<connection>
<GID>1875</GID>
<name>clock</name></connection>
<connection>
<GID>1872</GID>
<name>clock</name></connection>
<connection>
<GID>1869</GID>
<name>clock</name></connection>
<connection>
<GID>1866</GID>
<name>clock</name></connection>
<connection>
<GID>1863</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-6246.5,-112,-6099.5</points>
<intersection>-6246.5 3</intersection>
<intersection>-6228.5 1</intersection>
<intersection>-6099.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112,-6228.5,-9.5,-6228.5</points>
<connection>
<GID>1912</GID>
<name>IN_0</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6099.5,-112,-6099.5</points>
<connection>
<GID>1783</GID>
<name>OUT_2</name></connection>
<intersection>-112 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-112,-6246.5,-28,-6246.5</points>
<connection>
<GID>1913</GID>
<name>ENABLE_0</name></connection>
<intersection>-112 0</intersection></hsegment></shape></wire>
<wire>
<ID>1310</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-25.5,-6248.5,587,-6248.5</points>
<connection>
<GID>1913</GID>
<name>OUT_0</name></connection>
<intersection>32 38</intersection>
<intersection>106 43</intersection>
<intersection>190 42</intersection>
<intersection>264 45</intersection>
<intersection>355 47</intersection>
<intersection>429 49</intersection>
<intersection>513 51</intersection>
<intersection>587 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>32,-6248.5,32,-6236</points>
<connection>
<GID>1891</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>190,-6248.5,190,-6238</points>
<connection>
<GID>1897</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>106,-6248.5,106,-6236</points>
<connection>
<GID>1888</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>264,-6248.5,264,-6238</points>
<connection>
<GID>1894</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>355,-6248.5,355,-6239.5</points>
<connection>
<GID>1903</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>429,-6248.5,429,-6239.5</points>
<connection>
<GID>1900</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>513,-6248.5,513,-6241.5</points>
<connection>
<GID>1909</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>587,-6248.5,587,-6241.5</points>
<connection>
<GID>1906</GID>
<name>IN_1</name></connection>
<intersection>-6248.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-6235,47.5,-6235</points>
<connection>
<GID>1891</GID>
<name>OUT</name></connection>
<connection>
<GID>1890</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-6243.5,29,-6226.5</points>
<intersection>-6243.5 3</intersection>
<intersection>-6234 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-6234,32,-6234</points>
<connection>
<GID>1891</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-6226.5,29,-6226.5</points>
<connection>
<GID>1889</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-6243.5,49.5,-6243.5</points>
<intersection>29 0</intersection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-6243.5,49.5,-6238</points>
<connection>
<GID>1890</GID>
<name>IN_0</name></connection>
<intersection>-6243.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1313</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112,-6235,121,-6235</points>
<connection>
<GID>1888</GID>
<name>OUT</name></connection>
<connection>
<GID>1893</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-6245,102.5,-6226.5</points>
<intersection>-6245 3</intersection>
<intersection>-6234 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-6234,106,-6234</points>
<connection>
<GID>1888</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-6226.5,102.5,-6226.5</points>
<connection>
<GID>1892</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-6245,123,-6245</points>
<intersection>102.5 0</intersection>
<intersection>123 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>123,-6245,123,-6238</points>
<connection>
<GID>1893</GID>
<name>IN_0</name></connection>
<intersection>-6245 3</intersection></vsegment></shape></wire>
<wire>
<ID>1315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,-6237,205.5,-6237</points>
<connection>
<GID>1897</GID>
<name>OUT</name></connection>
<connection>
<GID>1896</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-6245.5,187,-6226.5</points>
<intersection>-6245.5 3</intersection>
<intersection>-6236 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-6236,190,-6236</points>
<connection>
<GID>1897</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-6226.5,187,-6226.5</points>
<connection>
<GID>1895</GID>
<name>OUT_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,-6245.5,207.5,-6245.5</points>
<intersection>187 0</intersection>
<intersection>207.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207.5,-6245.5,207.5,-6240</points>
<connection>
<GID>1896</GID>
<name>IN_0</name></connection>
<intersection>-6245.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1317</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>270,-6237,279,-6237</points>
<connection>
<GID>1894</GID>
<name>OUT</name></connection>
<connection>
<GID>1899</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-6247,260.5,-6226.5</points>
<connection>
<GID>1898</GID>
<name>OUT_0</name></connection>
<intersection>-6247 3</intersection>
<intersection>-6236 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-6236,264,-6236</points>
<connection>
<GID>1894</GID>
<name>IN_0</name></connection>
<intersection>260.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>260.5,-6247,281,-6247</points>
<intersection>260.5 0</intersection>
<intersection>281 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>281,-6247,281,-6240</points>
<connection>
<GID>1899</GID>
<name>IN_0</name></connection>
<intersection>-6247 3</intersection></vsegment></shape></wire>
<wire>
<ID>1319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-6238.5,370.5,-6238.5</points>
<connection>
<GID>1903</GID>
<name>OUT</name></connection>
<connection>
<GID>1902</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-6247,352,-6226.5</points>
<intersection>-6247 3</intersection>
<intersection>-6237.5 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-6237.5,355,-6237.5</points>
<connection>
<GID>1903</GID>
<name>IN_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-6226.5,352,-6226.5</points>
<connection>
<GID>1901</GID>
<name>OUT_0</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>352,-6247,372.5,-6247</points>
<intersection>352 0</intersection>
<intersection>372.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>372.5,-6247,372.5,-6241.5</points>
<connection>
<GID>1902</GID>
<name>IN_0</name></connection>
<intersection>-6247 3</intersection></vsegment></shape></wire>
<wire>
<ID>1321</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>435,-6238.5,444,-6238.5</points>
<connection>
<GID>1900</GID>
<name>OUT</name></connection>
<connection>
<GID>1905</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-6247,425.5,-6226.5</points>
<intersection>-6247 3</intersection>
<intersection>-6237.5 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,-6237.5,429,-6237.5</points>
<connection>
<GID>1900</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,-6226.5,425.5,-6226.5</points>
<connection>
<GID>1904</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>425.5,-6247,446,-6247</points>
<intersection>425.5 0</intersection>
<intersection>446 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>446,-6247,446,-6241.5</points>
<connection>
<GID>1905</GID>
<name>IN_0</name></connection>
<intersection>-6247 3</intersection></vsegment></shape></wire>
<wire>
<ID>1323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-6240.5,528.5,-6240.5</points>
<connection>
<GID>1909</GID>
<name>OUT</name></connection>
<connection>
<GID>1908</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,-6246.5,510,-6226.5</points>
<intersection>-6246.5 3</intersection>
<intersection>-6239.5 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,-6239.5,513,-6239.5</points>
<connection>
<GID>1909</GID>
<name>IN_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509,-6226.5,510,-6226.5</points>
<connection>
<GID>1907</GID>
<name>OUT_0</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>510,-6246.5,530.5,-6246.5</points>
<intersection>510 0</intersection>
<intersection>530.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>530.5,-6246.5,530.5,-6243.5</points>
<connection>
<GID>1908</GID>
<name>IN_0</name></connection>
<intersection>-6246.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1325</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>593,-6240.5,602,-6240.5</points>
<connection>
<GID>1906</GID>
<name>OUT</name></connection>
<connection>
<GID>1911</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,-6246.5,583.5,-6226.5</points>
<intersection>-6246.5 3</intersection>
<intersection>-6239.5 1</intersection>
<intersection>-6226.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583.5,-6239.5,587,-6239.5</points>
<connection>
<GID>1906</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>582.5,-6226.5,583.5,-6226.5</points>
<connection>
<GID>1910</GID>
<name>OUT_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>583.5,-6246.5,604,-6246.5</points>
<intersection>583.5 0</intersection>
<intersection>604 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>604,-6246.5,604,-6243.5</points>
<connection>
<GID>1911</GID>
<name>IN_0</name></connection>
<intersection>-6246.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3.5,-6229.5,576.5,-6229.5</points>
<connection>
<GID>1889</GID>
<name>clock</name></connection>
<connection>
<GID>1892</GID>
<name>clock</name></connection>
<connection>
<GID>1895</GID>
<name>clock</name></connection>
<connection>
<GID>1901</GID>
<name>clock</name></connection>
<connection>
<GID>1904</GID>
<name>clock</name></connection>
<connection>
<GID>1907</GID>
<name>clock</name></connection>
<connection>
<GID>1910</GID>
<name>clock</name></connection>
<connection>
<GID>1912</GID>
<name>OUT</name></connection>
<connection>
<GID>1898</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-6156.5,-111,-6098.5</points>
<intersection>-6156.5 3</intersection>
<intersection>-6138.5 1</intersection>
<intersection>-6098.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-6138.5,-12.5,-6138.5</points>
<connection>
<GID>1729</GID>
<name>IN_0</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6098.5,-111,-6098.5</points>
<connection>
<GID>1783</GID>
<name>OUT_3</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-111,-6156.5,-31,-6156.5</points>
<connection>
<GID>1730</GID>
<name>ENABLE_0</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>1329</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-28.5,-6158.5,584,-6158.5</points>
<connection>
<GID>1730</GID>
<name>OUT_0</name></connection>
<intersection>29 38</intersection>
<intersection>103 43</intersection>
<intersection>187 42</intersection>
<intersection>261 45</intersection>
<intersection>352 47</intersection>
<intersection>426 49</intersection>
<intersection>510 51</intersection>
<intersection>584 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>29,-6158.5,29,-6146</points>
<connection>
<GID>1917</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>187,-6158.5,187,-6148</points>
<connection>
<GID>1714</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>103,-6158.5,103,-6146</points>
<connection>
<GID>1914</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>261,-6158.5,261,-6148</points>
<connection>
<GID>1920</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>352,-6158.5,352,-6149.5</points>
<connection>
<GID>1720</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>426,-6158.5,426,-6149.5</points>
<connection>
<GID>1717</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>510,-6158.5,510,-6151.5</points>
<connection>
<GID>1726</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>584,-6158.5,584,-6151.5</points>
<connection>
<GID>1723</GID>
<name>IN_1</name></connection>
<intersection>-6158.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-6145,44.5,-6145</points>
<connection>
<GID>1917</GID>
<name>OUT</name></connection>
<connection>
<GID>1916</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-6153.5,26,-6136.5</points>
<intersection>-6153.5 3</intersection>
<intersection>-6144 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-6144,29,-6144</points>
<connection>
<GID>1917</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-6136.5,26,-6136.5</points>
<connection>
<GID>1915</GID>
<name>OUT_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26,-6153.5,46.5,-6153.5</points>
<intersection>26 0</intersection>
<intersection>46.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46.5,-6153.5,46.5,-6148</points>
<connection>
<GID>1916</GID>
<name>IN_0</name></connection>
<intersection>-6153.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1332</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>109,-6145,118,-6145</points>
<connection>
<GID>1914</GID>
<name>OUT</name></connection>
<connection>
<GID>1919</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-6155,99.5,-6136.5</points>
<intersection>-6155 3</intersection>
<intersection>-6144 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-6144,103,-6144</points>
<connection>
<GID>1914</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-6136.5,99.5,-6136.5</points>
<connection>
<GID>1918</GID>
<name>OUT_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-6155,120,-6155</points>
<intersection>99.5 0</intersection>
<intersection>120 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>120,-6155,120,-6148</points>
<connection>
<GID>1919</GID>
<name>IN_0</name></connection>
<intersection>-6155 3</intersection></vsegment></shape></wire>
<wire>
<ID>1334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>193,-6147,202.5,-6147</points>
<connection>
<GID>1714</GID>
<name>OUT</name></connection>
<connection>
<GID>1922</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-6155.5,184,-6136.5</points>
<intersection>-6155.5 3</intersection>
<intersection>-6146 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-6146,187,-6146</points>
<connection>
<GID>1714</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183,-6136.5,184,-6136.5</points>
<connection>
<GID>1921</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184,-6155.5,204.5,-6155.5</points>
<intersection>184 0</intersection>
<intersection>204.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>204.5,-6155.5,204.5,-6150</points>
<connection>
<GID>1922</GID>
<name>IN_0</name></connection>
<intersection>-6155.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1336</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>267,-6147,276,-6147</points>
<connection>
<GID>1920</GID>
<name>OUT</name></connection>
<connection>
<GID>1716</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-6157,257.5,-6136.5</points>
<connection>
<GID>1715</GID>
<name>OUT_0</name></connection>
<intersection>-6157 3</intersection>
<intersection>-6146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-6146,261,-6146</points>
<connection>
<GID>1920</GID>
<name>IN_0</name></connection>
<intersection>257.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257.5,-6157,278,-6157</points>
<intersection>257.5 0</intersection>
<intersection>278 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>278,-6157,278,-6150</points>
<connection>
<GID>1716</GID>
<name>IN_0</name></connection>
<intersection>-6157 3</intersection></vsegment></shape></wire>
<wire>
<ID>1338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358,-6148.5,367.5,-6148.5</points>
<connection>
<GID>1720</GID>
<name>OUT</name></connection>
<connection>
<GID>1719</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349,-6157,349,-6136.5</points>
<intersection>-6157 3</intersection>
<intersection>-6147.5 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349,-6147.5,352,-6147.5</points>
<connection>
<GID>1720</GID>
<name>IN_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348,-6136.5,349,-6136.5</points>
<connection>
<GID>1718</GID>
<name>OUT_0</name></connection>
<intersection>349 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>349,-6157,369.5,-6157</points>
<intersection>349 0</intersection>
<intersection>369.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>369.5,-6157,369.5,-6151.5</points>
<connection>
<GID>1719</GID>
<name>IN_0</name></connection>
<intersection>-6157 3</intersection></vsegment></shape></wire>
<wire>
<ID>1340</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>432,-6148.5,441,-6148.5</points>
<connection>
<GID>1717</GID>
<name>OUT</name></connection>
<connection>
<GID>1722</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422.5,-6157,422.5,-6136.5</points>
<intersection>-6157 3</intersection>
<intersection>-6147.5 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>422.5,-6147.5,426,-6147.5</points>
<connection>
<GID>1717</GID>
<name>IN_0</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,-6136.5,422.5,-6136.5</points>
<connection>
<GID>1721</GID>
<name>OUT_0</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>422.5,-6157,443,-6157</points>
<intersection>422.5 0</intersection>
<intersection>443 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>443,-6157,443,-6151.5</points>
<connection>
<GID>1722</GID>
<name>IN_0</name></connection>
<intersection>-6157 3</intersection></vsegment></shape></wire>
<wire>
<ID>1342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>516,-6150.5,525.5,-6150.5</points>
<connection>
<GID>1726</GID>
<name>OUT</name></connection>
<connection>
<GID>1725</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,-6156.5,507,-6136.5</points>
<intersection>-6156.5 3</intersection>
<intersection>-6149.5 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507,-6149.5,510,-6149.5</points>
<connection>
<GID>1726</GID>
<name>IN_0</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>506,-6136.5,507,-6136.5</points>
<connection>
<GID>1724</GID>
<name>OUT_0</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>507,-6156.5,527.5,-6156.5</points>
<intersection>507 0</intersection>
<intersection>527.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>527.5,-6156.5,527.5,-6153.5</points>
<connection>
<GID>1725</GID>
<name>IN_0</name></connection>
<intersection>-6156.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1344</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>590,-6150.5,599,-6150.5</points>
<connection>
<GID>1723</GID>
<name>OUT</name></connection>
<connection>
<GID>1728</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>580.5,-6156.5,580.5,-6136.5</points>
<intersection>-6156.5 3</intersection>
<intersection>-6149.5 1</intersection>
<intersection>-6136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>580.5,-6149.5,584,-6149.5</points>
<connection>
<GID>1723</GID>
<name>IN_0</name></connection>
<intersection>580.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>579.5,-6136.5,580.5,-6136.5</points>
<connection>
<GID>1727</GID>
<name>OUT_0</name></connection>
<intersection>580.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>580.5,-6156.5,601,-6156.5</points>
<intersection>580.5 0</intersection>
<intersection>601 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>601,-6156.5,601,-6153.5</points>
<connection>
<GID>1728</GID>
<name>IN_0</name></connection>
<intersection>-6156.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-6139.5,573.5,-6139.5</points>
<connection>
<GID>1921</GID>
<name>clock</name></connection>
<connection>
<GID>1918</GID>
<name>clock</name></connection>
<connection>
<GID>1915</GID>
<name>clock</name></connection>
<connection>
<GID>1729</GID>
<name>OUT</name></connection>
<connection>
<GID>1727</GID>
<name>clock</name></connection>
<connection>
<GID>1724</GID>
<name>clock</name></connection>
<connection>
<GID>1721</GID>
<name>clock</name></connection>
<connection>
<GID>1718</GID>
<name>clock</name></connection>
<connection>
<GID>1715</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-115,-6414.5,-115,-6101.5</points>
<intersection>-6414.5 3</intersection>
<intersection>-6396.5 1</intersection>
<intersection>-6101.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-115,-6396.5,-5.5,-6396.5</points>
<connection>
<GID>1755</GID>
<name>IN_0</name></connection>
<intersection>-115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6101.5,-115,-6101.5</points>
<connection>
<GID>1783</GID>
<name>OUT_0</name></connection>
<intersection>-115 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-115,-6414.5,-24,-6414.5</points>
<connection>
<GID>1756</GID>
<name>ENABLE_0</name></connection>
<intersection>-115 0</intersection></hsegment></shape></wire>
<wire>
<ID>1348</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-21.5,-6416.5,591,-6416.5</points>
<connection>
<GID>1756</GID>
<name>OUT_0</name></connection>
<intersection>36 38</intersection>
<intersection>110 43</intersection>
<intersection>194 42</intersection>
<intersection>268 45</intersection>
<intersection>359 47</intersection>
<intersection>433 49</intersection>
<intersection>517 51</intersection>
<intersection>591 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>36,-6416.5,36,-6404</points>
<connection>
<GID>1734</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>194,-6416.5,194,-6406</points>
<connection>
<GID>1740</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>110,-6416.5,110,-6404</points>
<connection>
<GID>1731</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>268,-6416.5,268,-6406</points>
<connection>
<GID>1737</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>359,-6416.5,359,-6407.5</points>
<connection>
<GID>1746</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>433,-6416.5,433,-6407.5</points>
<connection>
<GID>1743</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>517,-6416.5,517,-6409.5</points>
<connection>
<GID>1752</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>591,-6416.5,591,-6409.5</points>
<connection>
<GID>1749</GID>
<name>IN_1</name></connection>
<intersection>-6416.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-6403,51.5,-6403</points>
<connection>
<GID>1734</GID>
<name>OUT</name></connection>
<connection>
<GID>1733</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-6411.5,33,-6394.5</points>
<intersection>-6411.5 3</intersection>
<intersection>-6402 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-6402,36,-6402</points>
<connection>
<GID>1734</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-6394.5,33,-6394.5</points>
<connection>
<GID>1732</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-6411.5,53.5,-6411.5</points>
<intersection>33 0</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-6411.5,53.5,-6406</points>
<connection>
<GID>1733</GID>
<name>IN_0</name></connection>
<intersection>-6411.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1351</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116,-6403,125,-6403</points>
<connection>
<GID>1731</GID>
<name>OUT</name></connection>
<connection>
<GID>1736</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-6413,106.5,-6394.5</points>
<intersection>-6413 3</intersection>
<intersection>-6402 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-6402,110,-6402</points>
<connection>
<GID>1731</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-6394.5,106.5,-6394.5</points>
<connection>
<GID>1735</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,-6413,127,-6413</points>
<intersection>106.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-6413,127,-6406</points>
<connection>
<GID>1736</GID>
<name>IN_0</name></connection>
<intersection>-6413 3</intersection></vsegment></shape></wire>
<wire>
<ID>1353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-6405,209.5,-6405</points>
<connection>
<GID>1740</GID>
<name>OUT</name></connection>
<connection>
<GID>1739</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-6413.5,191,-6394.5</points>
<intersection>-6413.5 3</intersection>
<intersection>-6404 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-6404,194,-6404</points>
<connection>
<GID>1740</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,-6394.5,191,-6394.5</points>
<connection>
<GID>1738</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191,-6413.5,211.5,-6413.5</points>
<intersection>191 0</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>211.5,-6413.5,211.5,-6408</points>
<connection>
<GID>1739</GID>
<name>IN_0</name></connection>
<intersection>-6413.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1355</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>274,-6405,283,-6405</points>
<connection>
<GID>1737</GID>
<name>OUT</name></connection>
<connection>
<GID>1742</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-6415,264.5,-6394.5</points>
<connection>
<GID>1741</GID>
<name>OUT_0</name></connection>
<intersection>-6415 3</intersection>
<intersection>-6404 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-6404,268,-6404</points>
<connection>
<GID>1737</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>264.5,-6415,285,-6415</points>
<intersection>264.5 0</intersection>
<intersection>285 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>285,-6415,285,-6408</points>
<connection>
<GID>1742</GID>
<name>IN_0</name></connection>
<intersection>-6415 3</intersection></vsegment></shape></wire>
<wire>
<ID>1357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365,-6406.5,374.5,-6406.5</points>
<connection>
<GID>1746</GID>
<name>OUT</name></connection>
<connection>
<GID>1745</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356,-6415,356,-6394.5</points>
<intersection>-6415 3</intersection>
<intersection>-6405.5 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-6405.5,359,-6405.5</points>
<connection>
<GID>1746</GID>
<name>IN_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>355,-6394.5,356,-6394.5</points>
<connection>
<GID>1744</GID>
<name>OUT_0</name></connection>
<intersection>356 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>356,-6415,376.5,-6415</points>
<intersection>356 0</intersection>
<intersection>376.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>376.5,-6415,376.5,-6409.5</points>
<connection>
<GID>1745</GID>
<name>IN_0</name></connection>
<intersection>-6415 3</intersection></vsegment></shape></wire>
<wire>
<ID>1359</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>439,-6406.5,448,-6406.5</points>
<connection>
<GID>1743</GID>
<name>OUT</name></connection>
<connection>
<GID>1748</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-6415,429.5,-6394.5</points>
<intersection>-6415 3</intersection>
<intersection>-6405.5 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,-6405.5,433,-6405.5</points>
<connection>
<GID>1743</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,-6394.5,429.5,-6394.5</points>
<connection>
<GID>1747</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,-6415,450,-6415</points>
<intersection>429.5 0</intersection>
<intersection>450 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>450,-6415,450,-6409.5</points>
<connection>
<GID>1748</GID>
<name>IN_0</name></connection>
<intersection>-6415 3</intersection></vsegment></shape></wire>
<wire>
<ID>1361</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523,-6408.5,532.5,-6408.5</points>
<connection>
<GID>1752</GID>
<name>OUT</name></connection>
<connection>
<GID>1751</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-6414.5,514,-6394.5</points>
<intersection>-6414.5 3</intersection>
<intersection>-6407.5 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-6407.5,517,-6407.5</points>
<connection>
<GID>1752</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513,-6394.5,514,-6394.5</points>
<connection>
<GID>1750</GID>
<name>OUT_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>514,-6414.5,534.5,-6414.5</points>
<intersection>514 0</intersection>
<intersection>534.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>534.5,-6414.5,534.5,-6411.5</points>
<connection>
<GID>1751</GID>
<name>IN_0</name></connection>
<intersection>-6414.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1363</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>597,-6408.5,606,-6408.5</points>
<connection>
<GID>1749</GID>
<name>OUT</name></connection>
<connection>
<GID>1754</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,-6414.5,587.5,-6394.5</points>
<intersection>-6414.5 3</intersection>
<intersection>-6407.5 1</intersection>
<intersection>-6394.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>587.5,-6407.5,591,-6407.5</points>
<connection>
<GID>1749</GID>
<name>IN_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>586.5,-6394.5,587.5,-6394.5</points>
<connection>
<GID>1753</GID>
<name>OUT_0</name></connection>
<intersection>587.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>587.5,-6414.5,608,-6414.5</points>
<intersection>587.5 0</intersection>
<intersection>608 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>608,-6414.5,608,-6411.5</points>
<connection>
<GID>1754</GID>
<name>IN_0</name></connection>
<intersection>-6414.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-6397.5,580.5,-6397.5</points>
<connection>
<GID>1732</GID>
<name>clock</name></connection>
<connection>
<GID>1735</GID>
<name>clock</name></connection>
<connection>
<GID>1738</GID>
<name>clock</name></connection>
<connection>
<GID>1744</GID>
<name>clock</name></connection>
<connection>
<GID>1747</GID>
<name>clock</name></connection>
<connection>
<GID>1750</GID>
<name>clock</name></connection>
<connection>
<GID>1753</GID>
<name>clock</name></connection>
<connection>
<GID>1755</GID>
<name>OUT</name></connection>
<connection>
<GID>1741</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113,-6324.5,-113,-6100.5</points>
<intersection>-6324.5 3</intersection>
<intersection>-6306.5 1</intersection>
<intersection>-6100.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-113,-6306.5,-8.5,-6306.5</points>
<connection>
<GID>1781</GID>
<name>IN_0</name></connection>
<intersection>-113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121.5,-6100.5,-113,-6100.5</points>
<connection>
<GID>1783</GID>
<name>OUT_1</name></connection>
<intersection>-113 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-113,-6324.5,-27,-6324.5</points>
<connection>
<GID>1782</GID>
<name>ENABLE_0</name></connection>
<intersection>-113 0</intersection></hsegment></shape></wire>
<wire>
<ID>1367</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-24.5,-6326.5,588,-6326.5</points>
<connection>
<GID>1782</GID>
<name>OUT_0</name></connection>
<intersection>33 38</intersection>
<intersection>107 43</intersection>
<intersection>191 42</intersection>
<intersection>265 45</intersection>
<intersection>356 47</intersection>
<intersection>430 49</intersection>
<intersection>514 51</intersection>
<intersection>588 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>33,-6326.5,33,-6314</points>
<connection>
<GID>1760</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>191,-6326.5,191,-6316</points>
<connection>
<GID>1766</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>107,-6326.5,107,-6314</points>
<connection>
<GID>1757</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>265,-6326.5,265,-6316</points>
<connection>
<GID>1763</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>356,-6326.5,356,-6317.5</points>
<connection>
<GID>1772</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>430,-6326.5,430,-6317.5</points>
<connection>
<GID>1769</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>514,-6326.5,514,-6319.5</points>
<connection>
<GID>1778</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>588,-6326.5,588,-6319.5</points>
<connection>
<GID>1775</GID>
<name>IN_1</name></connection>
<intersection>-6326.5 33</intersection></vsegment></shape></wire>
<wire>
<ID>1368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-6313,48.5,-6313</points>
<connection>
<GID>1760</GID>
<name>OUT</name></connection>
<connection>
<GID>1759</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-6321.5,30,-6304.5</points>
<intersection>-6321.5 3</intersection>
<intersection>-6312 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-6312,33,-6312</points>
<connection>
<GID>1760</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-6304.5,30,-6304.5</points>
<connection>
<GID>1758</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30,-6321.5,50.5,-6321.5</points>
<intersection>30 0</intersection>
<intersection>50.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50.5,-6321.5,50.5,-6316</points>
<connection>
<GID>1759</GID>
<name>IN_0</name></connection>
<intersection>-6321.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1370</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113,-6313,122,-6313</points>
<connection>
<GID>1757</GID>
<name>OUT</name></connection>
<connection>
<GID>1762</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-6323,103.5,-6304.5</points>
<intersection>-6323 3</intersection>
<intersection>-6312 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-6312,107,-6312</points>
<connection>
<GID>1757</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-6304.5,103.5,-6304.5</points>
<connection>
<GID>1761</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,-6323,124,-6323</points>
<intersection>103.5 0</intersection>
<intersection>124 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124,-6323,124,-6316</points>
<connection>
<GID>1762</GID>
<name>IN_0</name></connection>
<intersection>-6323 3</intersection></vsegment></shape></wire>
<wire>
<ID>1372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-6315,206.5,-6315</points>
<connection>
<GID>1766</GID>
<name>OUT</name></connection>
<connection>
<GID>1765</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-6323.5,188,-6304.5</points>
<intersection>-6323.5 3</intersection>
<intersection>-6314 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188,-6314,191,-6314</points>
<connection>
<GID>1766</GID>
<name>IN_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-6304.5,188,-6304.5</points>
<connection>
<GID>1764</GID>
<name>OUT_0</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188,-6323.5,208.5,-6323.5</points>
<intersection>188 0</intersection>
<intersection>208.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>208.5,-6323.5,208.5,-6318</points>
<connection>
<GID>1765</GID>
<name>IN_0</name></connection>
<intersection>-6323.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1374</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>271,-6315,280,-6315</points>
<connection>
<GID>1763</GID>
<name>OUT</name></connection>
<connection>
<GID>1768</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-6325,261.5,-6304.5</points>
<connection>
<GID>1767</GID>
<name>OUT_0</name></connection>
<intersection>-6325 3</intersection>
<intersection>-6314 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-6314,265,-6314</points>
<connection>
<GID>1763</GID>
<name>IN_0</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>261.5,-6325,282,-6325</points>
<intersection>261.5 0</intersection>
<intersection>282 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282,-6325,282,-6318</points>
<connection>
<GID>1768</GID>
<name>IN_0</name></connection>
<intersection>-6325 3</intersection></vsegment></shape></wire>
<wire>
<ID>1376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362,-6316.5,371.5,-6316.5</points>
<connection>
<GID>1772</GID>
<name>OUT</name></connection>
<connection>
<GID>1771</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-6325,353,-6304.5</points>
<intersection>-6325 3</intersection>
<intersection>-6315.5 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>353,-6315.5,356,-6315.5</points>
<connection>
<GID>1772</GID>
<name>IN_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-6304.5,353,-6304.5</points>
<connection>
<GID>1770</GID>
<name>OUT_0</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353,-6325,373.5,-6325</points>
<intersection>353 0</intersection>
<intersection>373.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>373.5,-6325,373.5,-6319.5</points>
<connection>
<GID>1771</GID>
<name>IN_0</name></connection>
<intersection>-6325 3</intersection></vsegment></shape></wire>
<wire>
<ID>1378</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>436,-6316.5,445,-6316.5</points>
<connection>
<GID>1769</GID>
<name>OUT</name></connection>
<connection>
<GID>1774</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-6325,426.5,-6304.5</points>
<intersection>-6325 3</intersection>
<intersection>-6315.5 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426.5,-6315.5,430,-6315.5</points>
<connection>
<GID>1769</GID>
<name>IN_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>425.5,-6304.5,426.5,-6304.5</points>
<connection>
<GID>1773</GID>
<name>OUT_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>426.5,-6325,447,-6325</points>
<intersection>426.5 0</intersection>
<intersection>447 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447,-6325,447,-6319.5</points>
<connection>
<GID>1774</GID>
<name>IN_0</name></connection>
<intersection>-6325 3</intersection></vsegment></shape></wire>
<wire>
<ID>1380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>520,-6318.5,529.5,-6318.5</points>
<connection>
<GID>1778</GID>
<name>OUT</name></connection>
<connection>
<GID>1777</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,-6324.5,511,-6304.5</points>
<intersection>-6324.5 3</intersection>
<intersection>-6317.5 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,-6317.5,514,-6317.5</points>
<connection>
<GID>1778</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>510,-6304.5,511,-6304.5</points>
<connection>
<GID>1776</GID>
<name>OUT_0</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511,-6324.5,531.5,-6324.5</points>
<intersection>511 0</intersection>
<intersection>531.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531.5,-6324.5,531.5,-6321.5</points>
<connection>
<GID>1777</GID>
<name>IN_0</name></connection>
<intersection>-6324.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1382</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>594,-6318.5,603,-6318.5</points>
<connection>
<GID>1775</GID>
<name>OUT</name></connection>
<connection>
<GID>1780</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584.5,-6324.5,584.5,-6304.5</points>
<intersection>-6324.5 3</intersection>
<intersection>-6317.5 1</intersection>
<intersection>-6304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>584.5,-6317.5,588,-6317.5</points>
<connection>
<GID>1775</GID>
<name>IN_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583.5,-6304.5,584.5,-6304.5</points>
<connection>
<GID>1779</GID>
<name>OUT_0</name></connection>
<intersection>584.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>584.5,-6324.5,605,-6324.5</points>
<intersection>584.5 0</intersection>
<intersection>605 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>605,-6324.5,605,-6321.5</points>
<connection>
<GID>1780</GID>
<name>IN_0</name></connection>
<intersection>-6324.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1384</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-6307.5,577.5,-6307.5</points>
<connection>
<GID>1758</GID>
<name>clock</name></connection>
<connection>
<GID>1761</GID>
<name>clock</name></connection>
<connection>
<GID>1764</GID>
<name>clock</name></connection>
<connection>
<GID>1770</GID>
<name>clock</name></connection>
<connection>
<GID>1773</GID>
<name>clock</name></connection>
<connection>
<GID>1776</GID>
<name>clock</name></connection>
<connection>
<GID>1779</GID>
<name>clock</name></connection>
<connection>
<GID>1781</GID>
<name>OUT</name></connection>
<connection>
<GID>1767</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-170,39,-122.5,39</points>
<intersection>-170 15</intersection>
<intersection>-130 6</intersection>
<intersection>-122.5 14</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-130,-6099.5,-130,39</points>
<intersection>-6099.5 7</intersection>
<intersection>-5228 13</intersection>
<intersection>-4303.5 12</intersection>
<intersection>-3478 11</intersection>
<intersection>-2584 10</intersection>
<intersection>-1712.5 9</intersection>
<intersection>-788 8</intersection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-130,-6099.5,-127.5,-6099.5</points>
<connection>
<GID>1783</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-130,-788,-122.5,-788</points>
<connection>
<GID>529</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-130,-1712.5,-125,-1712.5</points>
<connection>
<GID>738</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-130,-2584,-125.5,-2584</points>
<connection>
<GID>947</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-130,-3478,-124.5,-3478</points>
<connection>
<GID>1295</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-130,-4303.5,-124.5,-4303.5</points>
<connection>
<GID>1365</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-130,-5228,-127,-5228</points>
<connection>
<GID>1574</GID>
<name>IN_2</name></connection>
<intersection>-130 6</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-122.5,37.5,-122.5,39</points>
<connection>
<GID>459</GID>
<name>IN_2</name></connection>
<intersection>39 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-170,39,-170,42</points>
<connection>
<GID>1926</GID>
<name>OUT_0</name></connection>
<intersection>39 1</intersection></vsegment></shape></wire>
<wire>
<ID>1386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-170,36.5,-122.5,36.5</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<connection>
<GID>1928</GID>
<name>OUT_0</name></connection>
<intersection>-129 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-129,-6100.5,-129,36.5</points>
<intersection>-6100.5 9</intersection>
<intersection>-5229 14</intersection>
<intersection>-4304.5 13</intersection>
<intersection>-3479 12</intersection>
<intersection>-2585 11</intersection>
<intersection>-1713.5 10</intersection>
<intersection>-789 8</intersection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-129,-789,-122.5,-789</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-129,-6100.5,-127.5,-6100.5</points>
<connection>
<GID>1783</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-129,-1713.5,-125,-1713.5</points>
<connection>
<GID>738</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-129,-2585,-125.5,-2585</points>
<connection>
<GID>947</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-129,-3479,-124.5,-3479</points>
<connection>
<GID>1295</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-129,-4304.5,-124.5,-4304.5</points>
<connection>
<GID>1365</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-129,-5229,-127,-5229</points>
<connection>
<GID>1574</GID>
<name>IN_1</name></connection>
<intersection>-129 7</intersection></hsegment></shape></wire>
<wire>
<ID>1387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-128,-6101.5,-128,35.5</points>
<intersection>-6101.5 3</intersection>
<intersection>-5230 9</intersection>
<intersection>-4305.5 8</intersection>
<intersection>-3480 7</intersection>
<intersection>-2586 6</intersection>
<intersection>-1714.5 5</intersection>
<intersection>-790 4</intersection>
<intersection>30 1</intersection>
<intersection>35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-170,30,-128,30</points>
<connection>
<GID>1930</GID>
<name>OUT_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-128,35.5,-122.5,35.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-128,-6101.5,-127.5,-6101.5</points>
<connection>
<GID>1783</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-128,-790,-122.5,-790</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,-1714.5,-125,-1714.5</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-128,-2586,-125.5,-2586</points>
<connection>
<GID>947</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-128,-3480,-124.5,-3480</points>
<connection>
<GID>1295</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-128,-4305.5,-124.5,-4305.5</points>
<connection>
<GID>1365</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-128,-5230,-127,-5230</points>
<connection>
<GID>1574</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment></shape></wire>
<wire>
<ID>1389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-170,21,-147,21</points>
<connection>
<GID>1935</GID>
<name>IN_2</name></connection>
<connection>
<GID>1937</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-149,16.5,-149,20</points>
<intersection>16.5 2</intersection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-149,20,-147,20</points>
<connection>
<GID>1935</GID>
<name>IN_1</name></connection>
<intersection>-149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-170.5,16.5,-149,16.5</points>
<connection>
<GID>1939</GID>
<name>OUT_0</name></connection>
<intersection>-149 0</intersection></hsegment></shape></wire>
<wire>
<ID>1391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148,12,-148,19</points>
<intersection>12 2</intersection>
<intersection>19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-148,19,-147,19</points>
<connection>
<GID>1935</GID>
<name>IN_0</name></connection>
<intersection>-148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-170,12,-148,12</points>
<connection>
<GID>1941</GID>
<name>OUT_0</name></connection>
<intersection>-148 0</intersection></hsegment></shape></wire>
<wire>
<ID>1392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-150.5,26,-147,26</points>
<connection>
<GID>1935</GID>
<name>ENABLE</name></connection>
<connection>
<GID>1943</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-134,26,-134,42.5</points>
<intersection>26 1</intersection>
<intersection>42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-141,26,-134,26</points>
<connection>
<GID>1935</GID>
<name>OUT_7</name></connection>
<intersection>-134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-134,42.5,-122.5,42.5</points>
<connection>
<GID>459</GID>
<name>ENABLE</name></connection>
<intersection>-134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-134,-783,-134,25</points>
<intersection>-783 1</intersection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-134,-783,-122.5,-783</points>
<connection>
<GID>529</GID>
<name>ENABLE</name></connection>
<intersection>-134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-141,25,-134,25</points>
<connection>
<GID>1935</GID>
<name>OUT_6</name></connection>
<intersection>-134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-135,-1707.5,-135,24</points>
<intersection>-1707.5 2</intersection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-141,24,-135,24</points>
<connection>
<GID>1935</GID>
<name>OUT_5</name></connection>
<intersection>-135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-135,-1707.5,-125,-1707.5</points>
<connection>
<GID>738</GID>
<name>ENABLE</name></connection>
<intersection>-135 0</intersection></hsegment></shape></wire>
<wire>
<ID>1396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-136,-2579,-136,23</points>
<intersection>-2579 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136,-2579,-125.5,-2579</points>
<connection>
<GID>947</GID>
<name>ENABLE</name></connection>
<intersection>-136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-141,23,-136,23</points>
<connection>
<GID>1935</GID>
<name>OUT_4</name></connection>
<intersection>-136 0</intersection></hsegment></shape></wire>
<wire>
<ID>1397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-137,-3473,-137,22</points>
<intersection>-3473 2</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-141,22,-137,22</points>
<connection>
<GID>1935</GID>
<name>OUT_3</name></connection>
<intersection>-137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-137,-3473,-124.5,-3473</points>
<connection>
<GID>1295</GID>
<name>ENABLE</name></connection>
<intersection>-137 0</intersection></hsegment></shape></wire>
<wire>
<ID>1398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-138,-4298.5,-138,21</points>
<intersection>-4298.5 1</intersection>
<intersection>21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-138,-4298.5,-124.5,-4298.5</points>
<connection>
<GID>1365</GID>
<name>ENABLE</name></connection>
<intersection>-138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-141,21,-138,21</points>
<connection>
<GID>1935</GID>
<name>OUT_2</name></connection>
<intersection>-138 0</intersection></hsegment></shape></wire>
<wire>
<ID>1399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-139,-5223,-139,20</points>
<intersection>-5223 1</intersection>
<intersection>20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-139,-5223,-127,-5223</points>
<connection>
<GID>1574</GID>
<name>ENABLE</name></connection>
<intersection>-139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-141,20,-139,20</points>
<connection>
<GID>1935</GID>
<name>OUT_1</name></connection>
<intersection>-139 0</intersection></hsegment></shape></wire>
<wire>
<ID>1400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-140,-6094.5,-140,19</points>
<intersection>-6094.5 2</intersection>
<intersection>19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-141,19,-140,19</points>
<connection>
<GID>1935</GID>
<name>OUT_0</name></connection>
<intersection>-140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-140,-6094.5,-127.5,-6094.5</points>
<connection>
<GID>1783</GID>
<name>ENABLE</name></connection>
<intersection>-140 0</intersection></hsegment></shape></wire>
<wire>
<ID>1403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-281.5,62,-281.5,66</points>
<connection>
<GID>2003</GID>
<name>N_in3</name></connection>
<connection>
<GID>2066</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-271,62,-271,66</points>
<connection>
<GID>2004</GID>
<name>N_in3</name></connection>
<connection>
<GID>2068</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-261,62,-261,66</points>
<connection>
<GID>2005</GID>
<name>N_in3</name></connection>
<connection>
<GID>2070</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-253.5,62,-253.5,66</points>
<connection>
<GID>2006</GID>
<name>N_in3</name></connection>
<connection>
<GID>2072</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-242,62,-242,66</points>
<connection>
<GID>2007</GID>
<name>N_in3</name></connection>
<connection>
<GID>2074</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233,62,-233,66</points>
<connection>
<GID>2024</GID>
<name>N_in3</name></connection>
<connection>
<GID>2076</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-223,62,-223,66</points>
<connection>
<GID>2022</GID>
<name>N_in3</name></connection>
<connection>
<GID>2078</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-215,62,-215,66</points>
<connection>
<GID>2026</GID>
<name>N_in3</name></connection>
<connection>
<GID>2080</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-6448.5,-15.5,372.5</points>
<intersection>-6448.5 3</intersection>
<intersection>-6398.5 1</intersection>
<intersection>-6308.5 69</intersection>
<intersection>-6230.5 68</intersection>
<intersection>-6140.5 67</intersection>
<intersection>-6022.5 66</intersection>
<intersection>-5932.5 65</intersection>
<intersection>-5854.5 64</intersection>
<intersection>-5764.5 63</intersection>
<intersection>-5527 62</intersection>
<intersection>-5437 61</intersection>
<intersection>-5359 60</intersection>
<intersection>-5269 59</intersection>
<intersection>-5151 58</intersection>
<intersection>-5061 51</intersection>
<intersection>-4983 50</intersection>
<intersection>-4893 49</intersection>
<intersection>-4602.5 48</intersection>
<intersection>-4512.5 47</intersection>
<intersection>-4434.5 46</intersection>
<intersection>-4344.5 45</intersection>
<intersection>-4226.5 44</intersection>
<intersection>-4136.5 43</intersection>
<intersection>-4058.5 42</intersection>
<intersection>-3968.5 41</intersection>
<intersection>-3777 40</intersection>
<intersection>-3687 39</intersection>
<intersection>-3609 38</intersection>
<intersection>-3519 37</intersection>
<intersection>-3401 36</intersection>
<intersection>-3311 35</intersection>
<intersection>-3233 34</intersection>
<intersection>-3143 33</intersection>
<intersection>-2883 32</intersection>
<intersection>-2793 31</intersection>
<intersection>-2715 30</intersection>
<intersection>-2625 29</intersection>
<intersection>-2507 28</intersection>
<intersection>-2339 27</intersection>
<intersection>-2249 26</intersection>
<intersection>-2011.5 25</intersection>
<intersection>-1921.5 24</intersection>
<intersection>-1843.5 23</intersection>
<intersection>-1753.5 22</intersection>
<intersection>-1545.5 21</intersection>
<intersection>-1467.5 20</intersection>
<intersection>-1377.5 19</intersection>
<intersection>-1087 18</intersection>
<intersection>-997 17</intersection>
<intersection>-919 16</intersection>
<intersection>-829 15</intersection>
<intersection>-711 14</intersection>
<intersection>-621 13</intersection>
<intersection>-543 12</intersection>
<intersection>-453 11</intersection>
<intersection>-261.5 10</intersection>
<intersection>-171.5 9</intersection>
<intersection>-93.5 8</intersection>
<intersection>-3.5 7</intersection>
<intersection>114.5 6</intersection>
<intersection>204.5 5</intersection>
<intersection>282.5 4</intersection>
<intersection>372.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-6398.5,-5.5,-6398.5</points>
<connection>
<GID>1755</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,372.5,-9.5,372.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-15.5,-6448.5,-8,-6448.5</points>
<connection>
<GID>2084</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-15.5,282.5,-6.5,282.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-15.5,204.5,-5.5,204.5</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-15.5,114.5,-2.5,114.5</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-15.5,-3.5,-7.5,-3.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-15.5,-93.5,-4.5,-93.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-15.5,-171.5,-3.5,-171.5</points>
<connection>
<GID>456</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-15.5,-261.5,-0.5,-261.5</points>
<connection>
<GID>430</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-15.5,-453,-9.5,-453</points>
<connection>
<GID>580</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-15.5,-543,-6.5,-543</points>
<connection>
<GID>554</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-15.5,-621,-5.5,-621</points>
<connection>
<GID>632</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-15.5,-711,-2.5,-711</points>
<connection>
<GID>606</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-15.5,-829,-7.5,-829</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-15.5,-919,-4.5,-919</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-15.5,-997,-3.5,-997</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-15.5,-1087,-0.5,-1087</points>
<connection>
<GID>501</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-15.5,-1377.5,-12,-1377.5</points>
<connection>
<GID>789</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-15.5,-1467.5,-9,-1467.5</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-15.5,-1545.5,-8,-1545.5</points>
<connection>
<GID>841</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-15.5,-1753.5,-10,-1753.5</points>
<connection>
<GID>684</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-15.5,-1843.5,-7,-1843.5</points>
<connection>
<GID>867</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-15.5,-1921.5,-6,-1921.5</points>
<connection>
<GID>736</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-15.5,-2011.5,-3,-2011.5</points>
<connection>
<GID>710</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-15.5,-2249,-12.5,-2249</points>
<connection>
<GID>998</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-15.5,-2339,-9.5,-2339</points>
<connection>
<GID>972</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-15.5,-2507,-5.5,-2507</points>
<connection>
<GID>1024</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-15.5,-2625,-10.5,-2625</points>
<connection>
<GID>893</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-15.5,-2715,-7.5,-2715</points>
<connection>
<GID>1076</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-15.5,-2793,-6.5,-2793</points>
<connection>
<GID>945</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-15.5,-2883,-3.5,-2883</points>
<connection>
<GID>919</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>-15.5,-3143,-11.5,-3143</points>
<connection>
<GID>1137</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-15.5,-3233,-8.5,-3233</points>
<connection>
<GID>1111</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-15.5,-3311,-7.5,-3311</points>
<connection>
<GID>1189</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-15.5,-3401,-4.5,-3401</points>
<connection>
<GID>1163</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-15.5,-3519,-9.5,-3519</points>
<connection>
<GID>1241</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>-15.5,-3609,-6.5,-3609</points>
<connection>
<GID>1215</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-15.5,-3687,-5.5,-3687</points>
<connection>
<GID>1293</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>-15.5,-3777,-2.5,-3777</points>
<connection>
<GID>1267</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>-15.5,-3968.5,-11.5,-3968.5</points>
<connection>
<GID>1416</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>-15.5,-4058.5,-8.5,-4058.5</points>
<connection>
<GID>1390</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>-15.5,-4136.5,-7.5,-4136.5</points>
<connection>
<GID>1468</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>-15.5,-4226.5,-4.5,-4226.5</points>
<connection>
<GID>1442</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-15.5,-4344.5,-9.5,-4344.5</points>
<connection>
<GID>1311</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>-15.5,-4434.5,-6.5,-4434.5</points>
<connection>
<GID>1494</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>-15.5,-4512.5,-5.5,-4512.5</points>
<connection>
<GID>1363</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-15.5,-4602.5,-2.5,-4602.5</points>
<connection>
<GID>1337</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>-15.5,-4893,-14,-4893</points>
<connection>
<GID>1625</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-15.5,-4983,-11,-4983</points>
<connection>
<GID>1599</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>-15.5,-5061,-10,-5061</points>
<connection>
<GID>1677</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>-15.5,-5151,-7,-5151</points>
<connection>
<GID>1651</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>-15.5,-5269,-12,-5269</points>
<connection>
<GID>1520</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>-15.5,-5359,-9,-5359</points>
<connection>
<GID>1703</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>-15.5,-5437,-8,-5437</points>
<connection>
<GID>1572</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>-15.5,-5527,-5,-5527</points>
<connection>
<GID>1546</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>-15.5,-5764.5,-14.5,-5764.5</points>
<connection>
<GID>1834</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>-15.5,-5854.5,-11.5,-5854.5</points>
<connection>
<GID>1808</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>-15.5,-5932.5,-10.5,-5932.5</points>
<connection>
<GID>1886</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>-15.5,-6022.5,-7.5,-6022.5</points>
<connection>
<GID>1860</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>-15.5,-6140.5,-12.5,-6140.5</points>
<connection>
<GID>1729</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>-15.5,-6230.5,-9.5,-6230.5</points>
<connection>
<GID>1912</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>-15.5,-6308.5,-8.5,-6308.5</points>
<connection>
<GID>1781</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-301,29,-297.5,29</points>
<connection>
<GID>2028</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2086</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-301,20.5,-298,20.5</points>
<connection>
<GID>2032</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2087</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-301,13,-298.5,13</points>
<connection>
<GID>2030</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2088</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-283,-13,-283,-10</points>
<connection>
<GID>1972</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2089</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-262.5,-13,-262.5,-10</points>
<connection>
<GID>1974</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2091</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-13,-255,-10</points>
<connection>
<GID>1975</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2092</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-244,-13.5,-244,-10.5</points>
<connection>
<GID>1961</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2093</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233,-13,-233,-10</points>
<connection>
<GID>1963</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2094</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-223,-13,-223,-10</points>
<connection>
<GID>1964</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2095</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-215,-13,-215,-10</points>
<connection>
<GID>1965</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2096</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-272.5,-13,-272.5,-10</points>
<connection>
<GID>1973</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2090</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-6452,13,-6444</points>
<connection>
<GID>2098</GID>
<name>IN_0</name></connection>
<connection>
<GID>2100</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-6453,75.5,-6444.5</points>
<connection>
<GID>2102</GID>
<name>IN_0</name></connection>
<connection>
<GID>2101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-6456,152,-6444.5</points>
<connection>
<GID>2104</GID>
<name>IN_0</name></connection>
<connection>
<GID>2103</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-6455.5,234.5,-6444.5</points>
<connection>
<GID>2105</GID>
<name>IN_0</name></connection>
<connection>
<GID>2106</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-6456,308,-6445</points>
<connection>
<GID>2107</GID>
<name>IN_0</name></connection>
<connection>
<GID>2108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,-6456,397,-6445</points>
<connection>
<GID>2110</GID>
<name>IN_0</name></connection>
<intersection>-6445 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>396.5,-6445,397,-6445</points>
<intersection>396.5 4</intersection>
<intersection>397 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>396.5,-6445.5,396.5,-6445</points>
<connection>
<GID>2109</GID>
<name>IN_0</name></connection>
<intersection>-6445 3</intersection></vsegment></shape></wire>
<wire>
<ID>1441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>478,-6456.5,478,-6445.5</points>
<connection>
<GID>2111</GID>
<name>IN_0</name></connection>
<connection>
<GID>2112</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>562,-6456.5,562,-6445.5</points>
<connection>
<GID>2113</GID>
<name>IN_0</name></connection>
<connection>
<GID>2114</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1444</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-6445.5,560,-6445.5</points>
<intersection>7.5 16</intersection>
<intersection>73.5 24</intersection>
<intersection>150 23</intersection>
<intersection>232.5 22</intersection>
<intersection>306 11</intersection>
<intersection>394.5 6</intersection>
<intersection>476 5</intersection>
<intersection>560 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>560,-6445.5,560,-6442.5</points>
<connection>
<GID>2113</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>476,-6445.5,476,-6442.5</points>
<connection>
<GID>2111</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>394.5,-6445.5,394.5,-6442.5</points>
<connection>
<GID>2109</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>306,-6445.5,306,-6442</points>
<connection>
<GID>2107</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>7.5,-6445.5,7.5,-6441</points>
<intersection>-6445.5 1</intersection>
<intersection>-6442 20</intersection>
<intersection>-6441 25</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>5.5,-6442,7.5,-6442</points>
<intersection>5.5 21</intersection>
<intersection>7.5 16</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>5.5,-6442,5.5,-6441</points>
<connection>
<GID>2116</GID>
<name>IN_0</name></connection>
<intersection>-6442 20</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>232.5,-6445.5,232.5,-6441.5</points>
<connection>
<GID>2105</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>150,-6445.5,150,-6441.5</points>
<connection>
<GID>2103</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>73.5,-6445.5,73.5,-6441.5</points>
<connection>
<GID>2101</GID>
<name>ENABLE_0</name></connection>
<intersection>-6445.5 1</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>7.5,-6441,11,-6441</points>
<connection>
<GID>2098</GID>
<name>ENABLE_0</name></connection>
<intersection>7.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>1445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,429,63,446.5</points>
<connection>
<GID>2118</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2127</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,428.5,143.5,445.5</points>
<connection>
<GID>2119</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,430.5,220,444.5</points>
<connection>
<GID>2132</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,429,288,446</points>
<connection>
<GID>2134</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,431,379.5,448</points>
<connection>
<GID>2136</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2137</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,430,458.5,447</points>
<connection>
<GID>2138</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543.5,427,543.5,444</points>
<connection>
<GID>2140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619.5,427.5,619.5,444.5</points>
<connection>
<GID>2144</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2145</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,433.5,617.5,433.5</points>
<intersection>61 15</intersection>
<intersection>141.5 13</intersection>
<intersection>218 11</intersection>
<intersection>286 9</intersection>
<intersection>377.5 5</intersection>
<intersection>456.5 3</intersection>
<intersection>541.5 6</intersection>
<intersection>617.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>456.5,427.5,456.5,433.5</points>
<connection>
<GID>2138</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>377.5,428.5,377.5,433.5</points>
<connection>
<GID>2136</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>541.5,424.5,541.5,433.5</points>
<connection>
<GID>2140</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>617.5,425,617.5,433.5</points>
<connection>
<GID>2144</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>286,426.5,286,433.5</points>
<connection>
<GID>2134</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>218,428,218,433.5</points>
<connection>
<GID>2132</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>141.5,426,141.5,433.5</points>
<connection>
<GID>2119</GID>
<name>ENABLE_0</name></connection>
<intersection>433.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>61,426.5,61,433.5</points>
<connection>
<GID>2118</GID>
<name>ENABLE_0</name></connection>
<intersection>426.5 16</intersection>
<intersection>433.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>14,426.5,61,426.5</points>
<connection>
<GID>2129</GID>
<name>IN_0</name></connection>
<intersection>61 15</intersection></hsegment></shape></wire>
<wire>
<ID>1456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-21.5,-35,400</points>
<connection>
<GID>2147</GID>
<name>IN_0</name></connection>
<intersection>-21.5 9</intersection>
<intersection>96.5 7</intersection>
<intersection>186.5 5</intersection>
<intersection>264.5 3</intersection>
<intersection>354.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,354.5,-31,354.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-35,264.5,-28,264.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-35,186.5,-27,186.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-35,96.5,-24,96.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-35,-21.5,-29,-21.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>-35 0</intersection>
<intersection>-34.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-34.5,-279.5,-34.5,-21.5</points>
<intersection>-279.5 15</intersection>
<intersection>-189.5 13</intersection>
<intersection>-111.5 11</intersection>
<intersection>-21.5 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-34.5,-111.5,-26,-111.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>-34.5 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-34.5,-189.5,-25,-189.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>-34.5 10</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-34.5,-279.5,-22,-279.5</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>-34.5 10</intersection>
<intersection>-34 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-34,-471,-34,-279.5</points>
<intersection>-471 17</intersection>
<intersection>-279.5 15</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-38.5,-471,-31,-471</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection>
<intersection>-34 16</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-38.5,-6416.5,-38.5,-471</points>
<intersection>-6416.5 21</intersection>
<intersection>-6326.5 83</intersection>
<intersection>-6248.5 82</intersection>
<intersection>-6158.5 81</intersection>
<intersection>-6040.5 80</intersection>
<intersection>-5950.5 79</intersection>
<intersection>-5872.5 78</intersection>
<intersection>-5782.5 77</intersection>
<intersection>-5545 76</intersection>
<intersection>-5455 75</intersection>
<intersection>-5377 74</intersection>
<intersection>-5287 73</intersection>
<intersection>-5169 72</intersection>
<intersection>-5079 65</intersection>
<intersection>-5001 64</intersection>
<intersection>-4911 63</intersection>
<intersection>-4620.5 62</intersection>
<intersection>-4530.5 61</intersection>
<intersection>-4452.5 60</intersection>
<intersection>-4362.5 59</intersection>
<intersection>-4244.5 58</intersection>
<intersection>-4154.5 57</intersection>
<intersection>-4076.5 56</intersection>
<intersection>-3986.5 53</intersection>
<intersection>-3795 52</intersection>
<intersection>-3705 51</intersection>
<intersection>-3627 50</intersection>
<intersection>-3537 49</intersection>
<intersection>-3419 48</intersection>
<intersection>-3329 47</intersection>
<intersection>-3251 46</intersection>
<intersection>-3161 45</intersection>
<intersection>-2901 44</intersection>
<intersection>-2811 43</intersection>
<intersection>-2733 42</intersection>
<intersection>-2643 41</intersection>
<intersection>-2525 40</intersection>
<intersection>-2435 39</intersection>
<intersection>-2357 38</intersection>
<intersection>-2267 37</intersection>
<intersection>-2029.5 36</intersection>
<intersection>-1939.5 35</intersection>
<intersection>-1861.5 34</intersection>
<intersection>-1771.5 33</intersection>
<intersection>-1653.5 32</intersection>
<intersection>-1635.5 31</intersection>
<intersection>-1563.5 30</intersection>
<intersection>-1485.5 29</intersection>
<intersection>-1396 28</intersection>
<intersection>-1105 27</intersection>
<intersection>-1015 26</intersection>
<intersection>-937 25</intersection>
<intersection>-847 24</intersection>
<intersection>-729 23</intersection>
<intersection>-639 22</intersection>
<intersection>-561 19</intersection>
<intersection>-471 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-38.5,-561,-28,-561</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-38.5,-6416.5,-27,-6416.5</points>
<connection>
<GID>1756</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-38.5,-639,-27,-639</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-38.5,-729,-24,-729</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-38.5,-847,-29,-847</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-38.5,-937,-26,-937</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-38.5,-1015,-25,-1015</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-38.5,-1105,-22,-1105</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-38.5,-1396,-29,-1396</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-38.5,-1485.5,-30.5,-1485.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-38.5,-1563.5,-29.5,-1563.5</points>
<connection>
<GID>842</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-38.5,-1635.5,-5,-1635.5</points>
<connection>
<GID>815</GID>
<name>IN_1</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-38.5,-1653.5,-26.5,-1653.5</points>
<connection>
<GID>816</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>-38.5,-1771.5,-31.5,-1771.5</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-38.5,-1861.5,-28.5,-1861.5</points>
<connection>
<GID>868</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-38.5,-1939.5,-27.5,-1939.5</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-38.5,-2029.5,-24.5,-2029.5</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-38.5,-2267,-34,-2267</points>
<connection>
<GID>999</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>-38.5,-2357,-31,-2357</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-38.5,-2435,-30,-2435</points>
<connection>
<GID>1051</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>-38.5,-2525,-27,-2525</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>-38.5,-2643,-32,-2643</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>-38.5,-2733,-29,-2733</points>
<connection>
<GID>1077</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>-38.5,-2811,-28,-2811</points>
<connection>
<GID>946</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>-38.5,-2901,-25,-2901</points>
<connection>
<GID>920</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-38.5,-3161,-33,-3161</points>
<connection>
<GID>1138</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>-38.5,-3251,-30,-3251</points>
<connection>
<GID>1112</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>-38.5,-3329,-29,-3329</points>
<connection>
<GID>1190</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-38.5,-3419,-26,-3419</points>
<connection>
<GID>1164</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>-38.5,-3537,-31,-3537</points>
<connection>
<GID>1242</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-38.5,-3627,-28,-3627</points>
<connection>
<GID>1216</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>-38.5,-3705,-27,-3705</points>
<connection>
<GID>1294</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>-38.5,-3795,-24,-3795</points>
<connection>
<GID>1268</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>-38.5,-3986.5,-33,-3986.5</points>
<connection>
<GID>1417</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>-38.5,-4076.5,-30,-4076.5</points>
<connection>
<GID>1391</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>-38.5,-4154.5,-29,-4154.5</points>
<connection>
<GID>1469</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>-38.5,-4244.5,-26,-4244.5</points>
<connection>
<GID>1443</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>-38.5,-4362.5,-31,-4362.5</points>
<connection>
<GID>1312</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>-38.5,-4452.5,-28,-4452.5</points>
<connection>
<GID>1495</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>-38.5,-4530.5,-27,-4530.5</points>
<connection>
<GID>1364</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>-38.5,-4620.5,-24,-4620.5</points>
<connection>
<GID>1338</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>-38.5,-4911,-35.5,-4911</points>
<connection>
<GID>1626</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>-38.5,-5001,-32.5,-5001</points>
<connection>
<GID>1600</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>-38.5,-5079,-31.5,-5079</points>
<connection>
<GID>1678</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>-38.5,-5169,-28.5,-5169</points>
<connection>
<GID>1652</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>-38.5,-5287,-33.5,-5287</points>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>-38.5,-5377,-30.5,-5377</points>
<connection>
<GID>1704</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>-38.5,-5455,-29.5,-5455</points>
<connection>
<GID>1573</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>-38.5,-5545,-26.5,-5545</points>
<connection>
<GID>1547</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>-38.5,-5782.5,-36,-5782.5</points>
<connection>
<GID>1835</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>-38.5,-5872.5,-33,-5872.5</points>
<connection>
<GID>1809</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>-38.5,-5950.5,-32,-5950.5</points>
<connection>
<GID>1887</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>80</ID>
<points>-38.5,-6040.5,-29,-6040.5</points>
<connection>
<GID>1861</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>81</ID>
<points>-38.5,-6158.5,-34,-6158.5</points>
<connection>
<GID>1730</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>82</ID>
<points>-38.5,-6248.5,-31,-6248.5</points>
<connection>
<GID>1913</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment>
<hsegment>
<ID>83</ID>
<points>-38.5,-6326.5,-30,-6326.5</points>
<connection>
<GID>1782</GID>
<name>IN_0</name></connection>
<intersection>-38.5 18</intersection></hsegment></shape></wire>
<wire>
<ID>1457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-263.5,63,423.5</points>
<connection>
<GID>2118</GID>
<name>IN_0</name></connection>
<intersection>-263.5 17</intersection>
<intersection>-173.5 15</intersection>
<intersection>-95.5 13</intersection>
<intersection>-5.5 11</intersection>
<intersection>112.5 9</intersection>
<intersection>202.5 7</intersection>
<intersection>280.5 5</intersection>
<intersection>370.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49.5,370.5,63,370.5</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>52.5,280.5,63,280.5</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>53.5,202.5,63,202.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>56.5,112.5,63,112.5</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>51.5,-5.5,63,-5.5</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>54.5,-95.5,63,-95.5</points>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>55.5,-173.5,63,-173.5</points>
<connection>
<GID>434</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>58.5,-263.5,63.5,-263.5</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection>
<intersection>63.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>63.5,-6400.5,63.5,-263.5</points>
<intersection>-6400.5 23</intersection>
<intersection>-6310.5 86</intersection>
<intersection>-6232.5 83</intersection>
<intersection>-6142.5 84</intersection>
<intersection>-6024.5 85</intersection>
<intersection>-5934.5 82</intersection>
<intersection>-5856.5 81</intersection>
<intersection>-5766.5 80</intersection>
<intersection>-5529 79</intersection>
<intersection>-5439 78</intersection>
<intersection>-5361 77</intersection>
<intersection>-5271 76</intersection>
<intersection>-5153 75</intersection>
<intersection>-5063.5 90</intersection>
<intersection>-4985 65</intersection>
<intersection>-4895 64</intersection>
<intersection>-4604.5 63</intersection>
<intersection>-4514.5 60</intersection>
<intersection>-4436.5 61</intersection>
<intersection>-4346.5 62</intersection>
<intersection>-4228.5 59</intersection>
<intersection>-4138.5 58</intersection>
<intersection>-4060.5 57</intersection>
<intersection>-3970.5 56</intersection>
<intersection>-3779 54</intersection>
<intersection>-3689 55</intersection>
<intersection>-3611 53</intersection>
<intersection>-3521 52</intersection>
<intersection>-3403 51</intersection>
<intersection>-3313 50</intersection>
<intersection>-3235 49</intersection>
<intersection>-3145 48</intersection>
<intersection>-2885 47</intersection>
<intersection>-2795 46</intersection>
<intersection>-2717 45</intersection>
<intersection>-2509 41</intersection>
<intersection>-2419 40</intersection>
<intersection>-2341 39</intersection>
<intersection>-2251 38</intersection>
<intersection>-2013.5 37</intersection>
<intersection>-1923.5 36</intersection>
<intersection>-1845.5 34</intersection>
<intersection>-1755.5 35</intersection>
<intersection>-1637.5 33</intersection>
<intersection>-1547.5 32</intersection>
<intersection>-1469.5 31</intersection>
<intersection>-1379.5 30</intersection>
<intersection>-1089 24</intersection>
<intersection>-999 26</intersection>
<intersection>-921 25</intersection>
<intersection>-831 27</intersection>
<intersection>-713 29</intersection>
<intersection>-623 28</intersection>
<intersection>-545 21</intersection>
<intersection>-455 19</intersection>
<intersection>-263.5 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>49.5,-455,63.5,-455</points>
<connection>
<GID>558</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>52.5,-545,63.5,-545</points>
<connection>
<GID>532</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>53.5,-6400.5,63.5,-6400.5</points>
<connection>
<GID>1733</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>58.5,-1089,63.5,-1089</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>54.5,-921,63.5,-921</points>
<connection>
<GID>636</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>55.5,-999,63.5,-999</points>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>51.5,-831,63.5,-831</points>
<connection>
<GID>662</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>53.5,-623,63.5,-623</points>
<connection>
<GID>610</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>56.5,-713,63.5,-713</points>
<connection>
<GID>584</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>47,-1379.5,63.5,-1379.5</points>
<connection>
<GID>767</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>50,-1469.5,63.5,-1469.5</points>
<connection>
<GID>741</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>51,-1547.5,63.5,-1547.5</points>
<connection>
<GID>819</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>54,-1637.5,63.5,-1637.5</points>
<connection>
<GID>793</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>52,-1845.5,63.5,-1845.5</points>
<connection>
<GID>845</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>49,-1755.5,63.5,-1755.5</points>
<connection>
<GID>871</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>53,-1923.5,63.5,-1923.5</points>
<connection>
<GID>714</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>56,-2013.5,63.5,-2013.5</points>
<connection>
<GID>688</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>46.5,-2251,63.5,-2251</points>
<connection>
<GID>976</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>49.5,-2341,63.5,-2341</points>
<connection>
<GID>950</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>50.5,-2419,63.5,-2419</points>
<connection>
<GID>1028</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>53.5,-2509,63.5,-2509</points>
<connection>
<GID>1002</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>37,-2629.5,46.5,-2629.5</points>
<connection>
<GID>1081</GID>
<name>OUT</name></connection>
<connection>
<GID>1080</GID>
<name>ENABLE_0</name></connection></hsegment>
<hsegment>
<ID>45</ID>
<points>51.5,-2717,63.5,-2717</points>
<connection>
<GID>1054</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>52.5,-2795,63.5,-2795</points>
<connection>
<GID>923</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>55.5,-2885,63.5,-2885</points>
<connection>
<GID>897</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>47.5,-3145,63.5,-3145</points>
<connection>
<GID>1115</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>50.5,-3235,63.5,-3235</points>
<connection>
<GID>1089</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>51.5,-3313,63.5,-3313</points>
<connection>
<GID>1167</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>54.5,-3403,63.5,-3403</points>
<connection>
<GID>1141</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>49.5,-3521,63.5,-3521</points>
<connection>
<GID>1219</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>52.5,-3611,63.5,-3611</points>
<connection>
<GID>1193</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>56.5,-3779,63.5,-3779</points>
<connection>
<GID>1245</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>53.5,-3689,63.5,-3689</points>
<connection>
<GID>1271</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>47.5,-3970.5,63.5,-3970.5</points>
<connection>
<GID>1394</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>50.5,-4060.5,63.5,-4060.5</points>
<connection>
<GID>1368</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>51.5,-4138.5,63.5,-4138.5</points>
<connection>
<GID>1446</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>54.5,-4228.5,63.5,-4228.5</points>
<connection>
<GID>1420</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>53.5,-4514.5,63.5,-4514.5</points>
<connection>
<GID>1341</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>52.5,-4436.5,63.5,-4436.5</points>
<connection>
<GID>1472</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>49.5,-4346.5,63.5,-4346.5</points>
<connection>
<GID>1498</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>56.5,-4604.5,63.5,-4604.5</points>
<connection>
<GID>1315</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>45,-4895,63.5,-4895</points>
<connection>
<GID>1603</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>48,-4985,63.5,-4985</points>
<connection>
<GID>1577</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>52,-5153,63.5,-5153</points>
<connection>
<GID>1629</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>47,-5271,63.5,-5271</points>
<connection>
<GID>1707</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>50,-5361,63.5,-5361</points>
<connection>
<GID>1681</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>51,-5439,63.5,-5439</points>
<connection>
<GID>1550</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>54,-5529,63.5,-5529</points>
<connection>
<GID>1524</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>80</ID>
<points>44.5,-5766.5,63.5,-5766.5</points>
<connection>
<GID>1812</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>81</ID>
<points>47.5,-5856.5,63.5,-5856.5</points>
<connection>
<GID>1786</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>82</ID>
<points>48.5,-5934.5,63.5,-5934.5</points>
<connection>
<GID>1864</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>83</ID>
<points>49.5,-6232.5,63.5,-6232.5</points>
<connection>
<GID>1890</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>84</ID>
<points>46.5,-6142.5,63.5,-6142.5</points>
<connection>
<GID>1916</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>85</ID>
<points>51.5,-6024.5,63.5,-6024.5</points>
<connection>
<GID>1838</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>86</ID>
<points>50.5,-6310.5,63.5,-6310.5</points>
<connection>
<GID>1759</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>42.5,-5063.5,63.5,-5063.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>63.5 18</intersection></hsegment></shape></wire>
<wire>
<ID>1458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,202.5,143.5,423</points>
<connection>
<GID>2119</GID>
<name>IN_0</name></connection>
<intersection>202.5 7</intersection>
<intersection>280.5 5</intersection>
<intersection>370.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,370.5,143.5,370.5</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>126,280.5,143.5,280.5</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>127,202.5,144,202.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>143.5 0</intersection>
<intersection>144 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>144,-545,144,202.5</points>
<intersection>-545 21</intersection>
<intersection>-455 19</intersection>
<intersection>-263.5 17</intersection>
<intersection>-173.5 15</intersection>
<intersection>-95.5 13</intersection>
<intersection>-5.5 11</intersection>
<intersection>112.5 9</intersection>
<intersection>202.5 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>130,112.5,144,112.5</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>125,-5.5,144,-5.5</points>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>128,-95.5,144,-95.5</points>
<connection>
<GID>359</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>129,-173.5,144,-173.5</points>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>132,-263.5,144,-263.5</points>
<connection>
<GID>411</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>123,-455,144,-455</points>
<connection>
<GID>561</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>126,-545,144.5,-545</points>
<connection>
<GID>535</GID>
<name>OUT_0</name></connection>
<intersection>144 8</intersection>
<intersection>144.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>144.5,-6400.5,144.5,-545</points>
<intersection>-6400.5 23</intersection>
<intersection>-6310.5 79</intersection>
<intersection>-6232.5 78</intersection>
<intersection>-6142.5 77</intersection>
<intersection>-6024.5 76</intersection>
<intersection>-5934.5 75</intersection>
<intersection>-5856.5 74</intersection>
<intersection>-5766.5 73</intersection>
<intersection>-5529 72</intersection>
<intersection>-5439 71</intersection>
<intersection>-5361 70</intersection>
<intersection>-5271 69</intersection>
<intersection>-5153 68</intersection>
<intersection>-5063 64</intersection>
<intersection>-4985 63</intersection>
<intersection>-4895 62</intersection>
<intersection>-4604.5 61</intersection>
<intersection>-4514.5 60</intersection>
<intersection>-4436.5 59</intersection>
<intersection>-4346.5 58</intersection>
<intersection>-4228.5 54</intersection>
<intersection>-4138.5 55</intersection>
<intersection>-4060.5 56</intersection>
<intersection>-3970.5 57</intersection>
<intersection>-3779 53</intersection>
<intersection>-3689 52</intersection>
<intersection>-3611 51</intersection>
<intersection>-3521 50</intersection>
<intersection>-3403 49</intersection>
<intersection>-3313 46</intersection>
<intersection>-3235 47</intersection>
<intersection>-3145 48</intersection>
<intersection>-2885 45</intersection>
<intersection>-2795 44</intersection>
<intersection>-2717 43</intersection>
<intersection>-2627 42</intersection>
<intersection>-2509 41</intersection>
<intersection>-2419 40</intersection>
<intersection>-2341 39</intersection>
<intersection>-2251 38</intersection>
<intersection>-2013.5 37</intersection>
<intersection>-1923.5 36</intersection>
<intersection>-1845.5 35</intersection>
<intersection>-1755.5 34</intersection>
<intersection>-1637.5 33</intersection>
<intersection>-1547.5 32</intersection>
<intersection>-1469.5 31</intersection>
<intersection>-1379.5 30</intersection>
<intersection>-1089 24</intersection>
<intersection>-999 27</intersection>
<intersection>-921 26</intersection>
<intersection>-831 25</intersection>
<intersection>-713 28</intersection>
<intersection>-623 29</intersection>
<intersection>-545 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>127,-6400.5,144.5,-6400.5</points>
<connection>
<GID>1736</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>132,-1089,144.5,-1089</points>
<connection>
<GID>482</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>125,-831,144.5,-831</points>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>129,-921,144.5,-921</points>
<connection>
<GID>639</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>129,-999,144.5,-999</points>
<connection>
<GID>508</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>130,-713,144.5,-713</points>
<connection>
<GID>587</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>127,-623,144.5,-623</points>
<connection>
<GID>613</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>120.5,-1379.5,144.5,-1379.5</points>
<connection>
<GID>770</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>123.5,-1469.5,144.5,-1469.5</points>
<connection>
<GID>744</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>124.5,-1547.5,144.5,-1547.5</points>
<connection>
<GID>822</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>127.5,-1637.5,144.5,-1637.5</points>
<connection>
<GID>796</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>122.5,-1755.5,144.5,-1755.5</points>
<connection>
<GID>874</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>125.5,-1845.5,144.5,-1845.5</points>
<connection>
<GID>848</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>126.5,-1923.5,144.5,-1923.5</points>
<connection>
<GID>717</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>129.5,-2013.5,144.5,-2013.5</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>120,-2251,144.5,-2251</points>
<connection>
<GID>979</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>123,-2341,144.5,-2341</points>
<connection>
<GID>953</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>124,-2419,144.5,-2419</points>
<connection>
<GID>1031</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>127,-2509,144.5,-2509</points>
<connection>
<GID>1005</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>122,-2627,144.5,-2627</points>
<connection>
<GID>1083</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>125,-2717,144.5,-2717</points>
<connection>
<GID>1057</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>126,-2795,144.5,-2795</points>
<connection>
<GID>926</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>129,-2885,144.5,-2885</points>
<connection>
<GID>900</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>125,-3313,144.5,-3313</points>
<connection>
<GID>1170</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>124,-3235,144.5,-3235</points>
<connection>
<GID>1092</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>121,-3145,144.5,-3145</points>
<connection>
<GID>1118</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>128,-3403,144.5,-3403</points>
<connection>
<GID>1144</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>123,-3521,144.5,-3521</points>
<connection>
<GID>1222</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>126,-3611,144.5,-3611</points>
<connection>
<GID>1196</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>127,-3689,144.5,-3689</points>
<connection>
<GID>1274</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>130,-3779,144.5,-3779</points>
<connection>
<GID>1248</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>128,-4228.5,144.5,-4228.5</points>
<connection>
<GID>1423</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>125,-4138.5,144.5,-4138.5</points>
<connection>
<GID>1449</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>124,-4060.5,144.5,-4060.5</points>
<connection>
<GID>1371</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>121,-3970.5,144.5,-3970.5</points>
<connection>
<GID>1397</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>123,-4346.5,144.5,-4346.5</points>
<connection>
<GID>1501</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>126,-4436.5,144.5,-4436.5</points>
<connection>
<GID>1475</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>127,-4514.5,144.5,-4514.5</points>
<connection>
<GID>1344</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>130,-4604.5,144.5,-4604.5</points>
<connection>
<GID>1318</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>118.5,-4895,144.5,-4895</points>
<connection>
<GID>1606</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>121.5,-4985,144.5,-4985</points>
<connection>
<GID>1580</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>122.5,-5063,144.5,-5063</points>
<connection>
<GID>1658</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>125.5,-5153,144.5,-5153</points>
<connection>
<GID>1632</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>120.5,-5271,144.5,-5271</points>
<connection>
<GID>1710</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>123.5,-5361,144.5,-5361</points>
<connection>
<GID>1684</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>124.5,-5439,144.5,-5439</points>
<connection>
<GID>1553</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>127.5,-5529,144.5,-5529</points>
<connection>
<GID>1527</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>118,-5766.5,144.5,-5766.5</points>
<connection>
<GID>1815</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>121,-5856.5,144.5,-5856.5</points>
<connection>
<GID>1789</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>122,-5934.5,144.5,-5934.5</points>
<connection>
<GID>1867</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>125,-6024.5,144.5,-6024.5</points>
<connection>
<GID>1841</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>120,-6142.5,144.5,-6142.5</points>
<connection>
<GID>1919</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>123,-6232.5,144.5,-6232.5</points>
<connection>
<GID>1893</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>124,-6310.5,144.5,-6310.5</points>
<connection>
<GID>1762</GID>
<name>OUT_0</name></connection>
<intersection>144.5 22</intersection></hsegment></shape></wire>
<wire>
<ID>1459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-7.5,220,425</points>
<connection>
<GID>2132</GID>
<name>IN_0</name></connection>
<intersection>-7.5 11</intersection>
<intersection>110.5 9</intersection>
<intersection>200.5 7</intersection>
<intersection>278.5 5</intersection>
<intersection>368.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>207.5,368.5,220,368.5</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>210.5,278.5,220,278.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>211.5,200.5,220,200.5</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>214.5,110.5,220,110.5</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>209.5,-7.5,220,-7.5</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<intersection>219.5 12</intersection>
<intersection>220 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>219.5,-265.5,219.5,-7.5</points>
<intersection>-265.5 17</intersection>
<intersection>-175.5 15</intersection>
<intersection>-97.5 13</intersection>
<intersection>-7.5 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>212.5,-97.5,219.5,-97.5</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<intersection>219.5 12</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>213.5,-175.5,219.5,-175.5</points>
<connection>
<GID>440</GID>
<name>OUT_0</name></connection>
<intersection>219.5 12</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>216.5,-265.5,220,-265.5</points>
<connection>
<GID>414</GID>
<name>OUT_0</name></connection>
<intersection>219.5 12</intersection>
<intersection>220 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>220,-457,220,-265.5</points>
<intersection>-457 19</intersection>
<intersection>-265.5 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>207.5,-457,220.5,-457</points>
<connection>
<GID>564</GID>
<name>OUT_0</name></connection>
<intersection>220 18</intersection>
<intersection>220.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>220.5,-547,220.5,-457</points>
<intersection>-547 21</intersection>
<intersection>-457 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>210.5,-547,221,-547</points>
<connection>
<GID>538</GID>
<name>OUT_0</name></connection>
<intersection>220.5 20</intersection>
<intersection>221 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>221,-6402.5,221,-547</points>
<intersection>-6402.5 23</intersection>
<intersection>-6312.5 77</intersection>
<intersection>-6234.5 74</intersection>
<intersection>-6144.5 75</intersection>
<intersection>-6026.5 76</intersection>
<intersection>-5936.5 73</intersection>
<intersection>-5858.5 72</intersection>
<intersection>-5768.5 71</intersection>
<intersection>-5531 69</intersection>
<intersection>-5441 70</intersection>
<intersection>-5363 68</intersection>
<intersection>-5273 67</intersection>
<intersection>-5155 66</intersection>
<intersection>-5065 62</intersection>
<intersection>-4987 61</intersection>
<intersection>-4897 60</intersection>
<intersection>-4606.5 59</intersection>
<intersection>-4516.5 58</intersection>
<intersection>-4438.5 57</intersection>
<intersection>-4348.5 56</intersection>
<intersection>-4230.5 55</intersection>
<intersection>-4140.5 54</intersection>
<intersection>-4062.5 53</intersection>
<intersection>-3972.5 52</intersection>
<intersection>-3781 51</intersection>
<intersection>-3691 50</intersection>
<intersection>-3613 48</intersection>
<intersection>-3523 47</intersection>
<intersection>-3405 49</intersection>
<intersection>-3315 46</intersection>
<intersection>-3237 45</intersection>
<intersection>-3147 44</intersection>
<intersection>-2887 43</intersection>
<intersection>-2797 42</intersection>
<intersection>-2719 41</intersection>
<intersection>-2629 40</intersection>
<intersection>-2511 39</intersection>
<intersection>-2421 38</intersection>
<intersection>-2343 37</intersection>
<intersection>-2253 36</intersection>
<intersection>-2015.5 35</intersection>
<intersection>-1925.5 34</intersection>
<intersection>-1757.5 33</intersection>
<intersection>-1639.5 32</intersection>
<intersection>-1549.5 31</intersection>
<intersection>-1471.5 30</intersection>
<intersection>-1091 24</intersection>
<intersection>-1001 27</intersection>
<intersection>-923 26</intersection>
<intersection>-833 25</intersection>
<intersection>-715 29</intersection>
<intersection>-625 28</intersection>
<intersection>-547 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>211.5,-6402.5,221,-6402.5</points>
<connection>
<GID>1739</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>216.5,-1091,221,-1091</points>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>209.5,-833,221,-833</points>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>212.5,-923,221,-923</points>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>213.5,-1001,221,-1001</points>
<connection>
<GID>511</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>211.5,-625,221,-625</points>
<connection>
<GID>616</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>214.5,-715,221,-715</points>
<connection>
<GID>590</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>208,-1471.5,221,-1471.5</points>
<connection>
<GID>747</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>209,-1549.5,221,-1549.5</points>
<connection>
<GID>825</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>212,-1639.5,221,-1639.5</points>
<connection>
<GID>799</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>207,-1757.5,221,-1757.5</points>
<connection>
<GID>877</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>211,-1925.5,221,-1925.5</points>
<connection>
<GID>720</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>214,-2015.5,221,-2015.5</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>204.5,-2253,221,-2253</points>
<connection>
<GID>982</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>207.5,-2343,221,-2343</points>
<connection>
<GID>956</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>208.5,-2421,221,-2421</points>
<connection>
<GID>1034</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>211.5,-2511,221,-2511</points>
<connection>
<GID>1008</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>206.5,-2629,221,-2629</points>
<connection>
<GID>1086</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>209.5,-2719,221,-2719</points>
<connection>
<GID>1060</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>210.5,-2797,221,-2797</points>
<connection>
<GID>929</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>213.5,-2887,221,-2887</points>
<connection>
<GID>903</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>205.5,-3147,221,-3147</points>
<connection>
<GID>1121</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>208.5,-3237,221,-3237</points>
<connection>
<GID>1095</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>209.5,-3315,221,-3315</points>
<connection>
<GID>1173</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>207.5,-3523,221,-3523</points>
<connection>
<GID>1225</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>210.5,-3613,221,-3613</points>
<connection>
<GID>1199</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>212.5,-3405,221,-3405</points>
<connection>
<GID>1147</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>211.5,-3691,221,-3691</points>
<connection>
<GID>1277</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>214.5,-3781,221,-3781</points>
<connection>
<GID>1251</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>205.5,-3972.5,221,-3972.5</points>
<connection>
<GID>1400</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>208.5,-4062.5,221,-4062.5</points>
<connection>
<GID>1374</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>209.5,-4140.5,221,-4140.5</points>
<connection>
<GID>1452</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>212.5,-4230.5,221,-4230.5</points>
<connection>
<GID>1426</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>207.5,-4348.5,221,-4348.5</points>
<connection>
<GID>1504</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>210.5,-4438.5,221,-4438.5</points>
<connection>
<GID>1478</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>211.5,-4516.5,221,-4516.5</points>
<connection>
<GID>1347</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>214.5,-4606.5,221,-4606.5</points>
<connection>
<GID>1321</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>203,-4897,221,-4897</points>
<connection>
<GID>1609</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>206,-4987,221,-4987</points>
<connection>
<GID>1583</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>207,-5065,221,-5065</points>
<connection>
<GID>1661</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>210,-5155,221,-5155</points>
<connection>
<GID>1635</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>205,-5273,221,-5273</points>
<connection>
<GID>1713</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>208,-5363,221,-5363</points>
<connection>
<GID>1687</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>212,-5531,221,-5531</points>
<connection>
<GID>1530</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>209,-5441,221,-5441</points>
<connection>
<GID>1556</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>202.5,-5768.5,221,-5768.5</points>
<connection>
<GID>1818</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>205.5,-5858.5,221,-5858.5</points>
<connection>
<GID>1792</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>206.5,-5936.5,221,-5936.5</points>
<connection>
<GID>1870</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>207.5,-6234.5,221,-6234.5</points>
<connection>
<GID>1896</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>204.5,-6144.5,221,-6144.5</points>
<connection>
<GID>1922</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>209.5,-6026.5,221,-6026.5</points>
<connection>
<GID>1844</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>208.5,-6312.5,221,-6312.5</points>
<connection>
<GID>1765</GID>
<name>OUT_0</name></connection>
<intersection>221 22</intersection></hsegment></shape></wire>
<wire>
<ID>1460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-7.5,298.5,423.5</points>
<intersection>-7.5 12</intersection>
<intersection>110.5 9</intersection>
<intersection>200.5 7</intersection>
<intersection>278.5 5</intersection>
<intersection>368.5 3</intersection>
<intersection>423.5 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>281,368.5,298.5,368.5</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>284,278.5,298.5,278.5</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>285,200.5,298.5,200.5</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>288,110.5,298.5,110.5</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>288,423.5,298.5,423.5</points>
<connection>
<GID>2134</GID>
<name>IN_0</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>283,-7.5,299,-7.5</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<intersection>298.5 0</intersection>
<intersection>299 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>299,-265.5,299,-7.5</points>
<intersection>-265.5 18</intersection>
<intersection>-175.5 16</intersection>
<intersection>-97.5 14</intersection>
<intersection>-7.5 12</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>286,-97.5,299,-97.5</points>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection>
<intersection>299 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>287,-175.5,299,-175.5</points>
<connection>
<GID>443</GID>
<name>OUT_0</name></connection>
<intersection>299 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>290,-265.5,299,-265.5</points>
<connection>
<GID>417</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection>
<intersection>299 13</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>298.5,-6402.5,298.5,-265.5</points>
<intersection>-6402.5 24</intersection>
<intersection>-6312.5 79</intersection>
<intersection>-6234.5 78</intersection>
<intersection>-6144.5 76</intersection>
<intersection>-6026.5 77</intersection>
<intersection>-5936.5 75</intersection>
<intersection>-5858.5 74</intersection>
<intersection>-5768.5 73</intersection>
<intersection>-5531 72</intersection>
<intersection>-5441 71</intersection>
<intersection>-5363 70</intersection>
<intersection>-5273 69</intersection>
<intersection>-5155 68</intersection>
<intersection>-5065 64</intersection>
<intersection>-4987 63</intersection>
<intersection>-4897 62</intersection>
<intersection>-4516.5 61</intersection>
<intersection>-4438.5 60</intersection>
<intersection>-4348.5 59</intersection>
<intersection>-4230.5 58</intersection>
<intersection>-4140.5 57</intersection>
<intersection>-4062.5 56</intersection>
<intersection>-3972.5 55</intersection>
<intersection>-3781 54</intersection>
<intersection>-3691 53</intersection>
<intersection>-3613 52</intersection>
<intersection>-3523 51</intersection>
<intersection>-3405 50</intersection>
<intersection>-3315 47</intersection>
<intersection>-3237 48</intersection>
<intersection>-3147 49</intersection>
<intersection>-2887 46</intersection>
<intersection>-2797 45</intersection>
<intersection>-2719 44</intersection>
<intersection>-2629 43</intersection>
<intersection>-2511 42</intersection>
<intersection>-2421 39</intersection>
<intersection>-2343 40</intersection>
<intersection>-2253 41</intersection>
<intersection>-2015.5 38</intersection>
<intersection>-1925.5 37</intersection>
<intersection>-1847.5 36</intersection>
<intersection>-1757.5 35</intersection>
<intersection>-1639.5 31</intersection>
<intersection>-1549.5 32</intersection>
<intersection>-1471.5 33</intersection>
<intersection>-1381.5 34</intersection>
<intersection>-1091 25</intersection>
<intersection>-1001 28</intersection>
<intersection>-923 27</intersection>
<intersection>-833 26</intersection>
<intersection>-715 29</intersection>
<intersection>-625 30</intersection>
<intersection>-547 22</intersection>
<intersection>-457 20</intersection>
<intersection>-265.5 18</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>281,-457,298.5,-457</points>
<connection>
<GID>567</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>284,-547,298.5,-547</points>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>285,-6402.5,298.5,-6402.5</points>
<connection>
<GID>1742</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>290,-1091,298.5,-1091</points>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>283,-833,298.5,-833</points>
<connection>
<GID>462</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>286,-923,298.5,-923</points>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>287,-1001,298.5,-1001</points>
<connection>
<GID>514</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>288,-715,298.5,-715</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>285,-625,298.5,-625</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>285.5,-1639.5,298.5,-1639.5</points>
<connection>
<GID>802</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>282.5,-1549.5,298.5,-1549.5</points>
<connection>
<GID>828</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>281.5,-1471.5,298.5,-1471.5</points>
<connection>
<GID>750</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>278.5,-1381.5,298.5,-1381.5</points>
<connection>
<GID>776</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>280.5,-1757.5,298.5,-1757.5</points>
<connection>
<GID>671</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>283.5,-1847.5,298.5,-1847.5</points>
<connection>
<GID>854</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>284.5,-1925.5,298.5,-1925.5</points>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>287.5,-2015.5,298.5,-2015.5</points>
<connection>
<GID>697</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>282,-2421,298.5,-2421</points>
<connection>
<GID>1037</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>281,-2343,298.5,-2343</points>
<connection>
<GID>959</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>278,-2253,298.5,-2253</points>
<connection>
<GID>985</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>285,-2511,298.5,-2511</points>
<connection>
<GID>1011</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>280,-2629,298.5,-2629</points>
<connection>
<GID>880</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>283,-2719,298.5,-2719</points>
<connection>
<GID>1063</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>284,-2797,298.5,-2797</points>
<connection>
<GID>932</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>287,-2887,298.5,-2887</points>
<connection>
<GID>906</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>283,-3315,298.5,-3315</points>
<connection>
<GID>1176</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>282,-3237,298.5,-3237</points>
<connection>
<GID>1098</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>279,-3147,298.5,-3147</points>
<connection>
<GID>1124</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>286,-3405,298.5,-3405</points>
<connection>
<GID>1150</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>281,-3523,298.5,-3523</points>
<connection>
<GID>1228</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>284,-3613,298.5,-3613</points>
<connection>
<GID>1202</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>285,-3691,298.5,-3691</points>
<connection>
<GID>1280</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>288,-3781,298.5,-3781</points>
<connection>
<GID>1254</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>279,-3972.5,298.5,-3972.5</points>
<connection>
<GID>1403</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>282,-4062.5,298.5,-4062.5</points>
<connection>
<GID>1377</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>283,-4140.5,298.5,-4140.5</points>
<connection>
<GID>1455</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>286,-4230.5,298.5,-4230.5</points>
<connection>
<GID>1429</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>281,-4348.5,298.5,-4348.5</points>
<connection>
<GID>1298</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>284,-4438.5,298.5,-4438.5</points>
<connection>
<GID>1481</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>285,-4516.5,298.5,-4516.5</points>
<connection>
<GID>1350</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>276.5,-4897,298.5,-4897</points>
<connection>
<GID>1612</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>279.5,-4987,298.5,-4987</points>
<connection>
<GID>1586</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>280.5,-5065,298.5,-5065</points>
<connection>
<GID>1664</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>283.5,-5155,298.5,-5155</points>
<connection>
<GID>1638</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>278.5,-5273,298.5,-5273</points>
<connection>
<GID>1507</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>281.5,-5363,298.5,-5363</points>
<connection>
<GID>1690</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>282.5,-5441,298.5,-5441</points>
<connection>
<GID>1559</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>285.5,-5531,298.5,-5531</points>
<connection>
<GID>1533</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>276,-5768.5,298.5,-5768.5</points>
<connection>
<GID>1821</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>279,-5858.5,298.5,-5858.5</points>
<connection>
<GID>1795</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>280,-5936.5,298.5,-5936.5</points>
<connection>
<GID>1873</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>278,-6144.5,298.5,-6144.5</points>
<connection>
<GID>1716</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>283,-6026.5,298.5,-6026.5</points>
<connection>
<GID>1847</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>281,-6234.5,298.5,-6234.5</points>
<connection>
<GID>1899</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>282,-6312.5,298.5,-6312.5</points>
<connection>
<GID>1768</GID>
<name>OUT_0</name></connection>
<intersection>298.5 19</intersection></hsegment></shape></wire>
<wire>
<ID>1461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-6404,396.5,425.5</points>
<intersection>-6404 24</intersection>
<intersection>-6314 80</intersection>
<intersection>-6236 79</intersection>
<intersection>-6146 78</intersection>
<intersection>-6028 77</intersection>
<intersection>-5938 76</intersection>
<intersection>-5860 75</intersection>
<intersection>-5770 74</intersection>
<intersection>-5532.5 73</intersection>
<intersection>-5442.5 72</intersection>
<intersection>-5364.5 71</intersection>
<intersection>-5274.5 70</intersection>
<intersection>-5156.5 69</intersection>
<intersection>-5066.5 65</intersection>
<intersection>-4988.5 64</intersection>
<intersection>-4898.5 63</intersection>
<intersection>-4608 62</intersection>
<intersection>-4518 61</intersection>
<intersection>-4440 60</intersection>
<intersection>-4350 59</intersection>
<intersection>-4232 58</intersection>
<intersection>-4142 57</intersection>
<intersection>-4064 56</intersection>
<intersection>-3974 55</intersection>
<intersection>-3782.5 54</intersection>
<intersection>-3692.5 53</intersection>
<intersection>-3614.5 52</intersection>
<intersection>-3524.5 51</intersection>
<intersection>-3406.5 50</intersection>
<intersection>-3316.5 49</intersection>
<intersection>-3238.5 48</intersection>
<intersection>-3148.5 47</intersection>
<intersection>-2888.5 46</intersection>
<intersection>-2798.5 45</intersection>
<intersection>-2720.5 44</intersection>
<intersection>-2630.5 43</intersection>
<intersection>-2512.5 42</intersection>
<intersection>-2422.5 41</intersection>
<intersection>-2344.5 39</intersection>
<intersection>-2254.5 40</intersection>
<intersection>-2017 38</intersection>
<intersection>-1927 37</intersection>
<intersection>-1849 35</intersection>
<intersection>-1759 36</intersection>
<intersection>-1641 34</intersection>
<intersection>-1551 33</intersection>
<intersection>-1473 32</intersection>
<intersection>-1383 31</intersection>
<intersection>-1092.5 25</intersection>
<intersection>-1002.5 28</intersection>
<intersection>-924.5 27</intersection>
<intersection>-834.5 26</intersection>
<intersection>-716.5 30</intersection>
<intersection>-626.5 29</intersection>
<intersection>-548.5 22</intersection>
<intersection>-458.5 20</intersection>
<intersection>-267 18</intersection>
<intersection>-177 16</intersection>
<intersection>-99 14</intersection>
<intersection>-9 12</intersection>
<intersection>108.5 10</intersection>
<intersection>199 7</intersection>
<intersection>277 5</intersection>
<intersection>367 3</intersection>
<intersection>425.5 9</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>372.5,367,396.5,367</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>375.5,277,396.5,277</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>376.5,199,396.5,199</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>379.5,425.5,396.5,425.5</points>
<connection>
<GID>2136</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>386,108.5,396.5,108.5</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>374.5,-9,396.5,-9</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>377.5,-99,396.5,-99</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>378.5,-177,396.5,-177</points>
<connection>
<GID>446</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>381.5,-267,396.5,-267</points>
<connection>
<GID>420</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>372.5,-458.5,396.5,-458.5</points>
<connection>
<GID>570</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>375.5,-548.5,396.5,-548.5</points>
<connection>
<GID>544</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>376.5,-6404,396.5,-6404</points>
<connection>
<GID>1745</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>381.5,-1092.5,396.5,-1092.5</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>374.5,-834.5,396.5,-834.5</points>
<connection>
<GID>465</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>377.5,-924.5,396.5,-924.5</points>
<connection>
<GID>648</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>378.5,-1002.5,396.5,-1002.5</points>
<connection>
<GID>517</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>376.5,-626.5,396.5,-626.5</points>
<connection>
<GID>622</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>379.5,-716.5,396.5,-716.5</points>
<connection>
<GID>596</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>370,-1383,396.5,-1383</points>
<connection>
<GID>779</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>373,-1473,396.5,-1473</points>
<connection>
<GID>753</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>374,-1551,396.5,-1551</points>
<connection>
<GID>831</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>377,-1641,396.5,-1641</points>
<connection>
<GID>805</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>375,-1849,396.5,-1849</points>
<connection>
<GID>857</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>372,-1759,396.5,-1759</points>
<connection>
<GID>674</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>376,-1927,396.5,-1927</points>
<connection>
<GID>726</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>379,-2017,396.5,-2017</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>372.5,-2344.5,396.5,-2344.5</points>
<connection>
<GID>962</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>369.5,-2254.5,396.5,-2254.5</points>
<connection>
<GID>988</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>373.5,-2422.5,396.5,-2422.5</points>
<connection>
<GID>1040</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>376.5,-2512.5,396.5,-2512.5</points>
<connection>
<GID>1014</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>371.5,-2630.5,396.5,-2630.5</points>
<connection>
<GID>883</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>374.5,-2720.5,396.5,-2720.5</points>
<connection>
<GID>1066</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>375.5,-2798.5,396.5,-2798.5</points>
<connection>
<GID>935</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>378.5,-2888.5,396.5,-2888.5</points>
<connection>
<GID>909</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>370.5,-3148.5,396.5,-3148.5</points>
<connection>
<GID>1127</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>373.5,-3238.5,396.5,-3238.5</points>
<connection>
<GID>1101</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>374.5,-3316.5,396.5,-3316.5</points>
<connection>
<GID>1179</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>377.5,-3406.5,396.5,-3406.5</points>
<connection>
<GID>1153</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>372.5,-3524.5,396.5,-3524.5</points>
<connection>
<GID>1231</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>375.5,-3614.5,396.5,-3614.5</points>
<connection>
<GID>1205</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>376.5,-3692.5,396.5,-3692.5</points>
<connection>
<GID>1283</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>379.5,-3782.5,396.5,-3782.5</points>
<connection>
<GID>1257</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>370.5,-3974,396.5,-3974</points>
<connection>
<GID>1406</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>373.5,-4064,396.5,-4064</points>
<connection>
<GID>1380</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>374.5,-4142,396.5,-4142</points>
<connection>
<GID>1458</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>377.5,-4232,396.5,-4232</points>
<connection>
<GID>1432</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>372.5,-4350,396.5,-4350</points>
<connection>
<GID>1301</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>375.5,-4440,396.5,-4440</points>
<connection>
<GID>1484</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>376.5,-4518,396.5,-4518</points>
<connection>
<GID>1353</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>379.5,-4608,396.5,-4608</points>
<connection>
<GID>1327</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>368,-4898.5,396.5,-4898.5</points>
<connection>
<GID>1615</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>371,-4988.5,396.5,-4988.5</points>
<connection>
<GID>1589</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>372,-5066.5,396.5,-5066.5</points>
<connection>
<GID>1667</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>375,-5156.5,396.5,-5156.5</points>
<connection>
<GID>1641</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>370,-5274.5,396.5,-5274.5</points>
<connection>
<GID>1510</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>373,-5364.5,396.5,-5364.5</points>
<connection>
<GID>1693</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>374,-5442.5,396.5,-5442.5</points>
<connection>
<GID>1562</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>377,-5532.5,396.5,-5532.5</points>
<connection>
<GID>1536</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>367.5,-5770,396.5,-5770</points>
<connection>
<GID>1824</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>370.5,-5860,396.5,-5860</points>
<connection>
<GID>1798</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>371.5,-5938,396.5,-5938</points>
<connection>
<GID>1876</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>374.5,-6028,396.5,-6028</points>
<connection>
<GID>1850</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>369.5,-6146,396.5,-6146</points>
<connection>
<GID>1719</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>372.5,-6236,396.5,-6236</points>
<connection>
<GID>1902</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>80</ID>
<points>373.5,-6314,396.5,-6314</points>
<connection>
<GID>1771</GID>
<name>OUT_0</name></connection>
<intersection>396.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-99,458.5,424.5</points>
<connection>
<GID>2138</GID>
<name>IN_0</name></connection>
<intersection>-99 13</intersection>
<intersection>-9 11</intersection>
<intersection>109 9</intersection>
<intersection>199 7</intersection>
<intersection>277 5</intersection>
<intersection>367 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>446,367,458.5,367</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>449,277,458.5,277</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>450,199,458.5,199</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>453,109,458.5,109</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>448,-9,458.5,-9</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>451,-99,459,-99</points>
<connection>
<GID>371</GID>
<name>OUT_0</name></connection>
<intersection>458.5 0</intersection>
<intersection>459 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>459,-458.5,459,-99</points>
<intersection>-458.5 19</intersection>
<intersection>-267 17</intersection>
<intersection>-177 15</intersection>
<intersection>-99 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>452,-177,459,-177</points>
<connection>
<GID>449</GID>
<name>OUT_0</name></connection>
<intersection>459 14</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>455,-267,459,-267</points>
<connection>
<GID>423</GID>
<name>OUT_0</name></connection>
<intersection>459 14</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>446,-458.5,459.5,-458.5</points>
<connection>
<GID>573</GID>
<name>OUT_0</name></connection>
<intersection>459 14</intersection>
<intersection>459.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>459.5,-6404,459.5,-458.5</points>
<intersection>-6404 23</intersection>
<intersection>-6314 75</intersection>
<intersection>-6236 74</intersection>
<intersection>-6146 73</intersection>
<intersection>-6028 72</intersection>
<intersection>-5938 71</intersection>
<intersection>-5860 70</intersection>
<intersection>-5770 69</intersection>
<intersection>-5532.5 68</intersection>
<intersection>-5442.5 67</intersection>
<intersection>-5364.5 65</intersection>
<intersection>-5274.5 64</intersection>
<intersection>-5156.5 66</intersection>
<intersection>-5066.5 63</intersection>
<intersection>-4988.5 62</intersection>
<intersection>-4898.5 61</intersection>
<intersection>-4608 60</intersection>
<intersection>-4518 57</intersection>
<intersection>-4440 58</intersection>
<intersection>-4350 59</intersection>
<intersection>-4232 56</intersection>
<intersection>-4142 54</intersection>
<intersection>-4064 55</intersection>
<intersection>-3974 53</intersection>
<intersection>-3782.5 52</intersection>
<intersection>-3692.5 51</intersection>
<intersection>-3614.5 50</intersection>
<intersection>-3524.5 49</intersection>
<intersection>-3406.5 48</intersection>
<intersection>-3316.5 47</intersection>
<intersection>-3238.5 46</intersection>
<intersection>-3148.5 45</intersection>
<intersection>-2888.5 44</intersection>
<intersection>-2798.5 43</intersection>
<intersection>-2720.5 42</intersection>
<intersection>-2512.5 41</intersection>
<intersection>-2422.5 40</intersection>
<intersection>-2344.5 38</intersection>
<intersection>-2254.5 39</intersection>
<intersection>-2017 37</intersection>
<intersection>-1927 36</intersection>
<intersection>-1849 35</intersection>
<intersection>-1759 34</intersection>
<intersection>-1641 33</intersection>
<intersection>-1551 32</intersection>
<intersection>-1473 31</intersection>
<intersection>-1383 30</intersection>
<intersection>-1092.5 24</intersection>
<intersection>-1002.5 25</intersection>
<intersection>-924.5 26</intersection>
<intersection>-834.5 27</intersection>
<intersection>-716.5 29</intersection>
<intersection>-626.5 28</intersection>
<intersection>-548.5 21</intersection>
<intersection>-458.5 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>449,-548.5,459.5,-548.5</points>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>450,-6404,459.5,-6404</points>
<connection>
<GID>1748</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>455,-1092.5,459.5,-1092.5</points>
<connection>
<GID>494</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>452,-1002.5,459.5,-1002.5</points>
<connection>
<GID>520</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>451,-924.5,459.5,-924.5</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>448,-834.5,459.5,-834.5</points>
<connection>
<GID>468</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>450,-626.5,459.5,-626.5</points>
<connection>
<GID>625</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>453,-716.5,459.5,-716.5</points>
<connection>
<GID>599</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>443.5,-1383,459.5,-1383</points>
<connection>
<GID>782</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>446.5,-1473,459.5,-1473</points>
<connection>
<GID>756</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>447.5,-1551,459.5,-1551</points>
<connection>
<GID>834</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>450.5,-1641,459.5,-1641</points>
<connection>
<GID>808</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>445.5,-1759,459.5,-1759</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>448.5,-1849,459.5,-1849</points>
<connection>
<GID>860</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>449.5,-1927,459.5,-1927</points>
<connection>
<GID>729</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>452.5,-2017,459.5,-2017</points>
<connection>
<GID>703</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>446,-2344.5,459.5,-2344.5</points>
<connection>
<GID>965</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>443,-2254.5,459.5,-2254.5</points>
<connection>
<GID>991</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>447,-2422.5,459.5,-2422.5</points>
<connection>
<GID>1043</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>450,-2512.5,459.5,-2512.5</points>
<connection>
<GID>1017</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>448,-2720.5,459.5,-2720.5</points>
<connection>
<GID>1069</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>449,-2798.5,459.5,-2798.5</points>
<connection>
<GID>938</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>452,-2888.5,459.5,-2888.5</points>
<connection>
<GID>912</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>444,-3148.5,459.5,-3148.5</points>
<connection>
<GID>1130</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>447,-3238.5,459.5,-3238.5</points>
<connection>
<GID>1104</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>448,-3316.5,459.5,-3316.5</points>
<connection>
<GID>1182</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>451,-3406.5,459.5,-3406.5</points>
<connection>
<GID>1156</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>446,-3524.5,459.5,-3524.5</points>
<connection>
<GID>1234</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>449,-3614.5,459.5,-3614.5</points>
<connection>
<GID>1208</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>450,-3692.5,459.5,-3692.5</points>
<connection>
<GID>1286</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>453,-3782.5,459.5,-3782.5</points>
<connection>
<GID>1260</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>444,-3974,459.5,-3974</points>
<connection>
<GID>1409</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>448,-4142,459.5,-4142</points>
<connection>
<GID>1461</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>447,-4064,459.5,-4064</points>
<connection>
<GID>1383</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>451,-4232,459.5,-4232</points>
<connection>
<GID>1435</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>450,-4518,459.5,-4518</points>
<connection>
<GID>1356</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>449,-4440,459.5,-4440</points>
<connection>
<GID>1487</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>446,-4350,459.5,-4350</points>
<connection>
<GID>1304</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>453,-4608,459.5,-4608</points>
<connection>
<GID>1330</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>441.5,-4898.5,459.5,-4898.5</points>
<connection>
<GID>1618</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>444.5,-4988.5,459.5,-4988.5</points>
<connection>
<GID>1592</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>445.5,-5066.5,459.5,-5066.5</points>
<connection>
<GID>1670</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>443.5,-5274.5,459.5,-5274.5</points>
<connection>
<GID>1513</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>446.5,-5364.5,459.5,-5364.5</points>
<connection>
<GID>1696</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>448.5,-5156.5,459.5,-5156.5</points>
<connection>
<GID>1644</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>447.5,-5442.5,459.5,-5442.5</points>
<connection>
<GID>1565</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>450.5,-5532.5,459.5,-5532.5</points>
<connection>
<GID>1539</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>441,-5770,459.5,-5770</points>
<connection>
<GID>1827</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>444,-5860,459.5,-5860</points>
<connection>
<GID>1801</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>445,-5938,459.5,-5938</points>
<connection>
<GID>1879</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>448,-6028,459.5,-6028</points>
<connection>
<GID>1853</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>443,-6146,459.5,-6146</points>
<connection>
<GID>1722</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>446,-6236,459.5,-6236</points>
<connection>
<GID>1905</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>447,-6314,459.5,-6314</points>
<connection>
<GID>1774</GID>
<name>OUT_0</name></connection>
<intersection>459.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>1463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543,-550.5,543,421.5</points>
<intersection>-550.5 23</intersection>
<intersection>-460.5 21</intersection>
<intersection>-269 19</intersection>
<intersection>-181.5 17</intersection>
<intersection>-101 14</intersection>
<intersection>-11 12</intersection>
<intersection>107 9</intersection>
<intersection>197 7</intersection>
<intersection>275 5</intersection>
<intersection>365 3</intersection>
<intersection>421.5 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>530.5,365,543,365</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>533.5,275,543,275</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>534.5,197,543,197</points>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>537.5,107,543,107</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>543,421.5,543.5,421.5</points>
<connection>
<GID>2140</GID>
<name>IN_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>532.5,-11,543,-11</points>
<connection>
<GID>400</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>535.5,-101,543,-101</points>
<connection>
<GID>374</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>525,-181.5,543,-181.5</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<connection>
<GID>452</GID>
<name>ENABLE_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>539.5,-269,543,-269</points>
<connection>
<GID>426</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>530.5,-460.5,543,-460.5</points>
<connection>
<GID>576</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>533.5,-550.5,543.5,-550.5</points>
<connection>
<GID>550</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection>
<intersection>543.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>543.5,-6406,543.5,-550.5</points>
<intersection>-6406 25</intersection>
<intersection>-6316 80</intersection>
<intersection>-6238 77</intersection>
<intersection>-6148 78</intersection>
<intersection>-6030 79</intersection>
<intersection>-5940 74</intersection>
<intersection>-5862 75</intersection>
<intersection>-5772 76</intersection>
<intersection>-5534.5 73</intersection>
<intersection>-5444.5 72</intersection>
<intersection>-5366.5 67</intersection>
<intersection>-5276.5 66</intersection>
<intersection>-5158.5 65</intersection>
<intersection>-4990.5 68</intersection>
<intersection>-4900.5 64</intersection>
<intersection>-4610 63</intersection>
<intersection>-4520 62</intersection>
<intersection>-4442 61</intersection>
<intersection>-4352 60</intersection>
<intersection>-4234 59</intersection>
<intersection>-4144 58</intersection>
<intersection>-3976 57</intersection>
<intersection>-3784.5 56</intersection>
<intersection>-3694.5 55</intersection>
<intersection>-3616.5 54</intersection>
<intersection>-3526.5 52</intersection>
<intersection>-3408.5 53</intersection>
<intersection>-3318.5 51</intersection>
<intersection>-3240.5 50</intersection>
<intersection>-3150.5 49</intersection>
<intersection>-2890.5 48</intersection>
<intersection>-2800.5 47</intersection>
<intersection>-2722.5 46</intersection>
<intersection>-2632.5 45</intersection>
<intersection>-2514.5 44</intersection>
<intersection>-2503 43</intersection>
<intersection>-2424.5 41</intersection>
<intersection>-2346.5 40</intersection>
<intersection>-2256.5 42</intersection>
<intersection>-2019 39</intersection>
<intersection>-1929 38</intersection>
<intersection>-1851 37</intersection>
<intersection>-1761 36</intersection>
<intersection>-1643 35</intersection>
<intersection>-1553 34</intersection>
<intersection>-1475 33</intersection>
<intersection>-1385 32</intersection>
<intersection>-1094.5 26</intersection>
<intersection>-1004.5 27</intersection>
<intersection>-926.5 28</intersection>
<intersection>-836.5 29</intersection>
<intersection>-718.5 31</intersection>
<intersection>-628.5 30</intersection>
<intersection>-550.5 23</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>534.5,-6406,543.5,-6406</points>
<connection>
<GID>1751</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>539.5,-1094.5,543.5,-1094.5</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>536.5,-1004.5,543.5,-1004.5</points>
<connection>
<GID>523</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>535.5,-926.5,543.5,-926.5</points>
<connection>
<GID>654</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>532.5,-836.5,543.5,-836.5</points>
<connection>
<GID>471</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>534.5,-628.5,543.5,-628.5</points>
<connection>
<GID>628</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>537.5,-718.5,543.5,-718.5</points>
<connection>
<GID>602</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>528,-1385,543.5,-1385</points>
<connection>
<GID>785</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>531,-1475,543.5,-1475</points>
<connection>
<GID>759</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>532,-1553,543.5,-1553</points>
<connection>
<GID>837</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>535,-1643,543.5,-1643</points>
<connection>
<GID>811</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>530,-1761,543.5,-1761</points>
<connection>
<GID>680</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>533,-1851,543.5,-1851</points>
<connection>
<GID>863</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>534,-1929,543.5,-1929</points>
<connection>
<GID>732</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>537,-2019,543.5,-2019</points>
<connection>
<GID>706</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>530.5,-2346.5,543.5,-2346.5</points>
<connection>
<GID>968</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>531.5,-2424.5,543.5,-2424.5</points>
<connection>
<GID>1046</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>527.5,-2256.5,543.5,-2256.5</points>
<connection>
<GID>994</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>543.5,-2503,580.5,-2503</points>
<connection>
<GID>1022</GID>
<name>IN_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>534.5,-2514.5,543.5,-2514.5</points>
<connection>
<GID>1020</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>529.5,-2632.5,543.5,-2632.5</points>
<connection>
<GID>889</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>532.5,-2722.5,543.5,-2722.5</points>
<connection>
<GID>1072</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>533.5,-2800.5,543.5,-2800.5</points>
<connection>
<GID>941</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>536.5,-2890.5,543.5,-2890.5</points>
<connection>
<GID>915</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>528.5,-3150.5,543.5,-3150.5</points>
<connection>
<GID>1133</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>531.5,-3240.5,543.5,-3240.5</points>
<connection>
<GID>1107</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>532.5,-3318.5,543.5,-3318.5</points>
<connection>
<GID>1185</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>530.5,-3526.5,543.5,-3526.5</points>
<connection>
<GID>1237</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>535.5,-3408.5,543.5,-3408.5</points>
<connection>
<GID>1159</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>533.5,-3616.5,543.5,-3616.5</points>
<connection>
<GID>1211</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>534.5,-3694.5,543.5,-3694.5</points>
<connection>
<GID>1289</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>537.5,-3784.5,543.5,-3784.5</points>
<connection>
<GID>1263</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>528.5,-3976,543.5,-3976</points>
<connection>
<GID>1412</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>532.5,-4144,543.5,-4144</points>
<connection>
<GID>1464</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>535.5,-4234,543.5,-4234</points>
<connection>
<GID>1438</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>530.5,-4352,543.5,-4352</points>
<connection>
<GID>1307</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>533.5,-4442,543.5,-4442</points>
<connection>
<GID>1490</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>534.5,-4520,543.5,-4520</points>
<connection>
<GID>1359</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>537.5,-4610,543.5,-4610</points>
<connection>
<GID>1333</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>526,-4900.5,543.5,-4900.5</points>
<connection>
<GID>1621</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>533,-5158.5,543.5,-5158.5</points>
<connection>
<GID>1647</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>528,-5276.5,543.5,-5276.5</points>
<connection>
<GID>1516</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>531,-5366.5,543.5,-5366.5</points>
<connection>
<GID>1699</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>529,-4990.5,543.5,-4990.5</points>
<connection>
<GID>1595</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>518.5,-5071,528,-5071</points>
<connection>
<GID>1674</GID>
<name>OUT</name></connection>
<connection>
<GID>1673</GID>
<name>ENABLE_0</name></connection></hsegment>
<hsegment>
<ID>72</ID>
<points>532,-5444.5,543.5,-5444.5</points>
<connection>
<GID>1568</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>535,-5534.5,543.5,-5534.5</points>
<connection>
<GID>1542</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>529.5,-5940,543.5,-5940</points>
<connection>
<GID>1882</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>528.5,-5862,543.5,-5862</points>
<connection>
<GID>1804</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>525.5,-5772,543.5,-5772</points>
<connection>
<GID>1830</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>530.5,-6238,543.5,-6238</points>
<connection>
<GID>1908</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>527.5,-6148,543.5,-6148</points>
<connection>
<GID>1725</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>532.5,-6030,543.5,-6030</points>
<connection>
<GID>1856</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment>
<hsegment>
<ID>80</ID>
<points>531.5,-6316,543.5,-6316</points>
<connection>
<GID>1777</GID>
<name>OUT_0</name></connection>
<intersection>543.5 24</intersection></hsegment></shape></wire>
<wire>
<ID>1464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619.5,-550.5,619.5,422</points>
<connection>
<GID>2144</GID>
<name>IN_0</name></connection>
<intersection>-550.5 21</intersection>
<intersection>-460.5 19</intersection>
<intersection>-269 17</intersection>
<intersection>-179 15</intersection>
<intersection>-101 13</intersection>
<intersection>-11 11</intersection>
<intersection>107 9</intersection>
<intersection>197 7</intersection>
<intersection>275 5</intersection>
<intersection>365 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>604,365,619.5,365</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>607,275,619.5,275</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>608,197,619.5,197</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>611,107,619.5,107</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>606,-11,619.5,-11</points>
<connection>
<GID>403</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>609,-101,619.5,-101</points>
<connection>
<GID>377</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>610,-179,619.5,-179</points>
<connection>
<GID>455</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>613,-269,619.5,-269</points>
<connection>
<GID>429</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>604,-460.5,619.5,-460.5</points>
<connection>
<GID>579</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>607,-550.5,620.5,-550.5</points>
<connection>
<GID>553</GID>
<name>OUT_0</name></connection>
<intersection>619.5 0</intersection>
<intersection>620.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>620.5,-6238,620.5,-550.5</points>
<intersection>-6238 23</intersection>
<intersection>-6148 77</intersection>
<intersection>-6030 78</intersection>
<intersection>-5940 76</intersection>
<intersection>-5862 75</intersection>
<intersection>-5772 74</intersection>
<intersection>-5534.5 73</intersection>
<intersection>-5444.5 72</intersection>
<intersection>-5366.5 71</intersection>
<intersection>-5276.5 70</intersection>
<intersection>-5158.5 69</intersection>
<intersection>-5068.5 68</intersection>
<intersection>-4990.5 67</intersection>
<intersection>-4900.5 66</intersection>
<intersection>-4610 65</intersection>
<intersection>-4520 62</intersection>
<intersection>-4442 63</intersection>
<intersection>-4352 64</intersection>
<intersection>-4234 61</intersection>
<intersection>-4144 60</intersection>
<intersection>-4066 59</intersection>
<intersection>-3976 58</intersection>
<intersection>-3784.5 56</intersection>
<intersection>-3694.5 57</intersection>
<intersection>-3616.5 55</intersection>
<intersection>-3526.5 54</intersection>
<intersection>-3408.5 53</intersection>
<intersection>-3318.5 52</intersection>
<intersection>-3240.5 51</intersection>
<intersection>-3150.5 50</intersection>
<intersection>-2890.5 49</intersection>
<intersection>-2800.5 48</intersection>
<intersection>-2722.5 47</intersection>
<intersection>-2632.5 46</intersection>
<intersection>-2514.5 45</intersection>
<intersection>-2424.5 44</intersection>
<intersection>-2346.5 43</intersection>
<intersection>-2256.5 42</intersection>
<intersection>-2019 41</intersection>
<intersection>-1929 40</intersection>
<intersection>-1851 39</intersection>
<intersection>-1761 38</intersection>
<intersection>-1643 37</intersection>
<intersection>-1553 36</intersection>
<intersection>-1475 35</intersection>
<intersection>-1385 34</intersection>
<intersection>-1094.5 29</intersection>
<intersection>-1004.5 28</intersection>
<intersection>-926.5 27</intersection>
<intersection>-836.5 26</intersection>
<intersection>-718.5 25</intersection>
<intersection>-628.5 24</intersection>
<intersection>-550.5 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>604,-6238,621,-6238</points>
<connection>
<GID>1911</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection>
<intersection>621 30</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>608,-628.5,620.5,-628.5</points>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>611,-718.5,620.5,-718.5</points>
<connection>
<GID>605</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>606,-836.5,620.5,-836.5</points>
<connection>
<GID>474</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>609,-926.5,620.5,-926.5</points>
<connection>
<GID>657</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>610,-1004.5,620.5,-1004.5</points>
<connection>
<GID>526</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>613,-1094.5,620.5,-1094.5</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>621,-6406,621,-6238</points>
<intersection>-6406 33</intersection>
<intersection>-6316 31</intersection>
<intersection>-6238 23</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>605,-6316,621,-6316</points>
<connection>
<GID>1780</GID>
<name>OUT_0</name></connection>
<intersection>621 30</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>608,-6406,621,-6406</points>
<connection>
<GID>1754</GID>
<name>OUT_0</name></connection>
<intersection>621 30</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>601.5,-1385,620.5,-1385</points>
<connection>
<GID>788</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>604.5,-1475,620.5,-1475</points>
<connection>
<GID>762</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>605.5,-1553,620.5,-1553</points>
<connection>
<GID>840</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>608.5,-1643,620.5,-1643</points>
<connection>
<GID>814</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>603.5,-1761,620.5,-1761</points>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>606.5,-1851,620.5,-1851</points>
<connection>
<GID>866</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>607.5,-1929,620.5,-1929</points>
<connection>
<GID>735</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>610.5,-2019,620.5,-2019</points>
<connection>
<GID>709</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>601,-2256.5,620.5,-2256.5</points>
<connection>
<GID>997</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>604,-2346.5,620.5,-2346.5</points>
<connection>
<GID>971</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>605,-2424.5,620.5,-2424.5</points>
<connection>
<GID>1049</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>608,-2514.5,620.5,-2514.5</points>
<connection>
<GID>1023</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>603,-2632.5,620.5,-2632.5</points>
<connection>
<GID>892</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>606,-2722.5,620.5,-2722.5</points>
<connection>
<GID>1075</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>607,-2800.5,620.5,-2800.5</points>
<connection>
<GID>944</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>610,-2890.5,620.5,-2890.5</points>
<connection>
<GID>918</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>602,-3150.5,620.5,-3150.5</points>
<connection>
<GID>1136</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>605,-3240.5,620.5,-3240.5</points>
<connection>
<GID>1110</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>606,-3318.5,620.5,-3318.5</points>
<connection>
<GID>1188</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>609,-3408.5,620.5,-3408.5</points>
<connection>
<GID>1162</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>604,-3526.5,620.5,-3526.5</points>
<connection>
<GID>1240</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>607,-3616.5,620.5,-3616.5</points>
<connection>
<GID>1214</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>611,-3784.5,620.5,-3784.5</points>
<connection>
<GID>1266</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>608,-3694.5,620.5,-3694.5</points>
<connection>
<GID>1292</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>602,-3976,620.5,-3976</points>
<connection>
<GID>1415</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>605,-4066,620.5,-4066</points>
<connection>
<GID>1389</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>606,-4144,620.5,-4144</points>
<connection>
<GID>1467</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>609,-4234,620.5,-4234</points>
<connection>
<GID>1441</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>608,-4520,620.5,-4520</points>
<connection>
<GID>1362</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>607,-4442,620.5,-4442</points>
<connection>
<GID>1493</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>604,-4352,620.5,-4352</points>
<connection>
<GID>1310</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>611,-4610,620.5,-4610</points>
<connection>
<GID>1336</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>599.5,-4900.5,620.5,-4900.5</points>
<connection>
<GID>1624</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>602.5,-4990.5,620.5,-4990.5</points>
<connection>
<GID>1598</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>603.5,-5068.5,620.5,-5068.5</points>
<connection>
<GID>1676</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>606.5,-5158.5,620.5,-5158.5</points>
<connection>
<GID>1650</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>601.5,-5276.5,620.5,-5276.5</points>
<connection>
<GID>1519</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>604.5,-5366.5,620.5,-5366.5</points>
<connection>
<GID>1702</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>605.5,-5444.5,620.5,-5444.5</points>
<connection>
<GID>1571</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>608.5,-5534.5,620.5,-5534.5</points>
<connection>
<GID>1545</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>599,-5772,620.5,-5772</points>
<connection>
<GID>1833</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>602,-5862,620.5,-5862</points>
<connection>
<GID>1807</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>603,-5940,620.5,-5940</points>
<connection>
<GID>1885</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>601,-6148,620.5,-6148</points>
<connection>
<GID>1728</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>606,-6030,620.5,-6030</points>
<connection>
<GID>1859</GID>
<name>OUT_0</name></connection>
<intersection>620.5 22</intersection></hsegment></shape></wire>
<wire>
<ID>1465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-6438.5,13,376.5</points>
<connection>
<GID>2098</GID>
<name>OUT_0</name></connection>
<intersection>-6394.5 70</intersection>
<intersection>-6304.5 69</intersection>
<intersection>-6226.5 66</intersection>
<intersection>-6136.5 67</intersection>
<intersection>-6018.5 68</intersection>
<intersection>-5928.5 65</intersection>
<intersection>-5850.5 64</intersection>
<intersection>-5760.5 63</intersection>
<intersection>-5523 62</intersection>
<intersection>-5433 61</intersection>
<intersection>-5355 60</intersection>
<intersection>-5265 59</intersection>
<intersection>-5147 58</intersection>
<intersection>-5057 51</intersection>
<intersection>-4979 50</intersection>
<intersection>-4889 49</intersection>
<intersection>-4598.5 48</intersection>
<intersection>-4508.5 47</intersection>
<intersection>-4430.5 45</intersection>
<intersection>-4340.5 46</intersection>
<intersection>-4222.5 44</intersection>
<intersection>-4132.5 42</intersection>
<intersection>-4054.5 43</intersection>
<intersection>-3964.5 41</intersection>
<intersection>-3773 40</intersection>
<intersection>-3683 39</intersection>
<intersection>-3605 38</intersection>
<intersection>-3515 37</intersection>
<intersection>-3397 36</intersection>
<intersection>-3307 35</intersection>
<intersection>-3229 34</intersection>
<intersection>-3139 33</intersection>
<intersection>-2879 32</intersection>
<intersection>-2789 31</intersection>
<intersection>-2711 30</intersection>
<intersection>-2621 29</intersection>
<intersection>-2503 28</intersection>
<intersection>-2413 27</intersection>
<intersection>-2335 26</intersection>
<intersection>-2245 25</intersection>
<intersection>-2007.5 24</intersection>
<intersection>-1917.5 23</intersection>
<intersection>-1839.5 21</intersection>
<intersection>-1749.5 22</intersection>
<intersection>-1631.5 18</intersection>
<intersection>-1541.5 19</intersection>
<intersection>-1463.5 20</intersection>
<intersection>-1373.5 17</intersection>
<intersection>-1083 16</intersection>
<intersection>-993 13</intersection>
<intersection>-915 14</intersection>
<intersection>-825 15</intersection>
<intersection>-707 12</intersection>
<intersection>-617 11</intersection>
<intersection>-539 9</intersection>
<intersection>-449 10</intersection>
<intersection>-257.5 8</intersection>
<intersection>-167.5 7</intersection>
<intersection>-89.5 6</intersection>
<intersection>0.5 5</intersection>
<intersection>118.5 4</intersection>
<intersection>208.5 3</intersection>
<intersection>286.5 2</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,376.5,22,376.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,286.5,25,286.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13,208.5,26,208.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>13,118.5,29,118.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>13,0.5,24,0.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>13,-89.5,27,-89.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>13,-167.5,28,-167.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>13,-257.5,31,-257.5</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>13,-539,25,-539</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>13,-449,22,-449</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>13,-617,26,-617</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>13,-707,29,-707</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>13,-993,28,-993</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>13,-915,27,-915</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>13,-825,24,-825</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>13,-1083,31,-1083</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>13,-1373.5,19.5,-1373.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>13,-1631.5,26.5,-1631.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>13,-1541.5,23.5,-1541.5</points>
<connection>
<GID>818</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>13,-1463.5,22.5,-1463.5</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>13,-1839.5,24.5,-1839.5</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>13,-1749.5,21.5,-1749.5</points>
<connection>
<GID>870</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>13,-1917.5,25.5,-1917.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>13,-2007.5,28.5,-2007.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>13,-2245,19,-2245</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>13,-2335,22,-2335</points>
<connection>
<GID>949</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>13,-2413,23,-2413</points>
<connection>
<GID>1027</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>13,-2503,26,-2503</points>
<connection>
<GID>1001</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>13,-2621,21,-2621</points>
<connection>
<GID>1079</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>13,-2711,24,-2711</points>
<connection>
<GID>1053</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>13,-2789,25,-2789</points>
<connection>
<GID>922</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>13,-2879,28,-2879</points>
<connection>
<GID>896</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>13,-3139,20,-3139</points>
<connection>
<GID>1114</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>13,-3229,23,-3229</points>
<connection>
<GID>1088</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>13,-3307,24,-3307</points>
<connection>
<GID>1166</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>13,-3397,27,-3397</points>
<connection>
<GID>1140</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>13,-3515,22,-3515</points>
<connection>
<GID>1218</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>13,-3605,25,-3605</points>
<connection>
<GID>1192</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>13,-3683,26,-3683</points>
<connection>
<GID>1270</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>13,-3773,29,-3773</points>
<connection>
<GID>1244</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>13,-3964.5,20,-3964.5</points>
<connection>
<GID>1393</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>13,-4132.5,24,-4132.5</points>
<connection>
<GID>1445</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>13,-4054.5,23,-4054.5</points>
<connection>
<GID>1367</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>13,-4222.5,27,-4222.5</points>
<connection>
<GID>1419</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>13,-4430.5,25,-4430.5</points>
<connection>
<GID>1471</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>13,-4340.5,22,-4340.5</points>
<connection>
<GID>1497</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>13,-4508.5,26,-4508.5</points>
<connection>
<GID>1340</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>13,-4598.5,29,-4598.5</points>
<connection>
<GID>1314</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>13,-4889,17.5,-4889</points>
<connection>
<GID>1602</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>13,-4979,20.5,-4979</points>
<connection>
<GID>1576</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>13,-5057,21.5,-5057</points>
<connection>
<GID>1654</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>13,-5147,24.5,-5147</points>
<connection>
<GID>1628</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>13,-5265,19.5,-5265</points>
<connection>
<GID>1706</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>13,-5355,22.5,-5355</points>
<connection>
<GID>1680</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>13,-5433,23.5,-5433</points>
<connection>
<GID>1549</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>13,-5523,26.5,-5523</points>
<connection>
<GID>1523</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>13,-5760.5,17,-5760.5</points>
<connection>
<GID>1811</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>13,-5850.5,20,-5850.5</points>
<connection>
<GID>1785</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>13,-5928.5,21,-5928.5</points>
<connection>
<GID>1863</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>13,-6226.5,22,-6226.5</points>
<connection>
<GID>1889</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>13,-6136.5,19,-6136.5</points>
<connection>
<GID>1915</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>13,-6018.5,24,-6018.5</points>
<connection>
<GID>1837</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>13,-6304.5,23,-6304.5</points>
<connection>
<GID>1758</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>13,-6394.5,26,-6394.5</points>
<connection>
<GID>1732</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>1466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-6439,74.5,376.5</points>
<intersection>-6439 2</intersection>
<intersection>-6394.5 68</intersection>
<intersection>-6304.5 67</intersection>
<intersection>-6226.5 66</intersection>
<intersection>-6136.5 65</intersection>
<intersection>-6018.5 64</intersection>
<intersection>-5928.5 63</intersection>
<intersection>-5850.5 62</intersection>
<intersection>-5760.5 61</intersection>
<intersection>-5523 60</intersection>
<intersection>-5433 59</intersection>
<intersection>-5355 58</intersection>
<intersection>-5265 57</intersection>
<intersection>-5147 56</intersection>
<intersection>-5057 52</intersection>
<intersection>-4979 51</intersection>
<intersection>-4889 50</intersection>
<intersection>-4598.5 49</intersection>
<intersection>-4508.5 48</intersection>
<intersection>-4430.5 47</intersection>
<intersection>-4340.5 46</intersection>
<intersection>-4222.5 44</intersection>
<intersection>-4132.5 45</intersection>
<intersection>-4054.5 43</intersection>
<intersection>-3964.5 42</intersection>
<intersection>-3773 41</intersection>
<intersection>-3683 40</intersection>
<intersection>-3605 39</intersection>
<intersection>-3515 38</intersection>
<intersection>-3397 37</intersection>
<intersection>-3307 34</intersection>
<intersection>-3229 35</intersection>
<intersection>-3139 36</intersection>
<intersection>-2879 33</intersection>
<intersection>-2789 32</intersection>
<intersection>-2711 31</intersection>
<intersection>-2621 30</intersection>
<intersection>-2503 29</intersection>
<intersection>-2413 28</intersection>
<intersection>-2335 27</intersection>
<intersection>-2245 26</intersection>
<intersection>-2007.5 25</intersection>
<intersection>-1917.5 24</intersection>
<intersection>-1839.5 23</intersection>
<intersection>-1749.5 22</intersection>
<intersection>-1631.5 21</intersection>
<intersection>-1541.5 20</intersection>
<intersection>-1463.5 19</intersection>
<intersection>-1373.5 18</intersection>
<intersection>-1083 17</intersection>
<intersection>-993 16</intersection>
<intersection>-915 15</intersection>
<intersection>-825 14</intersection>
<intersection>-707 13</intersection>
<intersection>-617 12</intersection>
<intersection>-539 11</intersection>
<intersection>-449 10</intersection>
<intersection>-257.5 9</intersection>
<intersection>-167.5 8</intersection>
<intersection>-89.5 7</intersection>
<intersection>0.5 6</intersection>
<intersection>118.5 5</intersection>
<intersection>208.5 4</intersection>
<intersection>286.5 3</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,376.5,95.5,376.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-6439,75.5,-6439</points>
<connection>
<GID>2101</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,286.5,98.5,286.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>74.5,208.5,99.5,208.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74.5,118.5,102.5,118.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>74.5,0.5,97.5,0.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>74.5,-89.5,97.5,-89.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>74.5,-167.5,101.5,-167.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>74.5,-257.5,104.5,-257.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>74.5,-449,95.5,-449</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>74.5,-539,98.5,-539</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>74.5,-617,99.5,-617</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>74.5,-707,102.5,-707</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>74.5,-825,97.5,-825</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>74.5,-915,100.5,-915</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>74.5,-993,101.5,-993</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>74.5,-1083,104.5,-1083</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>74.5,-1373.5,93,-1373.5</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>74.5,-1463.5,96,-1463.5</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>74.5,-1541.5,97,-1541.5</points>
<connection>
<GID>821</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>74.5,-1631.5,100,-1631.5</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>74.5,-1749.5,95,-1749.5</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>74.5,-1839.5,98,-1839.5</points>
<connection>
<GID>847</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>74.5,-1917.5,99,-1917.5</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>74.5,-2007.5,102,-2007.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>74.5,-2245,92.5,-2245</points>
<connection>
<GID>978</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>74.5,-2335,95.5,-2335</points>
<connection>
<GID>952</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>74.5,-2413,96.5,-2413</points>
<connection>
<GID>1030</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>74.5,-2503,99.5,-2503</points>
<connection>
<GID>1004</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>74.5,-2621,94.5,-2621</points>
<connection>
<GID>1082</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>74.5,-2711,97.5,-2711</points>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>74.5,-2789,98.5,-2789</points>
<connection>
<GID>925</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>74.5,-2879,101.5,-2879</points>
<connection>
<GID>899</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>74.5,-3307,97.5,-3307</points>
<connection>
<GID>1169</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>74.5,-3229,96.5,-3229</points>
<connection>
<GID>1091</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>74.5,-3139,93.5,-3139</points>
<connection>
<GID>1117</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>74.5,-3397,100.5,-3397</points>
<connection>
<GID>1143</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>74.5,-3515,95.5,-3515</points>
<connection>
<GID>1221</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>74.5,-3605,98.5,-3605</points>
<connection>
<GID>1195</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>74.5,-3683,99.5,-3683</points>
<connection>
<GID>1273</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>74.5,-3773,102.5,-3773</points>
<connection>
<GID>1247</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>74.5,-3964.5,93.5,-3964.5</points>
<connection>
<GID>1396</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>74.5,-4054.5,96.5,-4054.5</points>
<connection>
<GID>1370</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>74.5,-4222.5,100.5,-4222.5</points>
<connection>
<GID>1422</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>74.5,-4132.5,97.5,-4132.5</points>
<connection>
<GID>1448</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>74.5,-4340.5,95.5,-4340.5</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>74.5,-4430.5,98.5,-4430.5</points>
<connection>
<GID>1474</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>74.5,-4508.5,99.5,-4508.5</points>
<connection>
<GID>1343</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>74.5,-4598.5,102.5,-4598.5</points>
<connection>
<GID>1317</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>74.5,-4889,91,-4889</points>
<connection>
<GID>1605</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>74.5,-4979,94,-4979</points>
<connection>
<GID>1579</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>74.5,-5057,95,-5057</points>
<connection>
<GID>1657</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>74.5,-5147,98,-5147</points>
<connection>
<GID>1631</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>74.5,-5265,93,-5265</points>
<connection>
<GID>1709</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>74.5,-5355,96,-5355</points>
<connection>
<GID>1683</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>74.5,-5433,97,-5433</points>
<connection>
<GID>1552</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>74.5,-5523,100,-5523</points>
<connection>
<GID>1526</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>74.5,-5760.5,90.5,-5760.5</points>
<connection>
<GID>1814</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>74.5,-5850.5,93.5,-5850.5</points>
<connection>
<GID>1788</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>74.5,-5928.5,94.5,-5928.5</points>
<connection>
<GID>1866</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>74.5,-6018.5,97.5,-6018.5</points>
<connection>
<GID>1840</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>74.5,-6136.5,92.5,-6136.5</points>
<connection>
<GID>1918</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>74.5,-6226.5,95.5,-6226.5</points>
<connection>
<GID>1892</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>74.5,-6304.5,96.5,-6304.5</points>
<connection>
<GID>1761</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>74.5,-6394.5,99.5,-6394.5</points>
<connection>
<GID>1735</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-6439,152,376.5</points>
<connection>
<GID>2103</GID>
<name>OUT_0</name></connection>
<intersection>-6394.5 67</intersection>
<intersection>-6304.5 66</intersection>
<intersection>-6226.5 63</intersection>
<intersection>-6136.5 64</intersection>
<intersection>-6018.5 65</intersection>
<intersection>-5928.5 62</intersection>
<intersection>-5850.5 61</intersection>
<intersection>-5760.5 60</intersection>
<intersection>-5523 58</intersection>
<intersection>-5433 59</intersection>
<intersection>-5355 57</intersection>
<intersection>-5265 56</intersection>
<intersection>-5147 55</intersection>
<intersection>-5057 51</intersection>
<intersection>-4979 50</intersection>
<intersection>-4889 49</intersection>
<intersection>-4598.5 48</intersection>
<intersection>-4508.5 47</intersection>
<intersection>-4430.5 46</intersection>
<intersection>-4340.5 45</intersection>
<intersection>-4222.5 44</intersection>
<intersection>-4132.5 43</intersection>
<intersection>-4054.5 42</intersection>
<intersection>-3964.5 41</intersection>
<intersection>-3773 40</intersection>
<intersection>-3683 39</intersection>
<intersection>-3605 37</intersection>
<intersection>-3515 36</intersection>
<intersection>-3397 38</intersection>
<intersection>-3307 35</intersection>
<intersection>-3229 34</intersection>
<intersection>-3139 33</intersection>
<intersection>-2879 31</intersection>
<intersection>-2789 32</intersection>
<intersection>-2711 30</intersection>
<intersection>-2621 29</intersection>
<intersection>-2503 28</intersection>
<intersection>-2413 25</intersection>
<intersection>-2335 26</intersection>
<intersection>-2245 27</intersection>
<intersection>-2007.5 24</intersection>
<intersection>-1917.5 23</intersection>
<intersection>-1839.5 21</intersection>
<intersection>-1749.5 22</intersection>
<intersection>-1631.5 20</intersection>
<intersection>-1541.5 19</intersection>
<intersection>-1463.5 18</intersection>
<intersection>-1373.5 17</intersection>
<intersection>-1083 16</intersection>
<intersection>-993 13</intersection>
<intersection>-915 14</intersection>
<intersection>-825 15</intersection>
<intersection>-707 12</intersection>
<intersection>-617 11</intersection>
<intersection>-539 9</intersection>
<intersection>-449 10</intersection>
<intersection>-257.5 8</intersection>
<intersection>-167.5 7</intersection>
<intersection>-89.5 6</intersection>
<intersection>0.5 4</intersection>
<intersection>118.5 5</intersection>
<intersection>208.5 3</intersection>
<intersection>286.5 2</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,376.5,180,376.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,286.5,183,286.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>152,208.5,184,208.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>152,0.5,182,0.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>152,118.5,187,118.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>152,-89.5,185,-89.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>152,-167.5,186,-167.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>152,-257.5,189,-257.5</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-539,183,-539</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>152,-449,180,-449</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>152,-617,184,-617</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>152,-707,187,-707</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>152,-993,186,-993</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>152,-915,185,-915</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>152,-825,182,-825</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>152,-1083,189,-1083</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>152,-1373.5,177.5,-1373.5</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>152,-1463.5,180.5,-1463.5</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>152,-1541.5,181.5,-1541.5</points>
<connection>
<GID>824</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>152,-1631.5,184.5,-1631.5</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>152,-1839.5,182.5,-1839.5</points>
<connection>
<GID>850</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>152,-1749.5,179.5,-1749.5</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>152,-1917.5,183.5,-1917.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>152,-2007.5,186.5,-2007.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>152,-2413,181,-2413</points>
<connection>
<GID>1033</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>152,-2335,180,-2335</points>
<connection>
<GID>955</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>152,-2245,177,-2245</points>
<connection>
<GID>981</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>152,-2503,184,-2503</points>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>152,-2621,179,-2621</points>
<connection>
<GID>1085</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>152,-2711,182,-2711</points>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>152,-2879,186,-2879</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>152,-2789,183,-2789</points>
<connection>
<GID>928</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>152,-3139,178,-3139</points>
<connection>
<GID>1120</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>152,-3229,181,-3229</points>
<connection>
<GID>1094</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>152,-3307,182,-3307</points>
<connection>
<GID>1172</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>152,-3515,180,-3515</points>
<connection>
<GID>1224</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>152,-3605,183,-3605</points>
<connection>
<GID>1198</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>152,-3397,185,-3397</points>
<connection>
<GID>1146</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>152,-3683,184,-3683</points>
<connection>
<GID>1276</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>152,-3773,187,-3773</points>
<connection>
<GID>1250</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>152,-3964.5,178,-3964.5</points>
<connection>
<GID>1399</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>152,-4054.5,181,-4054.5</points>
<connection>
<GID>1373</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>152,-4132.5,182,-4132.5</points>
<connection>
<GID>1451</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>152,-4222.5,185,-4222.5</points>
<connection>
<GID>1425</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>152,-4340.5,180,-4340.5</points>
<connection>
<GID>1503</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>152,-4430.5,183,-4430.5</points>
<connection>
<GID>1477</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>152,-4508.5,184,-4508.5</points>
<connection>
<GID>1346</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>152,-4598.5,187,-4598.5</points>
<connection>
<GID>1320</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>152,-4889,175.5,-4889</points>
<connection>
<GID>1608</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>152,-4979,178.5,-4979</points>
<connection>
<GID>1582</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>152,-5057,179.5,-5057</points>
<connection>
<GID>1660</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>152,-5147,182.5,-5147</points>
<connection>
<GID>1634</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>152,-5265,177.5,-5265</points>
<connection>
<GID>1712</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>152,-5355,180.5,-5355</points>
<connection>
<GID>1686</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>152,-5523,184.5,-5523</points>
<connection>
<GID>1529</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>152,-5433,181.5,-5433</points>
<connection>
<GID>1555</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>152,-5760.5,175,-5760.5</points>
<connection>
<GID>1817</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>152,-5850.5,178,-5850.5</points>
<connection>
<GID>1791</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>152,-5928.5,179,-5928.5</points>
<connection>
<GID>1869</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>152,-6226.5,180,-6226.5</points>
<connection>
<GID>1895</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>152,-6136.5,177,-6136.5</points>
<connection>
<GID>1921</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>152,-6018.5,182,-6018.5</points>
<connection>
<GID>1843</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>152,-6304.5,181,-6304.5</points>
<connection>
<GID>1764</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>152,-6394.5,184,-6394.5</points>
<connection>
<GID>1738</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>1468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-6439,234.5,376.5</points>
<connection>
<GID>2105</GID>
<name>OUT_0</name></connection>
<intersection>-6394.5 65</intersection>
<intersection>-6304.5 66</intersection>
<intersection>-6226.5 64</intersection>
<intersection>-6136.5 63</intersection>
<intersection>-6018.5 62</intersection>
<intersection>-5928.5 61</intersection>
<intersection>-5850.5 60</intersection>
<intersection>-5760.5 59</intersection>
<intersection>-5523 58</intersection>
<intersection>-5433 57</intersection>
<intersection>-5355 56</intersection>
<intersection>-5265 55</intersection>
<intersection>-5147 54</intersection>
<intersection>-5057 50</intersection>
<intersection>-4979 49</intersection>
<intersection>-4889 48</intersection>
<intersection>-4508.5 47</intersection>
<intersection>-4430.5 46</intersection>
<intersection>-4340.5 45</intersection>
<intersection>-4222.5 44</intersection>
<intersection>-4132.5 43</intersection>
<intersection>-4054.5 42</intersection>
<intersection>-3964.5 41</intersection>
<intersection>-3773 39</intersection>
<intersection>-3683 40</intersection>
<intersection>-3605 38</intersection>
<intersection>-3515 37</intersection>
<intersection>-3397 36</intersection>
<intersection>-3307 33</intersection>
<intersection>-3229 34</intersection>
<intersection>-3139 35</intersection>
<intersection>-2879 32</intersection>
<intersection>-2789 31</intersection>
<intersection>-2711 30</intersection>
<intersection>-2621 29</intersection>
<intersection>-2503 28</intersection>
<intersection>-2413 27</intersection>
<intersection>-2335 26</intersection>
<intersection>-2245 25</intersection>
<intersection>-2007.5 24</intersection>
<intersection>-1917.5 23</intersection>
<intersection>-1839.5 22</intersection>
<intersection>-1749.5 21</intersection>
<intersection>-1631.5 17</intersection>
<intersection>-1541.5 18</intersection>
<intersection>-1463.5 19</intersection>
<intersection>-1373.5 20</intersection>
<intersection>-1083 16</intersection>
<intersection>-993 15</intersection>
<intersection>-915 14</intersection>
<intersection>-825 13</intersection>
<intersection>-707 12</intersection>
<intersection>-617 11</intersection>
<intersection>-539 10</intersection>
<intersection>-449 9</intersection>
<intersection>-257.5 8</intersection>
<intersection>-167.5 7</intersection>
<intersection>-89.5 6</intersection>
<intersection>0.5 5</intersection>
<intersection>118.5 4</intersection>
<intersection>208.5 3</intersection>
<intersection>286.5 2</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,376.5,254.5,376.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234.5,286.5,257.5,286.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>234.5,208.5,258.5,208.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>234.5,118.5,261.5,118.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>234.5,0.5,256.5,0.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>234.5,-89.5,259.5,-89.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>234.5,-167.5,260.5,-167.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>234.5,-257.5,263.5,-257.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>234.5,-449,254.5,-449</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>234.5,-539,257.5,-539</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>234.5,-617,258.5,-617</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>234.5,-707,261.5,-707</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>234.5,-825,256.5,-825</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>234.5,-915,259.5,-915</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>234.5,-993,260.5,-993</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>234.5,-1083,263.5,-1083</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>234.5,-1631.5,259,-1631.5</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>234.5,-1541.5,256,-1541.5</points>
<connection>
<GID>827</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>234.5,-1463.5,255,-1463.5</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>234.5,-1373.5,252,-1373.5</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>234.5,-1749.5,254,-1749.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>234.5,-1839.5,257,-1839.5</points>
<connection>
<GID>853</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>234.5,-1917.5,258,-1917.5</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>234.5,-2007.5,261,-2007.5</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>234.5,-2245,251.5,-2245</points>
<connection>
<GID>984</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>234.5,-2335,254.5,-2335</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>234.5,-2413,255.5,-2413</points>
<connection>
<GID>1036</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>234.5,-2503,258.5,-2503</points>
<connection>
<GID>1010</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>234.5,-2621,253.5,-2621</points>
<connection>
<GID>879</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>234.5,-2711,256.5,-2711</points>
<connection>
<GID>1062</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>234.5,-2789,257.5,-2789</points>
<connection>
<GID>931</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>234.5,-2879,260.5,-2879</points>
<connection>
<GID>905</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>234.5,-3307,256.5,-3307</points>
<connection>
<GID>1175</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>234.5,-3229,255.5,-3229</points>
<connection>
<GID>1097</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>234.5,-3139,252.5,-3139</points>
<connection>
<GID>1123</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>234.5,-3397,259.5,-3397</points>
<connection>
<GID>1149</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>234.5,-3515,254.5,-3515</points>
<connection>
<GID>1227</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>234.5,-3605,257.5,-3605</points>
<connection>
<GID>1201</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>234.5,-3773,261.5,-3773</points>
<connection>
<GID>1253</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>234.5,-3683,258.5,-3683</points>
<connection>
<GID>1279</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>234.5,-3964.5,252.5,-3964.5</points>
<connection>
<GID>1402</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>234.5,-4054.5,255.5,-4054.5</points>
<connection>
<GID>1376</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>234.5,-4132.5,256.5,-4132.5</points>
<connection>
<GID>1454</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>234.5,-4222.5,259.5,-4222.5</points>
<connection>
<GID>1428</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>234.5,-4340.5,254.5,-4340.5</points>
<connection>
<GID>1297</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>234.5,-4430.5,256.5,-4430.5</points>
<connection>
<GID>1480</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>234.5,-4508.5,258.5,-4508.5</points>
<connection>
<GID>1349</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>234.5,-4889,250,-4889</points>
<connection>
<GID>1611</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>234.5,-4979,253,-4979</points>
<connection>
<GID>1585</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>234.5,-5057,254,-5057</points>
<connection>
<GID>1663</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>234.5,-5147,257,-5147</points>
<connection>
<GID>1637</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>234.5,-5265,252,-5265</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>234.5,-5355,255,-5355</points>
<connection>
<GID>1689</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>234.5,-5433,256,-5433</points>
<connection>
<GID>1558</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>234.5,-5523,259,-5523</points>
<connection>
<GID>1532</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>234.5,-5760.5,249.5,-5760.5</points>
<connection>
<GID>1820</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>234.5,-5850.5,252.5,-5850.5</points>
<connection>
<GID>1794</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>234.5,-5928.5,253.5,-5928.5</points>
<connection>
<GID>1872</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>234.5,-6018.5,256.5,-6018.5</points>
<connection>
<GID>1846</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>234.5,-6136.5,251.5,-6136.5</points>
<connection>
<GID>1715</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>234.5,-6226.5,254.5,-6226.5</points>
<connection>
<GID>1898</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>234.5,-6394.5,258.5,-6394.5</points>
<connection>
<GID>1741</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>234.5,-6304.5,255.5,-6304.5</points>
<connection>
<GID>1767</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-6439.5,308,376.5</points>
<connection>
<GID>2107</GID>
<name>OUT_0</name></connection>
<intersection>-6394.5 67</intersection>
<intersection>-6304.5 66</intersection>
<intersection>-6226.5 65</intersection>
<intersection>-6136.5 64</intersection>
<intersection>-6018.5 63</intersection>
<intersection>-5928.5 62</intersection>
<intersection>-5850.5 61</intersection>
<intersection>-5760.5 60</intersection>
<intersection>-5523 59</intersection>
<intersection>-5433 58</intersection>
<intersection>-5355 57</intersection>
<intersection>-5265 56</intersection>
<intersection>-5147 55</intersection>
<intersection>-5057 51</intersection>
<intersection>-4979 50</intersection>
<intersection>-4889 49</intersection>
<intersection>-4598.5 48</intersection>
<intersection>-4508.5 47</intersection>
<intersection>-4430.5 46</intersection>
<intersection>-4340.5 45</intersection>
<intersection>-4222.5 44</intersection>
<intersection>-4132.5 43</intersection>
<intersection>-4054.5 42</intersection>
<intersection>-3964.5 41</intersection>
<intersection>-3773 40</intersection>
<intersection>-3683 39</intersection>
<intersection>-3605 38</intersection>
<intersection>-3515 37</intersection>
<intersection>-3397 36</intersection>
<intersection>-3307 35</intersection>
<intersection>-3229 34</intersection>
<intersection>-3139 33</intersection>
<intersection>-2879 32</intersection>
<intersection>-2789 31</intersection>
<intersection>-2711 30</intersection>
<intersection>-2621 29</intersection>
<intersection>-2503 28</intersection>
<intersection>-2413 27</intersection>
<intersection>-2335 25</intersection>
<intersection>-2245 26</intersection>
<intersection>-2007.5 24</intersection>
<intersection>-1917.5 23</intersection>
<intersection>-1839.5 21</intersection>
<intersection>-1749.5 22</intersection>
<intersection>-1631.5 20</intersection>
<intersection>-1541.5 19</intersection>
<intersection>-1463.5 18</intersection>
<intersection>-1373.5 17</intersection>
<intersection>-1083 16</intersection>
<intersection>-993 15</intersection>
<intersection>-915 14</intersection>
<intersection>-825 13</intersection>
<intersection>-707 12</intersection>
<intersection>-617 11</intersection>
<intersection>-539 10</intersection>
<intersection>-449 9</intersection>
<intersection>-257.5 8</intersection>
<intersection>-167.5 7</intersection>
<intersection>-89.5 6</intersection>
<intersection>0.5 5</intersection>
<intersection>118.5 4</intersection>
<intersection>208.5 3</intersection>
<intersection>286.5 2</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308,376.5,345,376.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,286.5,348,286.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>308,208.5,349,208.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>308,118.5,352,118.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>308,0.5,347,0.5</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>308,-89.5,350,-89.5</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>308,-167.5,351,-167.5</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>308,-257.5,354,-257.5</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>308,-449,345,-449</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>308,-539,348,-539</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>308,-617,349,-617</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>308,-707,352,-707</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>308,-825,347,-825</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>308,-915,350,-915</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>308,-993,351,-993</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>308,-1083,354,-1083</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>308,-1373.5,342.5,-1373.5</points>
<connection>
<GID>778</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>308,-1463.5,345.5,-1463.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>308,-1541.5,346.5,-1541.5</points>
<connection>
<GID>830</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>308,-1631.5,349.5,-1631.5</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>308,-1839.5,347.5,-1839.5</points>
<connection>
<GID>856</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>308,-1749.5,344.5,-1749.5</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>308,-1917.5,348.5,-1917.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>308,-2007.5,351.5,-2007.5</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>308,-2335,345,-2335</points>
<connection>
<GID>961</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>308,-2245,342,-2245</points>
<connection>
<GID>987</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>308,-2413,346,-2413</points>
<connection>
<GID>1039</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>308,-2503,349,-2503</points>
<connection>
<GID>1013</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>308,-2621,344,-2621</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>308,-2711,347,-2711</points>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>308,-2789,348,-2789</points>
<connection>
<GID>934</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>308,-2879,351,-2879</points>
<connection>
<GID>908</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>308,-3139,343,-3139</points>
<connection>
<GID>1126</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>308,-3229,346,-3229</points>
<connection>
<GID>1100</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>308,-3307,347,-3307</points>
<connection>
<GID>1178</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>308,-3397,350,-3397</points>
<connection>
<GID>1152</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>308,-3515,345,-3515</points>
<connection>
<GID>1230</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>308,-3605,348,-3605</points>
<connection>
<GID>1204</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>308,-3683,349,-3683</points>
<connection>
<GID>1282</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>308,-3773,352,-3773</points>
<connection>
<GID>1256</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>308,-3964.5,343,-3964.5</points>
<connection>
<GID>1405</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>308,-4054.5,346,-4054.5</points>
<connection>
<GID>1379</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>308,-4132.5,347,-4132.5</points>
<connection>
<GID>1457</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>308,-4222.5,350,-4222.5</points>
<connection>
<GID>1431</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>308,-4340.5,345,-4340.5</points>
<connection>
<GID>1300</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>308,-4430.5,348,-4430.5</points>
<connection>
<GID>1483</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>308,-4508.5,349,-4508.5</points>
<connection>
<GID>1352</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>308,-4598.5,352,-4598.5</points>
<connection>
<GID>1326</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>308,-4889,340.5,-4889</points>
<connection>
<GID>1614</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>308,-4979,343.5,-4979</points>
<connection>
<GID>1588</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>308,-5057,344.5,-5057</points>
<connection>
<GID>1666</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>308,-5147,347.5,-5147</points>
<connection>
<GID>1640</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>308,-5265,342.5,-5265</points>
<connection>
<GID>1509</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>308,-5355,345.5,-5355</points>
<connection>
<GID>1692</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>308,-5433,346.5,-5433</points>
<connection>
<GID>1561</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>308,-5523,349.5,-5523</points>
<connection>
<GID>1535</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>308,-5760.5,340,-5760.5</points>
<connection>
<GID>1823</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>308,-5850.5,343,-5850.5</points>
<connection>
<GID>1797</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>308,-5928.5,344,-5928.5</points>
<connection>
<GID>1875</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>308,-6018.5,347,-6018.5</points>
<connection>
<GID>1849</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>308,-6136.5,342,-6136.5</points>
<connection>
<GID>1718</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>308,-6226.5,345,-6226.5</points>
<connection>
<GID>1901</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>308,-6304.5,346,-6304.5</points>
<connection>
<GID>1770</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>308,-6394.5,349,-6394.5</points>
<connection>
<GID>1744</GID>
<name>IN_0</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>1470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404,-6440,404,376.5</points>
<intersection>-6440 2</intersection>
<intersection>-6394.5 68</intersection>
<intersection>-6304.5 67</intersection>
<intersection>-6226.5 66</intersection>
<intersection>-6136.5 65</intersection>
<intersection>-6018.5 64</intersection>
<intersection>-5928.5 63</intersection>
<intersection>-5850.5 62</intersection>
<intersection>-5760.5 61</intersection>
<intersection>-5523 60</intersection>
<intersection>-5433 59</intersection>
<intersection>-5355 58</intersection>
<intersection>-5265 57</intersection>
<intersection>-5147 53</intersection>
<intersection>-5057 52</intersection>
<intersection>-4979 51</intersection>
<intersection>-4889 50</intersection>
<intersection>-4598.5 49</intersection>
<intersection>-4508.5 46</intersection>
<intersection>-4430.5 47</intersection>
<intersection>-4340.5 48</intersection>
<intersection>-4222.5 45</intersection>
<intersection>-4132.5 43</intersection>
<intersection>-4054.5 44</intersection>
<intersection>-3964.5 42</intersection>
<intersection>-3773 41</intersection>
<intersection>-3683 40</intersection>
<intersection>-3605 39</intersection>
<intersection>-3515 38</intersection>
<intersection>-3397 37</intersection>
<intersection>-3307 36</intersection>
<intersection>-3229 35</intersection>
<intersection>-3139 34</intersection>
<intersection>-2879 33</intersection>
<intersection>-2789 32</intersection>
<intersection>-2711 31</intersection>
<intersection>-2621 30</intersection>
<intersection>-2503 29</intersection>
<intersection>-2413 26</intersection>
<intersection>-2335 27</intersection>
<intersection>-2245 28</intersection>
<intersection>-2007.5 25</intersection>
<intersection>-1917.5 24</intersection>
<intersection>-1839.5 23</intersection>
<intersection>-1749.5 22</intersection>
<intersection>-1631.5 21</intersection>
<intersection>-1541.5 20</intersection>
<intersection>-1463.5 19</intersection>
<intersection>-1373.5 18</intersection>
<intersection>-1083 17</intersection>
<intersection>-993 16</intersection>
<intersection>-915 15</intersection>
<intersection>-825 14</intersection>
<intersection>-707 13</intersection>
<intersection>-617 12</intersection>
<intersection>-539 11</intersection>
<intersection>-449 10</intersection>
<intersection>-257.5 9</intersection>
<intersection>-167.5 8</intersection>
<intersection>-89.5 7</intersection>
<intersection>0.5 5</intersection>
<intersection>118.5 6</intersection>
<intersection>208.5 4</intersection>
<intersection>286.5 3</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>404,376.5,418.5,376.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>396.5,-6440,404,-6440</points>
<connection>
<GID>2109</GID>
<name>OUT_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>404,286.5,421.5,286.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>404,208.5,422.5,208.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>404,0.5,420.5,0.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>404,118.5,425.5,118.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>404,-89.5,423.5,-89.5</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>404,-167.5,424.5,-167.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>404,-257.5,427.5,-257.5</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>404,-449,418.5,-449</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>404,-539,421.5,-539</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>404,-617,422.5,-617</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>404,-707,425.5,-707</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>404,-825,420.5,-825</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>404,-915,423.5,-915</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>404,-993,424.5,-993</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>404,-1083,427.5,-1083</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>404,-1373.5,416,-1373.5</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>404,-1463.5,419,-1463.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>404,-1541.5,420,-1541.5</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>404,-1631.5,423,-1631.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>404,-1749.5,418,-1749.5</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>404,-1839.5,421,-1839.5</points>
<connection>
<GID>859</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>404,-1917.5,422,-1917.5</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>404,-2007.5,425,-2007.5</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>404,-2413,419.5,-2413</points>
<connection>
<GID>1042</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>404,-2335,418.5,-2335</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>404,-2245,415.5,-2245</points>
<connection>
<GID>990</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>404,-2503,422.5,-2503</points>
<connection>
<GID>1016</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>404,-2621,417.5,-2621</points>
<connection>
<GID>885</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>404,-2711,420.5,-2711</points>
<connection>
<GID>1068</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>404,-2789,421.5,-2789</points>
<connection>
<GID>937</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>404,-2879,424.5,-2879</points>
<connection>
<GID>911</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>404,-3139,416.5,-3139</points>
<connection>
<GID>1129</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>404,-3229,419.5,-3229</points>
<connection>
<GID>1103</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>404,-3307,420.5,-3307</points>
<connection>
<GID>1181</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>404,-3397,423.5,-3397</points>
<connection>
<GID>1155</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>404,-3515,418.5,-3515</points>
<connection>
<GID>1233</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>404,-3605,421.5,-3605</points>
<connection>
<GID>1207</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>404,-3683,422.5,-3683</points>
<connection>
<GID>1285</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>404,-3773,425.5,-3773</points>
<connection>
<GID>1259</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>404,-3964.5,416.5,-3964.5</points>
<connection>
<GID>1408</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>404,-4132.5,420.5,-4132.5</points>
<connection>
<GID>1460</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>404,-4054.5,419.5,-4054.5</points>
<connection>
<GID>1382</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>404,-4222.5,423.5,-4222.5</points>
<connection>
<GID>1434</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>404,-4508.5,422.5,-4508.5</points>
<connection>
<GID>1355</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>404,-4430.5,421.5,-4430.5</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>404,-4340.5,418.5,-4340.5</points>
<connection>
<GID>1303</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>404,-4598.5,425.5,-4598.5</points>
<connection>
<GID>1329</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>404,-4889,414,-4889</points>
<connection>
<GID>1617</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>404,-4979,417,-4979</points>
<connection>
<GID>1591</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>404,-5057,418,-5057</points>
<connection>
<GID>1669</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>404,-5147,421,-5147</points>
<connection>
<GID>1643</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>404,-5265,416,-5265</points>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>404,-5355,419,-5355</points>
<connection>
<GID>1695</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>404,-5433,420,-5433</points>
<connection>
<GID>1564</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>404,-5523,423,-5523</points>
<connection>
<GID>1538</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>404,-5760.5,413.5,-5760.5</points>
<connection>
<GID>1826</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>404,-5850.5,416.5,-5850.5</points>
<connection>
<GID>1800</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>404,-5928.5,417.5,-5928.5</points>
<connection>
<GID>1878</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>404,-6018.5,420.5,-6018.5</points>
<connection>
<GID>1852</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>65</ID>
<points>404,-6136.5,415.5,-6136.5</points>
<connection>
<GID>1721</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>404,-6226.5,418.5,-6226.5</points>
<connection>
<GID>1904</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>67</ID>
<points>404,-6304.5,419.5,-6304.5</points>
<connection>
<GID>1773</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>404,-6394.5,422.5,-6394.5</points>
<connection>
<GID>1747</GID>
<name>IN_0</name></connection>
<intersection>404 0</intersection></hsegment></shape></wire>
<wire>
<ID>1471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>478,-6440,478,376.5</points>
<connection>
<GID>2111</GID>
<name>OUT_0</name></connection>
<intersection>-6394.5 62</intersection>
<intersection>-6304.5 63</intersection>
<intersection>-6226.5 59</intersection>
<intersection>-6136.5 60</intersection>
<intersection>-6018.5 61</intersection>
<intersection>-5928.5 56</intersection>
<intersection>-5850.5 57</intersection>
<intersection>-5760.5 58</intersection>
<intersection>-5523 55</intersection>
<intersection>-5433 54</intersection>
<intersection>-5355 51</intersection>
<intersection>-5265 50</intersection>
<intersection>-5147 49</intersection>
<intersection>-5057 53</intersection>
<intersection>-4979 52</intersection>
<intersection>-4889 48</intersection>
<intersection>-4598.5 47</intersection>
<intersection>-4508.5 46</intersection>
<intersection>-4430.5 45</intersection>
<intersection>-4340.5 44</intersection>
<intersection>-4222.5 43</intersection>
<intersection>-4132.5 41</intersection>
<intersection>-4054.5 42</intersection>
<intersection>-3964.5 40</intersection>
<intersection>-3773 39</intersection>
<intersection>-3683 38</intersection>
<intersection>-3605 37</intersection>
<intersection>-3515 35</intersection>
<intersection>-3397 36</intersection>
<intersection>-3307 34</intersection>
<intersection>-3229 33</intersection>
<intersection>-3139 32</intersection>
<intersection>-2879 31</intersection>
<intersection>-2789 30</intersection>
<intersection>-2711 29</intersection>
<intersection>-2621 28</intersection>
<intersection>-2503 27</intersection>
<intersection>-2413 26</intersection>
<intersection>-2335 25</intersection>
<intersection>-2007.5 24</intersection>
<intersection>-1917.5 23</intersection>
<intersection>-1839.5 22</intersection>
<intersection>-1749.5 21</intersection>
<intersection>-1631.5 20</intersection>
<intersection>-1541.5 19</intersection>
<intersection>-1463.5 18</intersection>
<intersection>-1373.5 17</intersection>
<intersection>-1083 16</intersection>
<intersection>-993 15</intersection>
<intersection>-915 14</intersection>
<intersection>-825 13</intersection>
<intersection>-707 12</intersection>
<intersection>-617 11</intersection>
<intersection>-539 10</intersection>
<intersection>-449 9</intersection>
<intersection>-257.5 8</intersection>
<intersection>-167.5 7</intersection>
<intersection>-89.5 6</intersection>
<intersection>0.5 5</intersection>
<intersection>118.5 4</intersection>
<intersection>208.5 3</intersection>
<intersection>286.5 2</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478,376.5,503,376.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>478,286.5,506,286.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>478,208.5,507,208.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>478,118.5,510,118.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>478,0.5,505,0.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>478,-89.5,508,-89.5</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>478,-167.5,509,-167.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>478,-257.5,512,-257.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>478,-449,503,-449</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>478,-539,506,-539</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>478,-617,507,-617</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>478,-707,510,-707</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>478,-825,505,-825</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>478,-915,508,-915</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>478,-993,509,-993</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>478,-1083,512,-1083</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>478,-1373.5,500.5,-1373.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>478,-1463.5,503.5,-1463.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>478,-1541.5,504.5,-1541.5</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>478,-1631.5,507.5,-1631.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>478,-1749.5,502.5,-1749.5</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>478,-1839.5,505.5,-1839.5</points>
<connection>
<GID>862</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>478,-1917.5,506.5,-1917.5</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>478,-2007.5,509.5,-2007.5</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>478,-2335,503,-2335</points>
<connection>
<GID>967</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>478,-2413,504,-2413</points>
<connection>
<GID>1045</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>478,-2503,507,-2503</points>
<connection>
<GID>1019</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>478,-2621,502,-2621</points>
<connection>
<GID>888</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>478,-2711,505,-2711</points>
<connection>
<GID>1071</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>478,-2789,506,-2789</points>
<connection>
<GID>940</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>478,-2879,509,-2879</points>
<connection>
<GID>914</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>478,-3139,501,-3139</points>
<connection>
<GID>1132</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>478,-3229,504,-3229</points>
<connection>
<GID>1106</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>478,-3307,505,-3307</points>
<connection>
<GID>1184</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>478,-3515,503,-3515</points>
<connection>
<GID>1236</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>478,-3397,508,-3397</points>
<connection>
<GID>1158</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>478,-3605,506,-3605</points>
<connection>
<GID>1210</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>478,-3683,507,-3683</points>
<connection>
<GID>1288</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>478,-3773,510,-3773</points>
<connection>
<GID>1262</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>478,-3964.5,501,-3964.5</points>
<connection>
<GID>1411</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>478,-4132.5,505,-4132.5</points>
<connection>
<GID>1463</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>478,-4054.5,504,-4054.5</points>
<connection>
<GID>1385</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>478,-4222.5,508,-4222.5</points>
<connection>
<GID>1437</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>478,-4340.5,503,-4340.5</points>
<connection>
<GID>1306</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>478,-4430.5,506,-4430.5</points>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>478,-4508.5,507,-4508.5</points>
<connection>
<GID>1358</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>478,-4598.5,510,-4598.5</points>
<connection>
<GID>1332</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>478,-4889,498.5,-4889</points>
<connection>
<GID>1620</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>478,-5147,505.5,-5147</points>
<connection>
<GID>1646</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>478,-5265,500.5,-5265</points>
<connection>
<GID>1515</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>478,-5355,503.5,-5355</points>
<connection>
<GID>1698</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>478,-4979,501.5,-4979</points>
<connection>
<GID>1594</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>478,-5057,502.5,-5057</points>
<connection>
<GID>1672</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>478,-5433,504.5,-5433</points>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>478,-5523,507.5,-5523</points>
<connection>
<GID>1541</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>478,-5928.5,502,-5928.5</points>
<connection>
<GID>1881</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>478,-5850.5,501,-5850.5</points>
<connection>
<GID>1803</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>478,-5760.5,498,-5760.5</points>
<connection>
<GID>1829</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>478,-6226.5,503,-6226.5</points>
<connection>
<GID>1907</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>478,-6136.5,500,-6136.5</points>
<connection>
<GID>1724</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>478,-6018.5,505,-6018.5</points>
<connection>
<GID>1855</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>478,-6394.5,507,-6394.5</points>
<connection>
<GID>1750</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>478,-6304.5,504,-6304.5</points>
<connection>
<GID>1776</GID>
<name>IN_0</name></connection>
<intersection>478 0</intersection></hsegment></shape></wire>
<wire>
<ID>1472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>562,-6440,562,376.5</points>
<connection>
<GID>2113</GID>
<name>OUT_0</name></connection>
<intersection>-6394.5 62</intersection>
<intersection>-6304.5 63</intersection>
<intersection>-6226.5 61</intersection>
<intersection>-6136.5 60</intersection>
<intersection>-6018.5 59</intersection>
<intersection>-5928.5 58</intersection>
<intersection>-5850.5 57</intersection>
<intersection>-5760.5 56</intersection>
<intersection>-5523 55</intersection>
<intersection>-5433 54</intersection>
<intersection>-5355 53</intersection>
<intersection>-5265 52</intersection>
<intersection>-5147 51</intersection>
<intersection>-5057 50</intersection>
<intersection>-4979 49</intersection>
<intersection>-4889 48</intersection>
<intersection>-4598.5 47</intersection>
<intersection>-4508.5 44</intersection>
<intersection>-4430.5 45</intersection>
<intersection>-4340.5 46</intersection>
<intersection>-4222.5 43</intersection>
<intersection>-4132.5 42</intersection>
<intersection>-4054.5 41</intersection>
<intersection>-3964.5 40</intersection>
<intersection>-3773 38</intersection>
<intersection>-3683 39</intersection>
<intersection>-3605 37</intersection>
<intersection>-3515 36</intersection>
<intersection>-3397 35</intersection>
<intersection>-3307 34</intersection>
<intersection>-3229 33</intersection>
<intersection>-3139 32</intersection>
<intersection>-2879 31</intersection>
<intersection>-2789 30</intersection>
<intersection>-2711 29</intersection>
<intersection>-2621 28</intersection>
<intersection>-2413 27</intersection>
<intersection>-2335 26</intersection>
<intersection>-2245 25</intersection>
<intersection>-2007.5 24</intersection>
<intersection>-1917.5 23</intersection>
<intersection>-1839.5 22</intersection>
<intersection>-1749.5 21</intersection>
<intersection>-1631.5 20</intersection>
<intersection>-1541.5 19</intersection>
<intersection>-1463.5 18</intersection>
<intersection>-1373.5 17</intersection>
<intersection>-1083 16</intersection>
<intersection>-993 15</intersection>
<intersection>-915 14</intersection>
<intersection>-825 13</intersection>
<intersection>-707 12</intersection>
<intersection>-617 11</intersection>
<intersection>-539 10</intersection>
<intersection>-449 9</intersection>
<intersection>-257.5 8</intersection>
<intersection>-167.5 7</intersection>
<intersection>-89.5 6</intersection>
<intersection>0.5 4</intersection>
<intersection>118.5 5</intersection>
<intersection>208.5 3</intersection>
<intersection>286.5 2</intersection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562,376.5,576.5,376.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>562,286.5,579.5,286.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>562,208.5,580.5,208.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>562,0.5,578.5,0.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>562,118.5,583.5,118.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>562,-89.5,581.5,-89.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>562,-167.5,582.5,-167.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>562,-257.5,585.5,-257.5</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>562,-449,576.5,-449</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>562,-539,579.5,-539</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>562,-617,580.5,-617</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>562,-707,583.5,-707</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>562,-825,578.5,-825</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>562,-915,581.5,-915</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>562,-993,582.5,-993</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>562,-1083,585.5,-1083</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>562,-1373.5,574,-1373.5</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>562,-1463.5,577,-1463.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>562,-1541.5,578,-1541.5</points>
<connection>
<GID>839</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>562,-1631.5,581,-1631.5</points>
<connection>
<GID>813</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>562,-1749.5,576,-1749.5</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>562,-1839.5,579,-1839.5</points>
<connection>
<GID>865</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>562,-1917.5,580,-1917.5</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>562,-2007.5,583,-2007.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>562,-2245,573.5,-2245</points>
<connection>
<GID>996</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>562,-2335,576.5,-2335</points>
<connection>
<GID>970</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>562,-2413,577.5,-2413</points>
<connection>
<GID>1048</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>562,-2621,575.5,-2621</points>
<connection>
<GID>891</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>562,-2711,578.5,-2711</points>
<connection>
<GID>1074</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>562,-2789,579.5,-2789</points>
<connection>
<GID>943</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>562,-2879,582.5,-2879</points>
<connection>
<GID>917</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>562,-3139,574.5,-3139</points>
<connection>
<GID>1135</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>562,-3229,577.5,-3229</points>
<connection>
<GID>1109</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>562,-3307,578.5,-3307</points>
<connection>
<GID>1187</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>562,-3397,581.5,-3397</points>
<connection>
<GID>1161</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>562,-3515,576.5,-3515</points>
<connection>
<GID>1239</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>562,-3605,579.5,-3605</points>
<connection>
<GID>1213</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>562,-3773,583.5,-3773</points>
<connection>
<GID>1265</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>562,-3683,580.5,-3683</points>
<connection>
<GID>1291</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>562,-3964.5,574.5,-3964.5</points>
<connection>
<GID>1414</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>562,-4054.5,577.5,-4054.5</points>
<connection>
<GID>1388</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>562,-4132.5,578.5,-4132.5</points>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>562,-4222.5,581.5,-4222.5</points>
<connection>
<GID>1440</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>562,-4508.5,580.5,-4508.5</points>
<connection>
<GID>1361</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>562,-4430.5,579.5,-4430.5</points>
<connection>
<GID>1492</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>562,-4340.5,576.5,-4340.5</points>
<connection>
<GID>1309</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>562,-4598.5,583.5,-4598.5</points>
<connection>
<GID>1335</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>562,-4889,572,-4889</points>
<connection>
<GID>1623</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>562,-4979,575,-4979</points>
<connection>
<GID>1597</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>562,-5057,576,-5057</points>
<connection>
<GID>1675</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>562,-5147,579,-5147</points>
<connection>
<GID>1649</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>562,-5265,574,-5265</points>
<connection>
<GID>1518</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>562,-5355,577,-5355</points>
<connection>
<GID>1701</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>562,-5433,578,-5433</points>
<connection>
<GID>1570</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>562,-5523,581,-5523</points>
<connection>
<GID>1544</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>562,-5760.5,571.5,-5760.5</points>
<connection>
<GID>1832</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>562,-5850.5,574.5,-5850.5</points>
<connection>
<GID>1806</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>562,-5928.5,575.5,-5928.5</points>
<connection>
<GID>1884</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>562,-6018.5,578.5,-6018.5</points>
<connection>
<GID>1858</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>562,-6136.5,573.5,-6136.5</points>
<connection>
<GID>1727</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>562,-6226.5,576.5,-6226.5</points>
<connection>
<GID>1910</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>562,-6394.5,580.5,-6394.5</points>
<connection>
<GID>1753</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>562,-6304.5,577.5,-6304.5</points>
<connection>
<GID>1779</GID>
<name>IN_0</name></connection>
<intersection>562 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,181.954,1224,-423.046</PageViewport></page 2>
<page 3>
<PageViewport>0,181.954,1224,-423.046</PageViewport></page 3>
<page 4>
<PageViewport>0,181.954,1224,-423.046</PageViewport></page 4>
<page 5>
<PageViewport>0,181.954,1224,-423.046</PageViewport></page 5>
<page 6>
<PageViewport>74.986,-19.9309,211.487,-87.4007</PageViewport>
<gate>
<ID>51</ID>
<type>HA_JUNC_2</type>
<position>86,-43</position>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate></page 6>
<page 7>
<PageViewport>108.001,-5.85821,184.783,-43.8103</PageViewport>
<gate>
<ID>68</ID>
<type>BE_DECODER_3x8</type>
<position>123.5,-21</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate></page 7>
<page 8>
<PageViewport>67.8032,8.24731,391.365,-151.683</PageViewport>
<gate>
<ID>1958</ID>
<type>AA_TOGGLE</type>
<position>85,-42.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate></page 8>
<page 9>
<PageViewport>-141.018,810.696,1082.98,205.696</PageViewport>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>129,-26.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AE_DFF_LOW</type>
<position>45,-20</position>
<output>
<ID>OUT_0</ID>132 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>202</ID>
<type>BA_TRI_STATE</type>
<position>69.5,-26.5</position>
<input>
<ID>ENABLE_0</ID>131 </input>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_AND2</type>
<position>55,-26.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_DFF_LOW</type>
<position>118.5,-20</position>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>205</ID>
<type>BA_TRI_STATE</type>
<position>143,-26.5</position>
<input>
<ID>ENABLE_0</ID>133 </input>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND2</type>
<position>287,-28.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_DFF_LOW</type>
<position>203,-20</position>
<output>
<ID>OUT_0</ID>137 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>208</ID>
<type>BA_TRI_STATE</type>
<position>227.5,-28.5</position>
<input>
<ID>ENABLE_0</ID>136 </input>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND2</type>
<position>213,-28.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_DFF_LOW</type>
<position>277.5,-20</position>
<output>
<ID>OUT_0</ID>139 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>211</ID>
<type>BA_TRI_STATE</type>
<position>301,-28.5</position>
<input>
<ID>ENABLE_0</ID>138 </input>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_AND2</type>
<position>452,-30</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_DFF_LOW</type>
<position>368,-20</position>
<output>
<ID>OUT_0</ID>142 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>214</ID>
<type>BA_TRI_STATE</type>
<position>392.5,-30</position>
<input>
<ID>ENABLE_0</ID>141 </input>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>378,-30</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_DFF_LOW</type>
<position>441.5,-20</position>
<output>
<ID>OUT_0</ID>144 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>217</ID>
<type>BA_TRI_STATE</type>
<position>466,-30</position>
<input>
<ID>ENABLE_0</ID>143 </input>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>610,-32</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_DFF_LOW</type>
<position>526,-20</position>
<output>
<ID>OUT_0</ID>146 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>220</ID>
<type>BA_TRI_STATE</type>
<position>550.5,-32</position>
<input>
<ID>ENABLE_0</ID>145 </input>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>536,-32</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AE_DFF_LOW</type>
<position>599.5,-20</position>
<output>
<ID>OUT_0</ID>148 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>223</ID>
<type>BA_TRI_STATE</type>
<position>624,-32</position>
<input>
<ID>ENABLE_0</ID>147 </input>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>13.5,-21</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>BA_TRI_STATE</type>
<position>-8,-40</position>
<input>
<ID>ENABLE_0</ID>90 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-38,-8,-20</points>
<connection>
<GID>151</GID>
<name>ENABLE_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-20,10.5,-20</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>33</ID>
<points>-5.5,-40,607,-40</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>52 38</intersection>
<intersection>126 43</intersection>
<intersection>210 42</intersection>
<intersection>284 45</intersection>
<intersection>375 47</intersection>
<intersection>449 49</intersection>
<intersection>533 51</intersection>
<intersection>607 53</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>52,-40,52,-27.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>210,-40,210,-29.5</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>126,-40,126,-27.5</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>284,-40,284,-29.5</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>375,-40,375,-31</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>449,-40,449,-31</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>533,-40,533,-33</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>607,-40,607,-33</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>-40 33</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-26.5,67.5,-26.5</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<connection>
<GID>202</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-35,49,-18</points>
<intersection>-35 3</intersection>
<intersection>-25.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-25.5,52,-25.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-18,49,-18</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>49,-35,69.5,-35</points>
<intersection>49 0</intersection>
<intersection>69.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>69.5,-35,69.5,-29.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-35 3</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>132,-26.5,141,-26.5</points>
<connection>
<GID>205</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>200</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-36.5,122.5,-18</points>
<intersection>-36.5 3</intersection>
<intersection>-25.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-25.5,126,-25.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-18,122.5,-18</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>122.5,-36.5,143,-36.5</points>
<intersection>122.5 0</intersection>
<intersection>143 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>143,-36.5,143,-29.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-36.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-28.5,225.5,-28.5</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<connection>
<GID>208</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-37,207,-18</points>
<intersection>-37 3</intersection>
<intersection>-27.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-27.5,210,-27.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206,-18,207,-18</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,-37,227.5,-37</points>
<intersection>207 0</intersection>
<intersection>227.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>227.5,-37,227.5,-31.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-37 3</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>290,-28.5,299,-28.5</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<connection>
<GID>211</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-38.5,280.5,-18</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 3</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280.5,-27.5,284,-27.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280.5,-38.5,301,-38.5</points>
<intersection>280.5 0</intersection>
<intersection>301 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>301,-38.5,301,-31.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-38.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381,-30,390.5,-30</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-38.5,372,-18</points>
<intersection>-38.5 3</intersection>
<intersection>-29 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372,-29,375,-29</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>371,-18,372,-18</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>372,-38.5,392.5,-38.5</points>
<intersection>372 0</intersection>
<intersection>392.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>392.5,-38.5,392.5,-33</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-38.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>455,-30,464,-30</points>
<connection>
<GID>217</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>212</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,-38.5,445.5,-18</points>
<intersection>-38.5 3</intersection>
<intersection>-29 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,-29,449,-29</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444.5,-18,445.5,-18</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>445.5,-38.5,466,-38.5</points>
<intersection>445.5 0</intersection>
<intersection>466 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>466,-38.5,466,-33</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-38.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>539,-32,548.5,-32</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>220</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,-38,530,-18</points>
<intersection>-38 3</intersection>
<intersection>-31 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-31,533,-31</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,-18,530,-18</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>530,-38,550.5,-38</points>
<intersection>530 0</intersection>
<intersection>550.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>550.5,-38,550.5,-35</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-38 3</intersection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>613,-32,622,-32</points>
<connection>
<GID>223</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>218</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603.5,-38,603.5,-18</points>
<intersection>-38 3</intersection>
<intersection>-31 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>603.5,-31,607,-31</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>603.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>602.5,-18,603.5,-18</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>603.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>603.5,-38,624,-38</points>
<intersection>603.5 0</intersection>
<intersection>624 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>624,-38,624,-35</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-38 3</intersection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-21,596.5,-21</points>
<connection>
<GID>219</GID>
<name>clock</name></connection>
<connection>
<GID>213</GID>
<name>clock</name></connection>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<connection>
<GID>204</GID>
<name>clock</name></connection>
<connection>
<GID>201</GID>
<name>clock</name></connection>
<connection>
<GID>207</GID>
<name>clock</name></connection>
<connection>
<GID>210</GID>
<name>clock</name></connection>
<connection>
<GID>216</GID>
<name>clock</name></connection>
<connection>
<GID>222</GID>
<name>clock</name></connection></hsegment></shape></wire></page 9></circuit>