<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>105.173,494.287,243.029,426.148</PageViewport>
<gate>
<ID>2</ID>
<type>BA_TRI_STATE</type>
<position>492.5,537.5</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_TRI_STATE</type>
<position>462,536.5</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_TRI_STATE</type>
<position>431,536.5</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_TRI_STATE</type>
<position>400,537</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_TRI_STATE</type>
<position>369.5,536</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>BA_TRI_STATE</type>
<position>339,536.5</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_TRI_STATE</type>
<position>307,535.5</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>BA_TRI_STATE</type>
<position>276,536</position>
<input>
<ID>ENABLE_0</ID>2 </input>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>492.5,550.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O8</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>462,551</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O7</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>431,551</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O6</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>400,551</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O5</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>369.5,551</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O4</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>339,551</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O3</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>307,551</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O2</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>276,550.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O1</lparam></gate>
<gate>
<ID>31</ID>
<type>DE_TO</type>
<position>216,-937</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>35</ID>
<type>BA_TRI_STATE</type>
<position>241.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>BA_TRI_STATE</type>
<position>272.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>39</ID>
<type>BA_TRI_STATE</type>
<position>304.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>41</ID>
<type>BA_TRI_STATE</type>
<position>335.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>43</ID>
<type>BA_TRI_STATE</type>
<position>365.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>BA_TRI_STATE</type>
<position>396.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>BA_TRI_STATE</type>
<position>427.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_TRI_STATE</type>
<position>458.5,-911.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>225,-902</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>3130</ID>
<type>AA_AND2</type>
<position>263.5,-358</position>
<input>
<ID>IN_0</ID>2250 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3131</ID>
<type>BA_TRI_STATE</type>
<position>270.5,-358</position>
<input>
<ID>ENABLE_0</ID>2249 </input>
<input>
<ID>IN_0</ID>2250 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>241.5,-919</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>3132</ID>
<type>AE_DFF_LOW</type>
<position>251.5,-350.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2250 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3133</ID>
<type>HA_JUNC_2</type>
<position>247.5,-369</position>
<input>
<ID>N_in0</ID>4162 </input>
<input>
<ID>N_in1</ID>2414 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>272.5,-919</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>3134</ID>
<type>HA_JUNC_2</type>
<position>278.5,-369.5</position>
<input>
<ID>N_in0</ID>4164 </input>
<input>
<ID>N_in1</ID>2327 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3135</ID>
<type>HA_JUNC_2</type>
<position>310.5,-369.5</position>
<input>
<ID>N_in0</ID>4166 </input>
<input>
<ID>N_in1</ID>2328 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>304.5,-919.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>3136</ID>
<type>HA_JUNC_2</type>
<position>341.5,-368.5</position>
<input>
<ID>N_in0</ID>4168 </input>
<input>
<ID>N_in1</ID>2329 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3137</ID>
<type>HA_JUNC_2</type>
<position>371.5,-367.5</position>
<input>
<ID>N_in0</ID>4170 </input>
<input>
<ID>N_in1</ID>2330 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>335.5,-919.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>3138</ID>
<type>HA_JUNC_2</type>
<position>402.5,-367</position>
<input>
<ID>N_in0</ID>4172 </input>
<input>
<ID>N_in1</ID>2331 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3139</ID>
<type>HA_JUNC_2</type>
<position>464.5,-368</position>
<input>
<ID>N_in0</ID>4176 </input>
<input>
<ID>N_in1</ID>2333 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>61</ID>
<type>DE_TO</type>
<position>365.5,-919.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>3140</ID>
<type>HA_JUNC_2</type>
<position>433.5,-366</position>
<input>
<ID>N_in0</ID>4174 </input>
<input>
<ID>N_in1</ID>2332 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3141</ID>
<type>HA_JUNC_2</type>
<position>247.5,-227.5</position>
<input>
<ID>N_in0</ID>2414 </input>
<input>
<ID>N_in1</ID>4161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>63</ID>
<type>DE_TO</type>
<position>396.5,-920</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>3142</ID>
<type>HA_JUNC_2</type>
<position>278.5,-227.5</position>
<input>
<ID>N_in0</ID>2327 </input>
<input>
<ID>N_in1</ID>4160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3143</ID>
<type>HA_JUNC_2</type>
<position>310.5,-227.5</position>
<input>
<ID>N_in0</ID>2328 </input>
<input>
<ID>N_in1</ID>4158 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>427.5,-920.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>3144</ID>
<type>AA_AND2</type>
<position>295,-358</position>
<input>
<ID>IN_0</ID>2262 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3145</ID>
<type>BA_TRI_STATE</type>
<position>302,-358</position>
<input>
<ID>ENABLE_0</ID>2261 </input>
<input>
<ID>IN_0</ID>2262 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>458.5,-920.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>3146</ID>
<type>AE_DFF_LOW</type>
<position>282.5,-350.5</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2262 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3147</ID>
<type>AA_AND2</type>
<position>325.5,-358</position>
<input>
<ID>IN_0</ID>2264 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>136.5,449</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3148</ID>
<type>BA_TRI_STATE</type>
<position>332.5,-358</position>
<input>
<ID>ENABLE_0</ID>2263 </input>
<input>
<ID>IN_0</ID>2264 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>131,453</position>
<gparam>LABEL_TEXT i/p 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3149</ID>
<type>AE_DFF_LOW</type>
<position>313.5,-350.5</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2264 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3150</ID>
<type>AA_AND2</type>
<position>357,-358</position>
<input>
<ID>IN_0</ID>2266 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>136.5,445.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3151</ID>
<type>BA_TRI_STATE</type>
<position>364,-358</position>
<input>
<ID>ENABLE_0</ID>2265 </input>
<input>
<ID>IN_0</ID>2266 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>131,450</position>
<gparam>LABEL_TEXT i/p 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3152</ID>
<type>AE_DFF_LOW</type>
<position>344.5,-350.5</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2266 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3153</ID>
<type>AA_AND2</type>
<position>386.5,-358</position>
<input>
<ID>IN_0</ID>2268 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>136.5,452.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3154</ID>
<type>BA_TRI_STATE</type>
<position>393.5,-358</position>
<input>
<ID>ENABLE_0</ID>2267 </input>
<input>
<ID>IN_0</ID>2268 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>131,446</position>
<gparam>LABEL_TEXT i/p 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3155</ID>
<type>AE_DFF_LOW</type>
<position>374.5,-350.5</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2268 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3156</ID>
<type>AA_AND2</type>
<position>418,-358</position>
<input>
<ID>IN_0</ID>2270 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2269 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3157</ID>
<type>BA_TRI_STATE</type>
<position>425,-358</position>
<input>
<ID>ENABLE_0</ID>2269 </input>
<input>
<ID>IN_0</ID>2270 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3158</ID>
<type>AE_DFF_LOW</type>
<position>405.5,-350.5</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2270 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3159</ID>
<type>AA_AND2</type>
<position>448.5,-358</position>
<input>
<ID>IN_0</ID>2272 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2271 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3160</ID>
<type>BA_TRI_STATE</type>
<position>455.5,-358</position>
<input>
<ID>ENABLE_0</ID>2271 </input>
<input>
<ID>IN_0</ID>2272 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3161</ID>
<type>AE_DFF_LOW</type>
<position>436.5,-350.5</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2272 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3162</ID>
<type>AA_AND2</type>
<position>480,-358</position>
<input>
<ID>IN_0</ID>2274 </input>
<input>
<ID>IN_1</ID>2326 </input>
<output>
<ID>OUT</ID>2273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3163</ID>
<type>BA_TRI_STATE</type>
<position>487,-358</position>
<input>
<ID>ENABLE_0</ID>2273 </input>
<input>
<ID>IN_0</ID>2274 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3164</ID>
<type>AE_DFF_LOW</type>
<position>467.5,-350.5</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2274 </output>
<input>
<ID>clock</ID>2325 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3165</ID>
<type>AA_AND2</type>
<position>264,-341</position>
<input>
<ID>IN_0</ID>2276 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3166</ID>
<type>BA_TRI_STATE</type>
<position>271,-341</position>
<input>
<ID>ENABLE_0</ID>2275 </input>
<input>
<ID>IN_0</ID>2276 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3167</ID>
<type>AE_DFF_LOW</type>
<position>252,-333.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2276 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3168</ID>
<type>AA_AND2</type>
<position>295.5,-341</position>
<input>
<ID>IN_0</ID>2278 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3169</ID>
<type>BA_TRI_STATE</type>
<position>302.5,-341</position>
<input>
<ID>ENABLE_0</ID>2277 </input>
<input>
<ID>IN_0</ID>2278 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3170</ID>
<type>AE_DFF_LOW</type>
<position>283,-333.5</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2278 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3171</ID>
<type>AA_AND2</type>
<position>326,-341</position>
<input>
<ID>IN_0</ID>2280 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2279 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3172</ID>
<type>BA_TRI_STATE</type>
<position>333,-341</position>
<input>
<ID>ENABLE_0</ID>2279 </input>
<input>
<ID>IN_0</ID>2280 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3173</ID>
<type>AE_DFF_LOW</type>
<position>314,-333.5</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2280 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3174</ID>
<type>AA_AND2</type>
<position>357.5,-341</position>
<input>
<ID>IN_0</ID>2282 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3175</ID>
<type>BA_TRI_STATE</type>
<position>364.5,-341</position>
<input>
<ID>ENABLE_0</ID>2281 </input>
<input>
<ID>IN_0</ID>2282 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3176</ID>
<type>AE_DFF_LOW</type>
<position>345,-333.5</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2282 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3177</ID>
<type>AA_AND2</type>
<position>387,-341</position>
<input>
<ID>IN_0</ID>2284 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3178</ID>
<type>BA_TRI_STATE</type>
<position>394,-341</position>
<input>
<ID>ENABLE_0</ID>2283 </input>
<input>
<ID>IN_0</ID>2284 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3179</ID>
<type>AE_DFF_LOW</type>
<position>375,-333.5</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2284 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3180</ID>
<type>AA_AND2</type>
<position>418.5,-341</position>
<input>
<ID>IN_0</ID>2286 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2285 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3181</ID>
<type>BA_TRI_STATE</type>
<position>425.5,-341</position>
<input>
<ID>ENABLE_0</ID>2285 </input>
<input>
<ID>IN_0</ID>2286 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3182</ID>
<type>AE_DFF_LOW</type>
<position>406,-333.5</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2286 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3183</ID>
<type>AA_AND2</type>
<position>449,-341</position>
<input>
<ID>IN_0</ID>2288 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3184</ID>
<type>BA_TRI_STATE</type>
<position>456,-341</position>
<input>
<ID>ENABLE_0</ID>2287 </input>
<input>
<ID>IN_0</ID>2288 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3185</ID>
<type>AE_DFF_LOW</type>
<position>437,-333.5</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2288 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3186</ID>
<type>AA_AND2</type>
<position>480.5,-341</position>
<input>
<ID>IN_0</ID>2290 </input>
<input>
<ID>IN_1</ID>2324 </input>
<output>
<ID>OUT</ID>2289 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3187</ID>
<type>BA_TRI_STATE</type>
<position>487.5,-341</position>
<input>
<ID>ENABLE_0</ID>2289 </input>
<input>
<ID>IN_0</ID>2290 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3188</ID>
<type>AE_DFF_LOW</type>
<position>468,-333.5</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2290 </output>
<input>
<ID>clock</ID>2323 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3189</ID>
<type>AA_AND2</type>
<position>264.5,-325</position>
<input>
<ID>IN_0</ID>2292 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2291 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3190</ID>
<type>BA_TRI_STATE</type>
<position>271.5,-325</position>
<input>
<ID>ENABLE_0</ID>2291 </input>
<input>
<ID>IN_0</ID>2292 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3191</ID>
<type>AE_DFF_LOW</type>
<position>252.5,-317.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2292 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3192</ID>
<type>AA_AND2</type>
<position>296,-325</position>
<input>
<ID>IN_0</ID>2294 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2293 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3193</ID>
<type>BA_TRI_STATE</type>
<position>303,-325</position>
<input>
<ID>ENABLE_0</ID>2293 </input>
<input>
<ID>IN_0</ID>2294 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3194</ID>
<type>AE_DFF_LOW</type>
<position>283.5,-317.5</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2294 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3195</ID>
<type>AA_AND2</type>
<position>326.5,-325</position>
<input>
<ID>IN_0</ID>2296 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2295 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3196</ID>
<type>BA_TRI_STATE</type>
<position>333.5,-325</position>
<input>
<ID>ENABLE_0</ID>2295 </input>
<input>
<ID>IN_0</ID>2296 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3197</ID>
<type>AE_DFF_LOW</type>
<position>314.5,-317.5</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2296 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3198</ID>
<type>AA_AND2</type>
<position>358,-325</position>
<input>
<ID>IN_0</ID>2298 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2297 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3199</ID>
<type>BA_TRI_STATE</type>
<position>365,-325</position>
<input>
<ID>ENABLE_0</ID>2297 </input>
<input>
<ID>IN_0</ID>2298 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3200</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-317.5</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2298 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>122</ID>
<type>BE_DECODER_3x8</type>
<position>164.5,439</position>
<input>
<ID>ENABLE</ID>62 </input>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>63 </input>
<output>
<ID>OUT_0</ID>74 </output>
<output>
<ID>OUT_1</ID>73 </output>
<output>
<ID>OUT_2</ID>72 </output>
<output>
<ID>OUT_3</ID>70 </output>
<output>
<ID>OUT_4</ID>69 </output>
<output>
<ID>OUT_5</ID>68 </output>
<output>
<ID>OUT_6</ID>67 </output>
<output>
<ID>OUT_7</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>3201</ID>
<type>AA_AND2</type>
<position>387.5,-325</position>
<input>
<ID>IN_0</ID>2300 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2299 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3202</ID>
<type>BA_TRI_STATE</type>
<position>394.5,-325</position>
<input>
<ID>ENABLE_0</ID>2299 </input>
<input>
<ID>IN_0</ID>2300 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>154.5,442.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3203</ID>
<type>AE_DFF_LOW</type>
<position>375.5,-317.5</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2300 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3204</ID>
<type>AA_AND2</type>
<position>419,-325</position>
<input>
<ID>IN_0</ID>2302 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2301 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>151.5,443</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3205</ID>
<type>BA_TRI_STATE</type>
<position>426,-325</position>
<input>
<ID>ENABLE_0</ID>2301 </input>
<input>
<ID>IN_0</ID>2302 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3206</ID>
<type>AE_DFF_LOW</type>
<position>406.5,-317.5</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2302 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_TOGGLE</type>
<position>136.5,440</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3207</ID>
<type>AA_AND2</type>
<position>449.5,-325</position>
<input>
<ID>IN_0</ID>2304 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2303 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3208</ID>
<type>BA_TRI_STATE</type>
<position>456.5,-325</position>
<input>
<ID>ENABLE_0</ID>2303 </input>
<input>
<ID>IN_0</ID>2304 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>136.5,436</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3209</ID>
<type>AE_DFF_LOW</type>
<position>437.5,-317.5</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2304 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3210</ID>
<type>AA_AND2</type>
<position>481,-325</position>
<input>
<ID>IN_0</ID>2306 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>136.5,432</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3211</ID>
<type>BA_TRI_STATE</type>
<position>488,-325</position>
<input>
<ID>ENABLE_0</ID>2305 </input>
<input>
<ID>IN_0</ID>2306 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>131,440.5</position>
<gparam>LABEL_TEXT i/p 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3212</ID>
<type>AE_DFF_LOW</type>
<position>468.5,-317.5</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2306 </output>
<input>
<ID>clock</ID>2259 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>131,436.5</position>
<gparam>LABEL_TEXT i/p 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3213</ID>
<type>AA_AND2</type>
<position>265,-309.5</position>
<input>
<ID>IN_0</ID>2308 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2307 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>131,432.5</position>
<gparam>LABEL_TEXT i/p 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3214</ID>
<type>BA_TRI_STATE</type>
<position>272,-309.5</position>
<input>
<ID>ENABLE_0</ID>2307 </input>
<input>
<ID>IN_0</ID>2308 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3215</ID>
<type>AE_DFF_LOW</type>
<position>253,-302</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2308 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3216</ID>
<type>AA_AND2</type>
<position>296.5,-309.5</position>
<input>
<ID>IN_0</ID>2310 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2309 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_TOGGLE</type>
<position>114,449.5</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3217</ID>
<type>BA_TRI_STATE</type>
<position>303.5,-309.5</position>
<input>
<ID>ENABLE_0</ID>2309 </input>
<input>
<ID>IN_0</ID>2310 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>114,433.5</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3218</ID>
<type>AE_DFF_LOW</type>
<position>284,-302</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2310 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>113.5,441</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3219</ID>
<type>AA_AND2</type>
<position>327,-309.5</position>
<input>
<ID>IN_0</ID>2312 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2311 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>108,449.5</position>
<gparam>LABEL_TEXT Read</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3220</ID>
<type>BA_TRI_STATE</type>
<position>334,-309.5</position>
<input>
<ID>ENABLE_0</ID>2311 </input>
<input>
<ID>IN_0</ID>2312 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>108,441.5</position>
<gparam>LABEL_TEXT Write</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3221</ID>
<type>AE_DFF_LOW</type>
<position>315,-302</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2312 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>109.5,434</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3222</ID>
<type>AA_AND2</type>
<position>358.5,-309.5</position>
<input>
<ID>IN_0</ID>2314 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2313 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>121.5,449.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>3223</ID>
<type>BA_TRI_STATE</type>
<position>365.5,-309.5</position>
<input>
<ID>ENABLE_0</ID>2313 </input>
<input>
<ID>IN_0</ID>2314 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>121,441</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W</lparam></gate>
<gate>
<ID>3224</ID>
<type>AE_DFF_LOW</type>
<position>346,-302</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2314 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>120.5,433.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>3225</ID>
<type>AA_AND2</type>
<position>388,-309.5</position>
<input>
<ID>IN_0</ID>2316 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2315 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>124,461</position>
<input>
<ID>N_in3</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3226</ID>
<type>BA_TRI_STATE</type>
<position>395,-309.5</position>
<input>
<ID>ENABLE_0</ID>2315 </input>
<input>
<ID>IN_0</ID>2316 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>134.5,461</position>
<input>
<ID>N_in3</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3227</ID>
<type>AE_DFF_LOW</type>
<position>376,-302</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2316 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>144.5,461</position>
<input>
<ID>N_in3</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3228</ID>
<type>AA_AND2</type>
<position>419.5,-309.5</position>
<input>
<ID>IN_0</ID>2318 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2317 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>152,461</position>
<input>
<ID>N_in3</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3229</ID>
<type>BA_TRI_STATE</type>
<position>426.5,-309.5</position>
<input>
<ID>ENABLE_0</ID>2317 </input>
<input>
<ID>IN_0</ID>2318 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>163.5,461</position>
<input>
<ID>N_in3</ID>82 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3230</ID>
<type>AE_DFF_LOW</type>
<position>407,-302</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2318 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>182.5,461</position>
<input>
<ID>N_in3</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3231</ID>
<type>AA_AND2</type>
<position>450,-309.5</position>
<input>
<ID>IN_0</ID>2320 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2319 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>172.5,461</position>
<input>
<ID>N_in3</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3232</ID>
<type>BA_TRI_STATE</type>
<position>457,-309.5</position>
<input>
<ID>ENABLE_0</ID>2319 </input>
<input>
<ID>IN_0</ID>2320 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>190.5,461</position>
<input>
<ID>N_in3</ID>85 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3233</ID>
<type>AE_DFF_LOW</type>
<position>438,-302</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2320 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>108,461.5</position>
<gparam>LABEL_TEXT Data out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3234</ID>
<type>AA_AND2</type>
<position>481.5,-309.5</position>
<input>
<ID>IN_0</ID>2322 </input>
<input>
<ID>IN_1</ID>2258 </input>
<output>
<ID>OUT</ID>2321 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>124,468</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O1</lparam></gate>
<gate>
<ID>3235</ID>
<type>BA_TRI_STATE</type>
<position>488.5,-309.5</position>
<input>
<ID>ENABLE_0</ID>2321 </input>
<input>
<ID>IN_0</ID>2322 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>134.5,468</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O2</lparam></gate>
<gate>
<ID>3236</ID>
<type>AE_DFF_LOW</type>
<position>469,-302</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2322 </output>
<input>
<ID>clock</ID>2257 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>144.5,468</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O3</lparam></gate>
<gate>
<ID>3237</ID>
<type>HA_JUNC_2</type>
<position>341.5,-227.5</position>
<input>
<ID>N_in0</ID>2329 </input>
<input>
<ID>N_in1</ID>4156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>152,468</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O4</lparam></gate>
<gate>
<ID>3238</ID>
<type>HA_JUNC_2</type>
<position>372.5,-228</position>
<input>
<ID>N_in0</ID>2330 </input>
<input>
<ID>N_in1</ID>4154 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>163.5,468</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O5</lparam></gate>
<gate>
<ID>3239</ID>
<type>HA_JUNC_2</type>
<position>402.5,-227.5</position>
<input>
<ID>N_in0</ID>2331 </input>
<input>
<ID>N_in1</ID>4151 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>172.5,468</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O6</lparam></gate>
<gate>
<ID>3240</ID>
<type>HA_JUNC_2</type>
<position>433.5,-227.5</position>
<input>
<ID>N_in0</ID>2332 </input>
<input>
<ID>N_in1</ID>4149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>182.5,468</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O7</lparam></gate>
<gate>
<ID>3241</ID>
<type>HA_JUNC_2</type>
<position>464.5,-228</position>
<input>
<ID>N_in0</ID>2333 </input>
<input>
<ID>N_in1</ID>4147 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>190.5,468</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID O8</lparam></gate>
<gate>
<ID>3242</ID>
<type>HA_JUNC_2</type>
<position>276.5,-220.5</position>
<input>
<ID>N_in0</ID>2334 </input>
<input>
<ID>N_in1</ID>4159 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_TOGGLE</type>
<position>163,476</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3243</ID>
<type>HA_JUNC_2</type>
<position>276.5,-377.5</position>
<input>
<ID>N_in0</ID>4163 </input>
<input>
<ID>N_in1</ID>2334 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_TOGGLE</type>
<position>172.5,476</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3244</ID>
<type>HA_JUNC_2</type>
<position>339.5,-376.5</position>
<input>
<ID>N_in0</ID>4167 </input>
<input>
<ID>N_in1</ID>2336 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_TOGGLE</type>
<position>182,476</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3245</ID>
<type>HA_JUNC_2</type>
<position>370,-376</position>
<input>
<ID>N_in0</ID>4169 </input>
<input>
<ID>N_in1</ID>2337 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>190.5,476</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3246</ID>
<type>HA_JUNC_2</type>
<position>400.5,-376</position>
<input>
<ID>N_in0</ID>4171 </input>
<input>
<ID>N_in1</ID>2338 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>124,476</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3247</ID>
<type>HA_JUNC_2</type>
<position>431.5,-376</position>
<input>
<ID>N_in0</ID>4173 </input>
<input>
<ID>N_in1</ID>2339 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_TOGGLE</type>
<position>133.5,476</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3248</ID>
<type>HA_JUNC_2</type>
<position>462.5,-376.5</position>
<input>
<ID>N_in0</ID>4175 </input>
<input>
<ID>N_in1</ID>2340 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>144,476</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3249</ID>
<type>HA_JUNC_2</type>
<position>493,-376</position>
<input>
<ID>N_in0</ID>4177 </input>
<input>
<ID>N_in1</ID>2341 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>152,476</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3250</ID>
<type>HA_JUNC_2</type>
<position>493,-219</position>
<input>
<ID>N_in0</ID>2341 </input>
<input>
<ID>N_in1</ID>4146 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>108.5,477</position>
<gparam>LABEL_TEXT Data in</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3251</ID>
<type>HA_JUNC_2</type>
<position>462.5,-219.5</position>
<input>
<ID>N_in0</ID>2340 </input>
<input>
<ID>N_in1</ID>4148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>124,483</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>3252</ID>
<type>HA_JUNC_2</type>
<position>431.5,-220.5</position>
<input>
<ID>N_in0</ID>2339 </input>
<input>
<ID>N_in1</ID>4150 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>134,483</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>3253</ID>
<type>HA_JUNC_2</type>
<position>400.5,-220.5</position>
<input>
<ID>N_in0</ID>2338 </input>
<input>
<ID>N_in1</ID>4152 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>144,483</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>3254</ID>
<type>HA_JUNC_2</type>
<position>370,-220.5</position>
<input>
<ID>N_in0</ID>2337 </input>
<input>
<ID>N_in1</ID>4153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>176</ID>
<type>DE_TO</type>
<position>152,483</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>3255</ID>
<type>HA_JUNC_2</type>
<position>339.5,-220.5</position>
<input>
<ID>N_in0</ID>2336 </input>
<input>
<ID>N_in1</ID>4155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>177</ID>
<type>DE_TO</type>
<position>163,483</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>3256</ID>
<type>HA_JUNC_2</type>
<position>307.5,-220.5</position>
<input>
<ID>N_in0</ID>2335 </input>
<input>
<ID>N_in1</ID>4157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>178</ID>
<type>DE_TO</type>
<position>172.5,483</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>3257</ID>
<type>BE_DECODER_3x8</type>
<position>197.5,-293</position>
<input>
<ID>ENABLE</ID>70 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>2349 </output>
<output>
<ID>OUT_1</ID>2348 </output>
<output>
<ID>OUT_2</ID>2347 </output>
<output>
<ID>OUT_3</ID>2346 </output>
<output>
<ID>OUT_4</ID>2345 </output>
<output>
<ID>OUT_5</ID>2344 </output>
<output>
<ID>OUT_6</ID>2343 </output>
<output>
<ID>OUT_7</ID>2342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>182.5,483</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>3258</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-307.5</position>
<input>
<ID>ENABLE_0</ID>2346 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2258 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_TO</type>
<position>190.5,483</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>3259</ID>
<type>AA_AND2</type>
<position>233.5,-303</position>
<input>
<ID>IN_0</ID>2346 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2257 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3260</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-323.5</position>
<input>
<ID>ENABLE_0</ID>2347 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3261</ID>
<type>AA_AND2</type>
<position>233.5,-318.5</position>
<input>
<ID>IN_0</ID>2347 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3262</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-339.5</position>
<input>
<ID>ENABLE_0</ID>2348 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2324 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3263</ID>
<type>AA_AND2</type>
<position>233.5,-334.5</position>
<input>
<ID>IN_0</ID>2348 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3264</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-356.5</position>
<input>
<ID>ENABLE_0</ID>2349 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2326 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>226.5,536</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>3265</ID>
<type>AA_AND2</type>
<position>233.5,-351.5</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3266</ID>
<type>AA_AND2</type>
<position>264.5,-293</position>
<input>
<ID>IN_0</ID>2351 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>201,523</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>3267</ID>
<type>BA_TRI_STATE</type>
<position>271.5,-293</position>
<input>
<ID>ENABLE_0</ID>2350 </input>
<input>
<ID>IN_0</ID>2351 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3268</ID>
<type>AE_DFF_LOW</type>
<position>252.5,-285.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2351 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3269</ID>
<type>BA_TRI_STATE</type>
<position>240.5,-242.5</position>
<input>
<ID>ENABLE_0</ID>2342 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3270</ID>
<type>AA_AND2</type>
<position>234,-238</position>
<input>
<ID>IN_0</ID>2342 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2416 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3271</ID>
<type>BA_TRI_STATE</type>
<position>240.5,-258.5</position>
<input>
<ID>ENABLE_0</ID>2343 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3272</ID>
<type>AA_AND2</type>
<position>296,-293</position>
<input>
<ID>IN_0</ID>2353 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2352 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3273</ID>
<type>AA_AND2</type>
<position>233.5,-253.5</position>
<input>
<ID>IN_0</ID>2343 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2252 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3274</ID>
<type>BA_TRI_STATE</type>
<position>303,-293</position>
<input>
<ID>ENABLE_0</ID>2352 </input>
<input>
<ID>IN_0</ID>2353 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3275</ID>
<type>BA_TRI_STATE</type>
<position>240.5,-274.5</position>
<input>
<ID>ENABLE_0</ID>2344 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3276</ID>
<type>AE_DFF_LOW</type>
<position>283.5,-285.5</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2353 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3277</ID>
<type>AA_AND2</type>
<position>233.5,-269.5</position>
<input>
<ID>IN_0</ID>2344 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3278</ID>
<type>AA_AND2</type>
<position>326.5,-293</position>
<input>
<ID>IN_0</ID>2355 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3279</ID>
<type>BA_TRI_STATE</type>
<position>240.5,-291.5</position>
<input>
<ID>ENABLE_0</ID>2345 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2256 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3280</ID>
<type>BA_TRI_STATE</type>
<position>333.5,-293</position>
<input>
<ID>ENABLE_0</ID>2354 </input>
<input>
<ID>IN_0</ID>2355 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3281</ID>
<type>AA_AND2</type>
<position>233.5,-286.5</position>
<input>
<ID>IN_0</ID>2345 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3282</ID>
<type>AE_DFF_LOW</type>
<position>314.5,-285.5</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2355 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3283</ID>
<type>AA_AND2</type>
<position>358,-293</position>
<input>
<ID>IN_0</ID>2357 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2356 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3284</ID>
<type>BA_TRI_STATE</type>
<position>365,-293</position>
<input>
<ID>ENABLE_0</ID>2356 </input>
<input>
<ID>IN_0</ID>2357 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3285</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-285.5</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2357 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3286</ID>
<type>AA_AND2</type>
<position>387.5,-293</position>
<input>
<ID>IN_0</ID>2359 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2358 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3287</ID>
<type>BA_TRI_STATE</type>
<position>394.5,-293</position>
<input>
<ID>ENABLE_0</ID>2358 </input>
<input>
<ID>IN_0</ID>2359 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3288</ID>
<type>AE_DFF_LOW</type>
<position>375.5,-285.5</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2359 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3289</ID>
<type>AA_AND2</type>
<position>419,-293</position>
<input>
<ID>IN_0</ID>2361 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3290</ID>
<type>BA_TRI_STATE</type>
<position>426,-293</position>
<input>
<ID>ENABLE_0</ID>2360 </input>
<input>
<ID>IN_0</ID>2361 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3291</ID>
<type>AE_DFF_LOW</type>
<position>406.5,-285.5</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2361 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3292</ID>
<type>AA_AND2</type>
<position>449.5,-293</position>
<input>
<ID>IN_0</ID>2363 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2362 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3293</ID>
<type>BA_TRI_STATE</type>
<position>456.5,-293</position>
<input>
<ID>ENABLE_0</ID>2362 </input>
<input>
<ID>IN_0</ID>2363 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3294</ID>
<type>AE_DFF_LOW</type>
<position>437.5,-285.5</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2363 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3295</ID>
<type>AA_AND2</type>
<position>481,-293</position>
<input>
<ID>IN_0</ID>2365 </input>
<input>
<ID>IN_1</ID>2256 </input>
<output>
<ID>OUT</ID>2364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3296</ID>
<type>BA_TRI_STATE</type>
<position>488,-293</position>
<input>
<ID>ENABLE_0</ID>2364 </input>
<input>
<ID>IN_0</ID>2365 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3297</ID>
<type>AE_DFF_LOW</type>
<position>468.5,-285.5</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2365 </output>
<input>
<ID>clock</ID>2255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3298</ID>
<type>AA_AND2</type>
<position>265,-276</position>
<input>
<ID>IN_0</ID>2367 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2366 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3299</ID>
<type>BA_TRI_STATE</type>
<position>272,-276</position>
<input>
<ID>ENABLE_0</ID>2366 </input>
<input>
<ID>IN_0</ID>2367 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3300</ID>
<type>AE_DFF_LOW</type>
<position>253,-268.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2367 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3301</ID>
<type>AA_AND2</type>
<position>296.5,-276</position>
<input>
<ID>IN_0</ID>2369 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2368 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3302</ID>
<type>BA_TRI_STATE</type>
<position>303.5,-276</position>
<input>
<ID>ENABLE_0</ID>2368 </input>
<input>
<ID>IN_0</ID>2369 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3303</ID>
<type>AE_DFF_LOW</type>
<position>284,-268.5</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2369 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3304</ID>
<type>AA_AND2</type>
<position>327,-276</position>
<input>
<ID>IN_0</ID>2371 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3305</ID>
<type>BA_TRI_STATE</type>
<position>334,-276</position>
<input>
<ID>ENABLE_0</ID>2370 </input>
<input>
<ID>IN_0</ID>2371 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3306</ID>
<type>AE_DFF_LOW</type>
<position>315,-268.5</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2371 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3307</ID>
<type>AA_AND2</type>
<position>358.5,-276</position>
<input>
<ID>IN_0</ID>2373 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2372 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3308</ID>
<type>BA_TRI_STATE</type>
<position>365.5,-276</position>
<input>
<ID>ENABLE_0</ID>2372 </input>
<input>
<ID>IN_0</ID>2373 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3309</ID>
<type>AE_DFF_LOW</type>
<position>346,-268.5</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2373 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3310</ID>
<type>AA_AND2</type>
<position>388,-276</position>
<input>
<ID>IN_0</ID>2375 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3311</ID>
<type>BA_TRI_STATE</type>
<position>395,-276</position>
<input>
<ID>ENABLE_0</ID>2374 </input>
<input>
<ID>IN_0</ID>2375 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3312</ID>
<type>AE_DFF_LOW</type>
<position>376,-268.5</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2375 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3313</ID>
<type>AA_AND2</type>
<position>419.5,-276</position>
<input>
<ID>IN_0</ID>2377 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2376 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3314</ID>
<type>BA_TRI_STATE</type>
<position>426.5,-276</position>
<input>
<ID>ENABLE_0</ID>2376 </input>
<input>
<ID>IN_0</ID>2377 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3315</ID>
<type>AE_DFF_LOW</type>
<position>407,-268.5</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2377 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3316</ID>
<type>AA_AND2</type>
<position>450,-276</position>
<input>
<ID>IN_0</ID>2379 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2378 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3317</ID>
<type>BA_TRI_STATE</type>
<position>457,-276</position>
<input>
<ID>ENABLE_0</ID>2378 </input>
<input>
<ID>IN_0</ID>2379 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3318</ID>
<type>AE_DFF_LOW</type>
<position>438,-268.5</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2379 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3319</ID>
<type>AA_AND2</type>
<position>481.5,-276</position>
<input>
<ID>IN_0</ID>2381 </input>
<input>
<ID>IN_1</ID>2253 </input>
<output>
<ID>OUT</ID>2380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3320</ID>
<type>BA_TRI_STATE</type>
<position>488.5,-276</position>
<input>
<ID>ENABLE_0</ID>2380 </input>
<input>
<ID>IN_0</ID>2381 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3321</ID>
<type>AE_DFF_LOW</type>
<position>469,-268.5</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2381 </output>
<input>
<ID>clock</ID>2254 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3322</ID>
<type>AA_AND2</type>
<position>265.5,-260</position>
<input>
<ID>IN_0</ID>2383 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3323</ID>
<type>BA_TRI_STATE</type>
<position>272.5,-260</position>
<input>
<ID>ENABLE_0</ID>2382 </input>
<input>
<ID>IN_0</ID>2383 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3324</ID>
<type>AE_DFF_LOW</type>
<position>253.5,-252.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2383 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3325</ID>
<type>AA_AND2</type>
<position>297,-260</position>
<input>
<ID>IN_0</ID>2385 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2384 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3326</ID>
<type>BA_TRI_STATE</type>
<position>304,-260</position>
<input>
<ID>ENABLE_0</ID>2384 </input>
<input>
<ID>IN_0</ID>2385 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3327</ID>
<type>AE_DFF_LOW</type>
<position>284.5,-252.5</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2385 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3328</ID>
<type>AA_AND2</type>
<position>327.5,-260</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2386 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3329</ID>
<type>BA_TRI_STATE</type>
<position>334.5,-260</position>
<input>
<ID>ENABLE_0</ID>2386 </input>
<input>
<ID>IN_0</ID>2387 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3330</ID>
<type>AE_DFF_LOW</type>
<position>315.5,-252.5</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2387 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3331</ID>
<type>AA_AND2</type>
<position>359,-260</position>
<input>
<ID>IN_0</ID>2389 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2388 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3332</ID>
<type>BA_TRI_STATE</type>
<position>366,-260</position>
<input>
<ID>ENABLE_0</ID>2388 </input>
<input>
<ID>IN_0</ID>2389 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3333</ID>
<type>AE_DFF_LOW</type>
<position>346.5,-252.5</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2389 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3334</ID>
<type>AA_AND2</type>
<position>388.5,-260</position>
<input>
<ID>IN_0</ID>2391 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2390 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3335</ID>
<type>BA_TRI_STATE</type>
<position>395.5,-260</position>
<input>
<ID>ENABLE_0</ID>2390 </input>
<input>
<ID>IN_0</ID>2391 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3336</ID>
<type>AE_DFF_LOW</type>
<position>376.5,-252.5</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2391 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3337</ID>
<type>AA_AND2</type>
<position>420,-260</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3338</ID>
<type>BA_TRI_STATE</type>
<position>427,-260</position>
<input>
<ID>ENABLE_0</ID>2392 </input>
<input>
<ID>IN_0</ID>2393 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3339</ID>
<type>AE_DFF_LOW</type>
<position>407.5,-252.5</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2393 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3340</ID>
<type>AA_AND2</type>
<position>450.5,-260</position>
<input>
<ID>IN_0</ID>2395 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3341</ID>
<type>BA_TRI_STATE</type>
<position>457.5,-260</position>
<input>
<ID>ENABLE_0</ID>2394 </input>
<input>
<ID>IN_0</ID>2395 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3342</ID>
<type>AE_DFF_LOW</type>
<position>438.5,-252.5</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2395 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3343</ID>
<type>AA_AND2</type>
<position>482,-260</position>
<input>
<ID>IN_0</ID>2397 </input>
<input>
<ID>IN_1</ID>2251 </input>
<output>
<ID>OUT</ID>2396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3344</ID>
<type>BA_TRI_STATE</type>
<position>489,-260</position>
<input>
<ID>ENABLE_0</ID>2396 </input>
<input>
<ID>IN_0</ID>2397 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3345</ID>
<type>AE_DFF_LOW</type>
<position>469.5,-252.5</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2397 </output>
<input>
<ID>clock</ID>2252 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3346</ID>
<type>AA_AND2</type>
<position>266,-244.5</position>
<input>
<ID>IN_0</ID>2399 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2398 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3347</ID>
<type>BA_TRI_STATE</type>
<position>273,-244.5</position>
<input>
<ID>ENABLE_0</ID>2398 </input>
<input>
<ID>IN_0</ID>2399 </input>
<output>
<ID>OUT_0</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3348</ID>
<type>AE_DFF_LOW</type>
<position>254,-237</position>
<input>
<ID>IN_0</ID>2414 </input>
<output>
<ID>OUT_0</ID>2399 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3349</ID>
<type>AA_AND2</type>
<position>297.5,-244.5</position>
<input>
<ID>IN_0</ID>2401 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2400 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3350</ID>
<type>BA_TRI_STATE</type>
<position>304.5,-244.5</position>
<input>
<ID>ENABLE_0</ID>2400 </input>
<input>
<ID>IN_0</ID>2401 </input>
<output>
<ID>OUT_0</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3351</ID>
<type>AE_DFF_LOW</type>
<position>285,-237</position>
<input>
<ID>IN_0</ID>2327 </input>
<output>
<ID>OUT_0</ID>2401 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3352</ID>
<type>AA_AND2</type>
<position>328,-244.5</position>
<input>
<ID>IN_0</ID>2403 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2402 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3353</ID>
<type>BA_TRI_STATE</type>
<position>335,-244.5</position>
<input>
<ID>ENABLE_0</ID>2402 </input>
<input>
<ID>IN_0</ID>2403 </input>
<output>
<ID>OUT_0</ID>2336 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3354</ID>
<type>AE_DFF_LOW</type>
<position>316,-237</position>
<input>
<ID>IN_0</ID>2328 </input>
<output>
<ID>OUT_0</ID>2403 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3355</ID>
<type>AA_AND2</type>
<position>359.5,-244.5</position>
<input>
<ID>IN_0</ID>2405 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2404 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3356</ID>
<type>BA_TRI_STATE</type>
<position>366.5,-244.5</position>
<input>
<ID>ENABLE_0</ID>2404 </input>
<input>
<ID>IN_0</ID>2405 </input>
<output>
<ID>OUT_0</ID>2337 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3357</ID>
<type>AE_DFF_LOW</type>
<position>347,-237</position>
<input>
<ID>IN_0</ID>2329 </input>
<output>
<ID>OUT_0</ID>2405 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3358</ID>
<type>AA_AND2</type>
<position>389,-244.5</position>
<input>
<ID>IN_0</ID>2407 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2406 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3359</ID>
<type>BA_TRI_STATE</type>
<position>396,-244.5</position>
<input>
<ID>ENABLE_0</ID>2406 </input>
<input>
<ID>IN_0</ID>2407 </input>
<output>
<ID>OUT_0</ID>2338 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3360</ID>
<type>AE_DFF_LOW</type>
<position>377,-237</position>
<input>
<ID>IN_0</ID>2330 </input>
<output>
<ID>OUT_0</ID>2407 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3361</ID>
<type>AA_AND2</type>
<position>420.5,-244.5</position>
<input>
<ID>IN_0</ID>2409 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2408 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3362</ID>
<type>BA_TRI_STATE</type>
<position>427.5,-244.5</position>
<input>
<ID>ENABLE_0</ID>2408 </input>
<input>
<ID>IN_0</ID>2409 </input>
<output>
<ID>OUT_0</ID>2339 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3363</ID>
<type>AE_DFF_LOW</type>
<position>408,-237</position>
<input>
<ID>IN_0</ID>2331 </input>
<output>
<ID>OUT_0</ID>2409 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3364</ID>
<type>AA_AND2</type>
<position>451,-244.5</position>
<input>
<ID>IN_0</ID>2411 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3365</ID>
<type>BA_TRI_STATE</type>
<position>458,-244.5</position>
<input>
<ID>ENABLE_0</ID>2410 </input>
<input>
<ID>IN_0</ID>2411 </input>
<output>
<ID>OUT_0</ID>2340 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3366</ID>
<type>AE_DFF_LOW</type>
<position>439,-237</position>
<input>
<ID>IN_0</ID>2332 </input>
<output>
<ID>OUT_0</ID>2411 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3367</ID>
<type>AA_AND2</type>
<position>482.5,-244.5</position>
<input>
<ID>IN_0</ID>2413 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2412 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3368</ID>
<type>BA_TRI_STATE</type>
<position>489.5,-244.5</position>
<input>
<ID>ENABLE_0</ID>2412 </input>
<input>
<ID>IN_0</ID>2413 </input>
<output>
<ID>OUT_0</ID>2341 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3369</ID>
<type>AE_DFF_LOW</type>
<position>470,-237</position>
<input>
<ID>IN_0</ID>2333 </input>
<output>
<ID>OUT_0</ID>2413 </output>
<input>
<ID>clock</ID>2416 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3370</ID>
<type>AA_AND2</type>
<position>266.5,-531</position>
<input>
<ID>IN_0</ID>2417 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2417 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3371</ID>
<type>BA_TRI_STATE</type>
<position>273.5,-531</position>
<input>
<ID>ENABLE_0</ID>2417 </input>
<input>
<ID>IN_0</ID>2417 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3372</ID>
<type>AE_DFF_LOW</type>
<position>254.5,-523.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2417 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3373</ID>
<type>HA_JUNC_2</type>
<position>250.5,-542</position>
<input>
<ID>N_in0</ID>4178 </input>
<input>
<ID>N_in1</ID>2582 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3374</ID>
<type>HA_JUNC_2</type>
<position>281.5,-542.5</position>
<input>
<ID>N_in0</ID>4180 </input>
<input>
<ID>N_in1</ID>2495 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3375</ID>
<type>HA_JUNC_2</type>
<position>313.5,-542.5</position>
<input>
<ID>N_in0</ID>4182 </input>
<input>
<ID>N_in1</ID>2496 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3376</ID>
<type>HA_JUNC_2</type>
<position>344.5,-541.5</position>
<input>
<ID>N_in0</ID>4184 </input>
<input>
<ID>N_in1</ID>2497 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3377</ID>
<type>HA_JUNC_2</type>
<position>374.5,-540.5</position>
<input>
<ID>N_in0</ID>4186 </input>
<input>
<ID>N_in1</ID>2498 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3378</ID>
<type>HA_JUNC_2</type>
<position>405.5,-540</position>
<input>
<ID>N_in0</ID>4188 </input>
<input>
<ID>N_in1</ID>2499 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3379</ID>
<type>HA_JUNC_2</type>
<position>467.5,-541</position>
<input>
<ID>N_in0</ID>4192 </input>
<input>
<ID>N_in1</ID>2501 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3380</ID>
<type>HA_JUNC_2</type>
<position>436.5,-539</position>
<input>
<ID>N_in0</ID>4190 </input>
<input>
<ID>N_in1</ID>2500 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3381</ID>
<type>HA_JUNC_2</type>
<position>250.5,-400.5</position>
<input>
<ID>N_in0</ID>2582 </input>
<input>
<ID>N_in1</ID>4162 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3382</ID>
<type>HA_JUNC_2</type>
<position>281.5,-400.5</position>
<input>
<ID>N_in0</ID>2495 </input>
<input>
<ID>N_in1</ID>4164 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3383</ID>
<type>HA_JUNC_2</type>
<position>313.5,-400.5</position>
<input>
<ID>N_in0</ID>2496 </input>
<input>
<ID>N_in1</ID>4166 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3384</ID>
<type>AA_AND2</type>
<position>298,-531</position>
<input>
<ID>IN_0</ID>2430 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2429 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3385</ID>
<type>BA_TRI_STATE</type>
<position>305,-531</position>
<input>
<ID>ENABLE_0</ID>2429 </input>
<input>
<ID>IN_0</ID>2430 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3386</ID>
<type>AE_DFF_LOW</type>
<position>285.5,-523.5</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2430 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3387</ID>
<type>AA_AND2</type>
<position>328.5,-531</position>
<input>
<ID>IN_0</ID>2432 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3388</ID>
<type>BA_TRI_STATE</type>
<position>335.5,-531</position>
<input>
<ID>ENABLE_0</ID>2431 </input>
<input>
<ID>IN_0</ID>2432 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3389</ID>
<type>AE_DFF_LOW</type>
<position>316.5,-523.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2432 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3390</ID>
<type>AA_AND2</type>
<position>360,-531</position>
<input>
<ID>IN_0</ID>2434 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3391</ID>
<type>BA_TRI_STATE</type>
<position>367,-531</position>
<input>
<ID>ENABLE_0</ID>2433 </input>
<input>
<ID>IN_0</ID>2434 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3392</ID>
<type>AE_DFF_LOW</type>
<position>347.5,-523.5</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2434 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3393</ID>
<type>AA_AND2</type>
<position>389.5,-531</position>
<input>
<ID>IN_0</ID>2436 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3394</ID>
<type>BA_TRI_STATE</type>
<position>396.5,-531</position>
<input>
<ID>ENABLE_0</ID>2435 </input>
<input>
<ID>IN_0</ID>2436 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3395</ID>
<type>AE_DFF_LOW</type>
<position>377.5,-523.5</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2436 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3396</ID>
<type>AA_AND2</type>
<position>421,-531</position>
<input>
<ID>IN_0</ID>2438 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3397</ID>
<type>BA_TRI_STATE</type>
<position>428,-531</position>
<input>
<ID>ENABLE_0</ID>2437 </input>
<input>
<ID>IN_0</ID>2438 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3398</ID>
<type>AE_DFF_LOW</type>
<position>408.5,-523.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2438 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3399</ID>
<type>AA_AND2</type>
<position>451.5,-531</position>
<input>
<ID>IN_0</ID>2440 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3400</ID>
<type>BA_TRI_STATE</type>
<position>458.5,-531</position>
<input>
<ID>ENABLE_0</ID>2439 </input>
<input>
<ID>IN_0</ID>2440 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3401</ID>
<type>AE_DFF_LOW</type>
<position>439.5,-523.5</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2440 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3402</ID>
<type>AA_AND2</type>
<position>483,-531</position>
<input>
<ID>IN_0</ID>2442 </input>
<input>
<ID>IN_1</ID>2494 </input>
<output>
<ID>OUT</ID>2441 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3403</ID>
<type>BA_TRI_STATE</type>
<position>490,-531</position>
<input>
<ID>ENABLE_0</ID>2441 </input>
<input>
<ID>IN_0</ID>2442 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3404</ID>
<type>AE_DFF_LOW</type>
<position>470.5,-523.5</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2442 </output>
<input>
<ID>clock</ID>2493 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3405</ID>
<type>AA_AND2</type>
<position>267,-514</position>
<input>
<ID>IN_0</ID>2444 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2443 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3406</ID>
<type>BA_TRI_STATE</type>
<position>274,-514</position>
<input>
<ID>ENABLE_0</ID>2443 </input>
<input>
<ID>IN_0</ID>2444 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3407</ID>
<type>AE_DFF_LOW</type>
<position>255,-506.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2444 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3408</ID>
<type>AA_AND2</type>
<position>298.5,-514</position>
<input>
<ID>IN_0</ID>2446 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3409</ID>
<type>BA_TRI_STATE</type>
<position>305.5,-514</position>
<input>
<ID>ENABLE_0</ID>2445 </input>
<input>
<ID>IN_0</ID>2446 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3410</ID>
<type>AE_DFF_LOW</type>
<position>286,-506.5</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2446 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3411</ID>
<type>AA_AND2</type>
<position>329,-514</position>
<input>
<ID>IN_0</ID>2448 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2447 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3412</ID>
<type>BA_TRI_STATE</type>
<position>336,-514</position>
<input>
<ID>ENABLE_0</ID>2447 </input>
<input>
<ID>IN_0</ID>2448 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3413</ID>
<type>AE_DFF_LOW</type>
<position>317,-506.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2448 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3414</ID>
<type>AA_AND2</type>
<position>360.5,-514</position>
<input>
<ID>IN_0</ID>2450 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3415</ID>
<type>BA_TRI_STATE</type>
<position>367.5,-514</position>
<input>
<ID>ENABLE_0</ID>2449 </input>
<input>
<ID>IN_0</ID>2450 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3416</ID>
<type>AE_DFF_LOW</type>
<position>348,-506.5</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2450 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3417</ID>
<type>AA_AND2</type>
<position>390,-514</position>
<input>
<ID>IN_0</ID>2452 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3418</ID>
<type>BA_TRI_STATE</type>
<position>397,-514</position>
<input>
<ID>ENABLE_0</ID>2451 </input>
<input>
<ID>IN_0</ID>2452 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3419</ID>
<type>AE_DFF_LOW</type>
<position>378,-506.5</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2452 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3420</ID>
<type>AA_AND2</type>
<position>421.5,-514</position>
<input>
<ID>IN_0</ID>2454 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3421</ID>
<type>BA_TRI_STATE</type>
<position>428.5,-514</position>
<input>
<ID>ENABLE_0</ID>2453 </input>
<input>
<ID>IN_0</ID>2454 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3422</ID>
<type>AE_DFF_LOW</type>
<position>409,-506.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2454 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3423</ID>
<type>AA_AND2</type>
<position>452,-514</position>
<input>
<ID>IN_0</ID>2456 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2455 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3424</ID>
<type>BA_TRI_STATE</type>
<position>459,-514</position>
<input>
<ID>ENABLE_0</ID>2455 </input>
<input>
<ID>IN_0</ID>2456 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3425</ID>
<type>AE_DFF_LOW</type>
<position>440,-506.5</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2456 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3426</ID>
<type>AA_AND2</type>
<position>483.5,-514</position>
<input>
<ID>IN_0</ID>2458 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2457 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3427</ID>
<type>BA_TRI_STATE</type>
<position>490.5,-514</position>
<input>
<ID>ENABLE_0</ID>2457 </input>
<input>
<ID>IN_0</ID>2458 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3428</ID>
<type>AE_DFF_LOW</type>
<position>471,-506.5</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2458 </output>
<input>
<ID>clock</ID>2491 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3429</ID>
<type>AA_AND2</type>
<position>267.5,-498</position>
<input>
<ID>IN_0</ID>2460 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2459 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3430</ID>
<type>BA_TRI_STATE</type>
<position>274.5,-498</position>
<input>
<ID>ENABLE_0</ID>2459 </input>
<input>
<ID>IN_0</ID>2460 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3431</ID>
<type>AE_DFF_LOW</type>
<position>255.5,-490.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2460 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3432</ID>
<type>AA_AND2</type>
<position>299,-498</position>
<input>
<ID>IN_0</ID>2462 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2461 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3433</ID>
<type>BA_TRI_STATE</type>
<position>306,-498</position>
<input>
<ID>ENABLE_0</ID>2461 </input>
<input>
<ID>IN_0</ID>2462 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3434</ID>
<type>AE_DFF_LOW</type>
<position>286.5,-490.5</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2462 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3435</ID>
<type>AA_AND2</type>
<position>329.5,-498</position>
<input>
<ID>IN_0</ID>2464 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2463 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3436</ID>
<type>BA_TRI_STATE</type>
<position>336.5,-498</position>
<input>
<ID>ENABLE_0</ID>2463 </input>
<input>
<ID>IN_0</ID>2464 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3437</ID>
<type>AE_DFF_LOW</type>
<position>317.5,-490.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2464 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3438</ID>
<type>AA_AND2</type>
<position>361,-498</position>
<input>
<ID>IN_0</ID>2466 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2465 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3439</ID>
<type>BA_TRI_STATE</type>
<position>368,-498</position>
<input>
<ID>ENABLE_0</ID>2465 </input>
<input>
<ID>IN_0</ID>2466 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3440</ID>
<type>AE_DFF_LOW</type>
<position>348.5,-490.5</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2466 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3441</ID>
<type>AA_AND2</type>
<position>390.5,-498</position>
<input>
<ID>IN_0</ID>2468 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2467 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3442</ID>
<type>BA_TRI_STATE</type>
<position>397.5,-498</position>
<input>
<ID>ENABLE_0</ID>2467 </input>
<input>
<ID>IN_0</ID>2468 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3443</ID>
<type>AE_DFF_LOW</type>
<position>378.5,-490.5</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2468 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3444</ID>
<type>AA_AND2</type>
<position>422,-498</position>
<input>
<ID>IN_0</ID>2470 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2469 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3445</ID>
<type>BA_TRI_STATE</type>
<position>429,-498</position>
<input>
<ID>ENABLE_0</ID>2469 </input>
<input>
<ID>IN_0</ID>2470 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3446</ID>
<type>AE_DFF_LOW</type>
<position>409.5,-490.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2470 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3447</ID>
<type>AA_AND2</type>
<position>452.5,-498</position>
<input>
<ID>IN_0</ID>2472 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2471 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3448</ID>
<type>BA_TRI_STATE</type>
<position>459.5,-498</position>
<input>
<ID>ENABLE_0</ID>2471 </input>
<input>
<ID>IN_0</ID>2472 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3449</ID>
<type>AE_DFF_LOW</type>
<position>440.5,-490.5</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2472 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3450</ID>
<type>AA_AND2</type>
<position>484,-498</position>
<input>
<ID>IN_0</ID>2474 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2473 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3451</ID>
<type>BA_TRI_STATE</type>
<position>491,-498</position>
<input>
<ID>ENABLE_0</ID>2473 </input>
<input>
<ID>IN_0</ID>2474 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3452</ID>
<type>AE_DFF_LOW</type>
<position>471.5,-490.5</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2474 </output>
<input>
<ID>clock</ID>2427 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3453</ID>
<type>AA_AND2</type>
<position>268,-482.5</position>
<input>
<ID>IN_0</ID>2476 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2475 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3454</ID>
<type>BA_TRI_STATE</type>
<position>275,-482.5</position>
<input>
<ID>ENABLE_0</ID>2475 </input>
<input>
<ID>IN_0</ID>2476 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3455</ID>
<type>AE_DFF_LOW</type>
<position>256,-475</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2476 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3456</ID>
<type>AA_AND2</type>
<position>299.5,-482.5</position>
<input>
<ID>IN_0</ID>2478 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2477 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3457</ID>
<type>BA_TRI_STATE</type>
<position>306.5,-482.5</position>
<input>
<ID>ENABLE_0</ID>2477 </input>
<input>
<ID>IN_0</ID>2478 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3458</ID>
<type>AE_DFF_LOW</type>
<position>287,-475</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2478 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3459</ID>
<type>AA_AND2</type>
<position>330,-482.5</position>
<input>
<ID>IN_0</ID>2480 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3460</ID>
<type>BA_TRI_STATE</type>
<position>337,-482.5</position>
<input>
<ID>ENABLE_0</ID>2479 </input>
<input>
<ID>IN_0</ID>2480 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3461</ID>
<type>AE_DFF_LOW</type>
<position>318,-475</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2480 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3462</ID>
<type>AA_AND2</type>
<position>361.5,-482.5</position>
<input>
<ID>IN_0</ID>2482 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3463</ID>
<type>BA_TRI_STATE</type>
<position>368.5,-482.5</position>
<input>
<ID>ENABLE_0</ID>2481 </input>
<input>
<ID>IN_0</ID>2482 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3464</ID>
<type>AE_DFF_LOW</type>
<position>349,-475</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2482 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3465</ID>
<type>AA_AND2</type>
<position>391,-482.5</position>
<input>
<ID>IN_0</ID>2484 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3466</ID>
<type>BA_TRI_STATE</type>
<position>398,-482.5</position>
<input>
<ID>ENABLE_0</ID>2483 </input>
<input>
<ID>IN_0</ID>2484 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3467</ID>
<type>AE_DFF_LOW</type>
<position>379,-475</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2484 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3468</ID>
<type>AA_AND2</type>
<position>422.5,-482.5</position>
<input>
<ID>IN_0</ID>2486 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3469</ID>
<type>BA_TRI_STATE</type>
<position>429.5,-482.5</position>
<input>
<ID>ENABLE_0</ID>2485 </input>
<input>
<ID>IN_0</ID>2486 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3470</ID>
<type>AE_DFF_LOW</type>
<position>410,-475</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2486 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3471</ID>
<type>AA_AND2</type>
<position>453,-482.5</position>
<input>
<ID>IN_0</ID>2488 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3472</ID>
<type>BA_TRI_STATE</type>
<position>460,-482.5</position>
<input>
<ID>ENABLE_0</ID>2487 </input>
<input>
<ID>IN_0</ID>2488 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3473</ID>
<type>AE_DFF_LOW</type>
<position>441,-475</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2488 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3474</ID>
<type>AA_AND2</type>
<position>484.5,-482.5</position>
<input>
<ID>IN_0</ID>2490 </input>
<input>
<ID>IN_1</ID>2426 </input>
<output>
<ID>OUT</ID>2489 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3475</ID>
<type>BA_TRI_STATE</type>
<position>491.5,-482.5</position>
<input>
<ID>ENABLE_0</ID>2489 </input>
<input>
<ID>IN_0</ID>2490 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3476</ID>
<type>AE_DFF_LOW</type>
<position>472,-475</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2490 </output>
<input>
<ID>clock</ID>2425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3477</ID>
<type>HA_JUNC_2</type>
<position>344.5,-400.5</position>
<input>
<ID>N_in0</ID>2497 </input>
<input>
<ID>N_in1</ID>4168 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3478</ID>
<type>HA_JUNC_2</type>
<position>375.5,-401</position>
<input>
<ID>N_in0</ID>2498 </input>
<input>
<ID>N_in1</ID>4170 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3479</ID>
<type>HA_JUNC_2</type>
<position>405.5,-400.5</position>
<input>
<ID>N_in0</ID>2499 </input>
<input>
<ID>N_in1</ID>4172 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3480</ID>
<type>HA_JUNC_2</type>
<position>436.5,-400.5</position>
<input>
<ID>N_in0</ID>2500 </input>
<input>
<ID>N_in1</ID>4174 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3481</ID>
<type>HA_JUNC_2</type>
<position>467.5,-401</position>
<input>
<ID>N_in0</ID>2501 </input>
<input>
<ID>N_in1</ID>4176 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3482</ID>
<type>HA_JUNC_2</type>
<position>279.5,-393.5</position>
<input>
<ID>N_in0</ID>2502 </input>
<input>
<ID>N_in1</ID>4163 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3483</ID>
<type>HA_JUNC_2</type>
<position>279.5,-550.5</position>
<input>
<ID>N_in0</ID>4179 </input>
<input>
<ID>N_in1</ID>2502 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3484</ID>
<type>HA_JUNC_2</type>
<position>342.5,-549.5</position>
<input>
<ID>N_in0</ID>4183 </input>
<input>
<ID>N_in1</ID>2504 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3485</ID>
<type>HA_JUNC_2</type>
<position>373,-549</position>
<input>
<ID>N_in0</ID>4185 </input>
<input>
<ID>N_in1</ID>2505 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3486</ID>
<type>HA_JUNC_2</type>
<position>403.5,-549</position>
<input>
<ID>N_in0</ID>4187 </input>
<input>
<ID>N_in1</ID>2506 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3487</ID>
<type>HA_JUNC_2</type>
<position>434.5,-549</position>
<input>
<ID>N_in0</ID>4189 </input>
<input>
<ID>N_in1</ID>2507 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3488</ID>
<type>HA_JUNC_2</type>
<position>465.5,-549.5</position>
<input>
<ID>N_in0</ID>4191 </input>
<input>
<ID>N_in1</ID>2508 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3489</ID>
<type>HA_JUNC_2</type>
<position>496,-549</position>
<input>
<ID>N_in0</ID>4193 </input>
<input>
<ID>N_in1</ID>2509 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3490</ID>
<type>HA_JUNC_2</type>
<position>496,-392</position>
<input>
<ID>N_in0</ID>2509 </input>
<input>
<ID>N_in1</ID>4177 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3491</ID>
<type>HA_JUNC_2</type>
<position>465.5,-392.5</position>
<input>
<ID>N_in0</ID>2508 </input>
<input>
<ID>N_in1</ID>4175 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3492</ID>
<type>HA_JUNC_2</type>
<position>434.5,-393.5</position>
<input>
<ID>N_in0</ID>2507 </input>
<input>
<ID>N_in1</ID>4173 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3493</ID>
<type>HA_JUNC_2</type>
<position>403.5,-393.5</position>
<input>
<ID>N_in0</ID>2506 </input>
<input>
<ID>N_in1</ID>4171 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3494</ID>
<type>HA_JUNC_2</type>
<position>373,-393.5</position>
<input>
<ID>N_in0</ID>2505 </input>
<input>
<ID>N_in1</ID>4169 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3495</ID>
<type>HA_JUNC_2</type>
<position>342.5,-393.5</position>
<input>
<ID>N_in0</ID>2504 </input>
<input>
<ID>N_in1</ID>4167 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3496</ID>
<type>HA_JUNC_2</type>
<position>310.5,-393.5</position>
<input>
<ID>N_in0</ID>2503 </input>
<input>
<ID>N_in1</ID>4165 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3497</ID>
<type>BE_DECODER_3x8</type>
<position>200.5,-466</position>
<input>
<ID>ENABLE</ID>72 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>2517 </output>
<output>
<ID>OUT_1</ID>2516 </output>
<output>
<ID>OUT_2</ID>2515 </output>
<output>
<ID>OUT_3</ID>2514 </output>
<output>
<ID>OUT_4</ID>2513 </output>
<output>
<ID>OUT_5</ID>2512 </output>
<output>
<ID>OUT_6</ID>2511 </output>
<output>
<ID>OUT_7</ID>2510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>3498</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-480.5</position>
<input>
<ID>ENABLE_0</ID>2514 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2426 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3499</ID>
<type>AA_AND2</type>
<position>236.5,-476</position>
<input>
<ID>IN_0</ID>2514 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2425 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3500</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-496.5</position>
<input>
<ID>ENABLE_0</ID>2515 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3501</ID>
<type>AA_AND2</type>
<position>236.5,-491.5</position>
<input>
<ID>IN_0</ID>2515 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2427 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3502</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-512.5</position>
<input>
<ID>ENABLE_0</ID>2516 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3503</ID>
<type>AA_AND2</type>
<position>236.5,-507.5</position>
<input>
<ID>IN_0</ID>2516 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2491 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3504</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-529.5</position>
<input>
<ID>ENABLE_0</ID>2517 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3505</ID>
<type>AA_AND2</type>
<position>236.5,-524.5</position>
<input>
<ID>IN_0</ID>2517 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2493 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3506</ID>
<type>AA_AND2</type>
<position>267.5,-466</position>
<input>
<ID>IN_0</ID>2519 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3507</ID>
<type>BA_TRI_STATE</type>
<position>274.5,-466</position>
<input>
<ID>ENABLE_0</ID>2518 </input>
<input>
<ID>IN_0</ID>2519 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3508</ID>
<type>AE_DFF_LOW</type>
<position>255.5,-458.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2519 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3509</ID>
<type>BA_TRI_STATE</type>
<position>243.5,-415.5</position>
<input>
<ID>ENABLE_0</ID>2510 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2583 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3510</ID>
<type>AA_AND2</type>
<position>237,-411</position>
<input>
<ID>IN_0</ID>2510 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3511</ID>
<type>BA_TRI_STATE</type>
<position>243.5,-431.5</position>
<input>
<ID>ENABLE_0</ID>2511 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2419 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3512</ID>
<type>AA_AND2</type>
<position>299,-466</position>
<input>
<ID>IN_0</ID>2521 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3513</ID>
<type>AA_AND2</type>
<position>236.5,-426.5</position>
<input>
<ID>IN_0</ID>2511 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3514</ID>
<type>BA_TRI_STATE</type>
<position>306,-466</position>
<input>
<ID>ENABLE_0</ID>2520 </input>
<input>
<ID>IN_0</ID>2521 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3515</ID>
<type>BA_TRI_STATE</type>
<position>243.5,-447.5</position>
<input>
<ID>ENABLE_0</ID>2512 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2421 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3516</ID>
<type>AE_DFF_LOW</type>
<position>286.5,-458.5</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2521 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3517</ID>
<type>AA_AND2</type>
<position>236.5,-442.5</position>
<input>
<ID>IN_0</ID>2512 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2422 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3518</ID>
<type>AA_AND2</type>
<position>329.5,-466</position>
<input>
<ID>IN_0</ID>2523 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2522 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3519</ID>
<type>BA_TRI_STATE</type>
<position>243.5,-464.5</position>
<input>
<ID>ENABLE_0</ID>2513 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3520</ID>
<type>BA_TRI_STATE</type>
<position>336.5,-466</position>
<input>
<ID>ENABLE_0</ID>2522 </input>
<input>
<ID>IN_0</ID>2523 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3521</ID>
<type>AA_AND2</type>
<position>236.5,-459.5</position>
<input>
<ID>IN_0</ID>2513 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2423 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3522</ID>
<type>AE_DFF_LOW</type>
<position>317.5,-458.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2523 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3523</ID>
<type>AA_AND2</type>
<position>361,-466</position>
<input>
<ID>IN_0</ID>2525 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3524</ID>
<type>BA_TRI_STATE</type>
<position>368,-466</position>
<input>
<ID>ENABLE_0</ID>2524 </input>
<input>
<ID>IN_0</ID>2525 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3525</ID>
<type>AE_DFF_LOW</type>
<position>348.5,-458.5</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2525 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3526</ID>
<type>AA_AND2</type>
<position>390.5,-466</position>
<input>
<ID>IN_0</ID>2527 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2526 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3527</ID>
<type>BA_TRI_STATE</type>
<position>397.5,-466</position>
<input>
<ID>ENABLE_0</ID>2526 </input>
<input>
<ID>IN_0</ID>2527 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3528</ID>
<type>AE_DFF_LOW</type>
<position>378.5,-458.5</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2527 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3529</ID>
<type>AA_AND2</type>
<position>422,-466</position>
<input>
<ID>IN_0</ID>2529 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3530</ID>
<type>BA_TRI_STATE</type>
<position>429,-466</position>
<input>
<ID>ENABLE_0</ID>2528 </input>
<input>
<ID>IN_0</ID>2529 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3531</ID>
<type>AE_DFF_LOW</type>
<position>409.5,-458.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2529 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3532</ID>
<type>AA_AND2</type>
<position>452.5,-466</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2530 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3533</ID>
<type>BA_TRI_STATE</type>
<position>459.5,-466</position>
<input>
<ID>ENABLE_0</ID>2530 </input>
<input>
<ID>IN_0</ID>2531 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3534</ID>
<type>AE_DFF_LOW</type>
<position>440.5,-458.5</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2531 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3535</ID>
<type>AA_AND2</type>
<position>484,-466</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3536</ID>
<type>BA_TRI_STATE</type>
<position>491,-466</position>
<input>
<ID>ENABLE_0</ID>2532 </input>
<input>
<ID>IN_0</ID>2533 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3537</ID>
<type>AE_DFF_LOW</type>
<position>471.5,-458.5</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2533 </output>
<input>
<ID>clock</ID>2423 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3538</ID>
<type>AA_AND2</type>
<position>268,-449</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2534 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3539</ID>
<type>BA_TRI_STATE</type>
<position>275,-449</position>
<input>
<ID>ENABLE_0</ID>2534 </input>
<input>
<ID>IN_0</ID>2535 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3540</ID>
<type>AE_DFF_LOW</type>
<position>256,-441.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2535 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3541</ID>
<type>AA_AND2</type>
<position>299.5,-449</position>
<input>
<ID>IN_0</ID>2537 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2536 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3542</ID>
<type>BA_TRI_STATE</type>
<position>306.5,-449</position>
<input>
<ID>ENABLE_0</ID>2536 </input>
<input>
<ID>IN_0</ID>2537 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3543</ID>
<type>AE_DFF_LOW</type>
<position>287,-441.5</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2537 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3544</ID>
<type>AA_AND2</type>
<position>330,-449</position>
<input>
<ID>IN_0</ID>2539 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2538 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3545</ID>
<type>BA_TRI_STATE</type>
<position>337,-449</position>
<input>
<ID>ENABLE_0</ID>2538 </input>
<input>
<ID>IN_0</ID>2539 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3546</ID>
<type>AE_DFF_LOW</type>
<position>318,-441.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2539 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3547</ID>
<type>AA_AND2</type>
<position>361.5,-449</position>
<input>
<ID>IN_0</ID>2541 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2540 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3548</ID>
<type>BA_TRI_STATE</type>
<position>368.5,-449</position>
<input>
<ID>ENABLE_0</ID>2540 </input>
<input>
<ID>IN_0</ID>2541 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3549</ID>
<type>AE_DFF_LOW</type>
<position>349,-441.5</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2541 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3550</ID>
<type>AA_AND2</type>
<position>391,-449</position>
<input>
<ID>IN_0</ID>2543 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2542 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3551</ID>
<type>BA_TRI_STATE</type>
<position>398,-449</position>
<input>
<ID>ENABLE_0</ID>2542 </input>
<input>
<ID>IN_0</ID>2543 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3552</ID>
<type>AE_DFF_LOW</type>
<position>379,-441.5</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2543 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3553</ID>
<type>AA_AND2</type>
<position>422.5,-449</position>
<input>
<ID>IN_0</ID>2545 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2544 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3554</ID>
<type>BA_TRI_STATE</type>
<position>429.5,-449</position>
<input>
<ID>ENABLE_0</ID>2544 </input>
<input>
<ID>IN_0</ID>2545 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3555</ID>
<type>AE_DFF_LOW</type>
<position>410,-441.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2545 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3556</ID>
<type>AA_AND2</type>
<position>453,-449</position>
<input>
<ID>IN_0</ID>2547 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3557</ID>
<type>BA_TRI_STATE</type>
<position>460,-449</position>
<input>
<ID>ENABLE_0</ID>2546 </input>
<input>
<ID>IN_0</ID>2547 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3558</ID>
<type>AE_DFF_LOW</type>
<position>441,-441.5</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2547 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3559</ID>
<type>AA_AND2</type>
<position>484.5,-449</position>
<input>
<ID>IN_0</ID>2549 </input>
<input>
<ID>IN_1</ID>2421 </input>
<output>
<ID>OUT</ID>2548 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3560</ID>
<type>BA_TRI_STATE</type>
<position>491.5,-449</position>
<input>
<ID>ENABLE_0</ID>2548 </input>
<input>
<ID>IN_0</ID>2549 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3561</ID>
<type>AE_DFF_LOW</type>
<position>472,-441.5</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2549 </output>
<input>
<ID>clock</ID>2422 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3562</ID>
<type>AA_AND2</type>
<position>268.5,-433</position>
<input>
<ID>IN_0</ID>2551 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2550 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3563</ID>
<type>BA_TRI_STATE</type>
<position>275.5,-433</position>
<input>
<ID>ENABLE_0</ID>2550 </input>
<input>
<ID>IN_0</ID>2551 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3564</ID>
<type>AE_DFF_LOW</type>
<position>256.5,-425.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2551 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3565</ID>
<type>AA_AND2</type>
<position>300,-433</position>
<input>
<ID>IN_0</ID>2553 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2552 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3566</ID>
<type>BA_TRI_STATE</type>
<position>307,-433</position>
<input>
<ID>ENABLE_0</ID>2552 </input>
<input>
<ID>IN_0</ID>2553 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3567</ID>
<type>AE_DFF_LOW</type>
<position>287.5,-425.5</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2553 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3568</ID>
<type>AA_AND2</type>
<position>330.5,-433</position>
<input>
<ID>IN_0</ID>2555 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2554 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3569</ID>
<type>BA_TRI_STATE</type>
<position>337.5,-433</position>
<input>
<ID>ENABLE_0</ID>2554 </input>
<input>
<ID>IN_0</ID>2555 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3570</ID>
<type>AE_DFF_LOW</type>
<position>318.5,-425.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2555 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3571</ID>
<type>AA_AND2</type>
<position>362,-433</position>
<input>
<ID>IN_0</ID>2557 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3572</ID>
<type>BA_TRI_STATE</type>
<position>369,-433</position>
<input>
<ID>ENABLE_0</ID>2556 </input>
<input>
<ID>IN_0</ID>2557 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3573</ID>
<type>AE_DFF_LOW</type>
<position>349.5,-425.5</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2557 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3574</ID>
<type>AA_AND2</type>
<position>391.5,-433</position>
<input>
<ID>IN_0</ID>2559 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2558 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3575</ID>
<type>BA_TRI_STATE</type>
<position>398.5,-433</position>
<input>
<ID>ENABLE_0</ID>2558 </input>
<input>
<ID>IN_0</ID>2559 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3576</ID>
<type>AE_DFF_LOW</type>
<position>379.5,-425.5</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2559 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3577</ID>
<type>AA_AND2</type>
<position>423,-433</position>
<input>
<ID>IN_0</ID>2561 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2560 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3578</ID>
<type>BA_TRI_STATE</type>
<position>430,-433</position>
<input>
<ID>ENABLE_0</ID>2560 </input>
<input>
<ID>IN_0</ID>2561 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3579</ID>
<type>AE_DFF_LOW</type>
<position>410.5,-425.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2561 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3580</ID>
<type>AA_AND2</type>
<position>453.5,-433</position>
<input>
<ID>IN_0</ID>2563 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2562 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3581</ID>
<type>BA_TRI_STATE</type>
<position>460.5,-433</position>
<input>
<ID>ENABLE_0</ID>2562 </input>
<input>
<ID>IN_0</ID>2563 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3582</ID>
<type>AE_DFF_LOW</type>
<position>441.5,-425.5</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2563 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3583</ID>
<type>AA_AND2</type>
<position>485,-433</position>
<input>
<ID>IN_0</ID>2565 </input>
<input>
<ID>IN_1</ID>2419 </input>
<output>
<ID>OUT</ID>2564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3584</ID>
<type>BA_TRI_STATE</type>
<position>492,-433</position>
<input>
<ID>ENABLE_0</ID>2564 </input>
<input>
<ID>IN_0</ID>2565 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3585</ID>
<type>AE_DFF_LOW</type>
<position>472.5,-425.5</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2565 </output>
<input>
<ID>clock</ID>2420 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3586</ID>
<type>AA_AND2</type>
<position>269,-417.5</position>
<input>
<ID>IN_0</ID>2567 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2566 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3587</ID>
<type>BA_TRI_STATE</type>
<position>276,-417.5</position>
<input>
<ID>ENABLE_0</ID>2566 </input>
<input>
<ID>IN_0</ID>2567 </input>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3588</ID>
<type>AE_DFF_LOW</type>
<position>257,-410</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2567 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3589</ID>
<type>AA_AND2</type>
<position>300.5,-417.5</position>
<input>
<ID>IN_0</ID>2569 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2568 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3590</ID>
<type>BA_TRI_STATE</type>
<position>307.5,-417.5</position>
<input>
<ID>ENABLE_0</ID>2568 </input>
<input>
<ID>IN_0</ID>2569 </input>
<output>
<ID>OUT_0</ID>2503 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3591</ID>
<type>AE_DFF_LOW</type>
<position>288,-410</position>
<input>
<ID>IN_0</ID>2495 </input>
<output>
<ID>OUT_0</ID>2569 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3592</ID>
<type>AA_AND2</type>
<position>331,-417.5</position>
<input>
<ID>IN_0</ID>2571 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2570 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3593</ID>
<type>BA_TRI_STATE</type>
<position>338,-417.5</position>
<input>
<ID>ENABLE_0</ID>2570 </input>
<input>
<ID>IN_0</ID>2571 </input>
<output>
<ID>OUT_0</ID>2504 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3594</ID>
<type>AE_DFF_LOW</type>
<position>319,-410</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2571 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3595</ID>
<type>AA_AND2</type>
<position>362.5,-417.5</position>
<input>
<ID>IN_0</ID>2573 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2572 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3596</ID>
<type>BA_TRI_STATE</type>
<position>369.5,-417.5</position>
<input>
<ID>ENABLE_0</ID>2572 </input>
<input>
<ID>IN_0</ID>2573 </input>
<output>
<ID>OUT_0</ID>2505 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3597</ID>
<type>AE_DFF_LOW</type>
<position>350,-410</position>
<input>
<ID>IN_0</ID>2497 </input>
<output>
<ID>OUT_0</ID>2573 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3598</ID>
<type>AA_AND2</type>
<position>392,-417.5</position>
<input>
<ID>IN_0</ID>2575 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2574 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3599</ID>
<type>BA_TRI_STATE</type>
<position>399,-417.5</position>
<input>
<ID>ENABLE_0</ID>2574 </input>
<input>
<ID>IN_0</ID>2575 </input>
<output>
<ID>OUT_0</ID>2506 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3600</ID>
<type>AE_DFF_LOW</type>
<position>380,-410</position>
<input>
<ID>IN_0</ID>2498 </input>
<output>
<ID>OUT_0</ID>2575 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3601</ID>
<type>AA_AND2</type>
<position>423.5,-417.5</position>
<input>
<ID>IN_0</ID>2577 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2576 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3602</ID>
<type>BA_TRI_STATE</type>
<position>430.5,-417.5</position>
<input>
<ID>ENABLE_0</ID>2576 </input>
<input>
<ID>IN_0</ID>2577 </input>
<output>
<ID>OUT_0</ID>2507 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3603</ID>
<type>AE_DFF_LOW</type>
<position>411,-410</position>
<input>
<ID>IN_0</ID>2499 </input>
<output>
<ID>OUT_0</ID>2577 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3604</ID>
<type>AA_AND2</type>
<position>454,-417.5</position>
<input>
<ID>IN_0</ID>2579 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2578 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3605</ID>
<type>BA_TRI_STATE</type>
<position>461,-417.5</position>
<input>
<ID>ENABLE_0</ID>2578 </input>
<input>
<ID>IN_0</ID>2579 </input>
<output>
<ID>OUT_0</ID>2508 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3606</ID>
<type>AE_DFF_LOW</type>
<position>442,-410</position>
<input>
<ID>IN_0</ID>2500 </input>
<output>
<ID>OUT_0</ID>2579 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3607</ID>
<type>AA_AND2</type>
<position>485.5,-417.5</position>
<input>
<ID>IN_0</ID>2581 </input>
<input>
<ID>IN_1</ID>2583 </input>
<output>
<ID>OUT</ID>2580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3608</ID>
<type>BA_TRI_STATE</type>
<position>492.5,-417.5</position>
<input>
<ID>ENABLE_0</ID>2580 </input>
<input>
<ID>IN_0</ID>2581 </input>
<output>
<ID>OUT_0</ID>2509 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3609</ID>
<type>AE_DFF_LOW</type>
<position>473,-410</position>
<input>
<ID>IN_0</ID>2501 </input>
<output>
<ID>OUT_0</ID>2581 </output>
<input>
<ID>clock</ID>2584 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3850</ID>
<type>AA_AND2</type>
<position>262.5,-717</position>
<input>
<ID>IN_0</ID>2754 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2753 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3851</ID>
<type>BA_TRI_STATE</type>
<position>269.5,-717</position>
<input>
<ID>ENABLE_0</ID>2753 </input>
<input>
<ID>IN_0</ID>2754 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3852</ID>
<type>AE_DFF_LOW</type>
<position>250.5,-709.5</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2754 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3853</ID>
<type>HA_JUNC_2</type>
<position>246.5,-728</position>
<input>
<ID>N_in0</ID>4209 </input>
<input>
<ID>N_in1</ID>2918 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3854</ID>
<type>HA_JUNC_2</type>
<position>277.5,-728.5</position>
<input>
<ID>N_in0</ID>4208 </input>
<input>
<ID>N_in1</ID>2831 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3855</ID>
<type>HA_JUNC_2</type>
<position>309.5,-728.5</position>
<input>
<ID>N_in0</ID>4205 </input>
<input>
<ID>N_in1</ID>2832 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3856</ID>
<type>HA_JUNC_2</type>
<position>340.5,-727.5</position>
<input>
<ID>N_in0</ID>4204 </input>
<input>
<ID>N_in1</ID>2833 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3857</ID>
<type>HA_JUNC_2</type>
<position>370.5,-726.5</position>
<input>
<ID>N_in0</ID>4202 </input>
<input>
<ID>N_in1</ID>2834 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3858</ID>
<type>HA_JUNC_2</type>
<position>401.5,-726</position>
<input>
<ID>N_in0</ID>4200 </input>
<input>
<ID>N_in1</ID>2835 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3859</ID>
<type>HA_JUNC_2</type>
<position>463.5,-727</position>
<input>
<ID>N_in0</ID>4196 </input>
<input>
<ID>N_in1</ID>2837 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3860</ID>
<type>HA_JUNC_2</type>
<position>432.5,-725</position>
<input>
<ID>N_in0</ID>4198 </input>
<input>
<ID>N_in1</ID>2836 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3861</ID>
<type>HA_JUNC_2</type>
<position>246.5,-586.5</position>
<input>
<ID>N_in0</ID>2918 </input>
<input>
<ID>N_in1</ID>4178 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3862</ID>
<type>HA_JUNC_2</type>
<position>277.5,-586.5</position>
<input>
<ID>N_in0</ID>2831 </input>
<input>
<ID>N_in1</ID>4180 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3863</ID>
<type>HA_JUNC_2</type>
<position>309.5,-586.5</position>
<input>
<ID>N_in0</ID>2832 </input>
<input>
<ID>N_in1</ID>4182 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3864</ID>
<type>AA_AND2</type>
<position>294,-717</position>
<input>
<ID>IN_0</ID>2766 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2765 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3865</ID>
<type>BA_TRI_STATE</type>
<position>301,-717</position>
<input>
<ID>ENABLE_0</ID>2765 </input>
<input>
<ID>IN_0</ID>2766 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3866</ID>
<type>AE_DFF_LOW</type>
<position>281.5,-709.5</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2766 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3867</ID>
<type>AA_AND2</type>
<position>324.5,-717</position>
<input>
<ID>IN_0</ID>2768 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2767 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3868</ID>
<type>BA_TRI_STATE</type>
<position>331.5,-717</position>
<input>
<ID>ENABLE_0</ID>2767 </input>
<input>
<ID>IN_0</ID>2768 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3869</ID>
<type>AE_DFF_LOW</type>
<position>312.5,-709.5</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2768 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3870</ID>
<type>AA_AND2</type>
<position>356,-717</position>
<input>
<ID>IN_0</ID>2770 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2769 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3871</ID>
<type>BA_TRI_STATE</type>
<position>363,-717</position>
<input>
<ID>ENABLE_0</ID>2769 </input>
<input>
<ID>IN_0</ID>2770 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3872</ID>
<type>AE_DFF_LOW</type>
<position>343.5,-709.5</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2770 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3873</ID>
<type>AA_AND2</type>
<position>385.5,-717</position>
<input>
<ID>IN_0</ID>2772 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3874</ID>
<type>BA_TRI_STATE</type>
<position>392.5,-717</position>
<input>
<ID>ENABLE_0</ID>2771 </input>
<input>
<ID>IN_0</ID>2772 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3875</ID>
<type>AE_DFF_LOW</type>
<position>373.5,-709.5</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2772 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3876</ID>
<type>AA_AND2</type>
<position>417,-717</position>
<input>
<ID>IN_0</ID>2774 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2773 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3877</ID>
<type>BA_TRI_STATE</type>
<position>424,-717</position>
<input>
<ID>ENABLE_0</ID>2773 </input>
<input>
<ID>IN_0</ID>2774 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3878</ID>
<type>AE_DFF_LOW</type>
<position>404.5,-709.5</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2774 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3879</ID>
<type>AA_AND2</type>
<position>447.5,-717</position>
<input>
<ID>IN_0</ID>2776 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3880</ID>
<type>BA_TRI_STATE</type>
<position>454.5,-717</position>
<input>
<ID>ENABLE_0</ID>2775 </input>
<input>
<ID>IN_0</ID>2776 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3881</ID>
<type>AE_DFF_LOW</type>
<position>435.5,-709.5</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2776 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3882</ID>
<type>AA_AND2</type>
<position>479,-717</position>
<input>
<ID>IN_0</ID>2778 </input>
<input>
<ID>IN_1</ID>2830 </input>
<output>
<ID>OUT</ID>2777 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3883</ID>
<type>BA_TRI_STATE</type>
<position>486,-717</position>
<input>
<ID>ENABLE_0</ID>2777 </input>
<input>
<ID>IN_0</ID>2778 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3884</ID>
<type>AE_DFF_LOW</type>
<position>466.5,-709.5</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2778 </output>
<input>
<ID>clock</ID>2829 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3885</ID>
<type>AA_AND2</type>
<position>263,-700</position>
<input>
<ID>IN_0</ID>2780 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2779 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3886</ID>
<type>BA_TRI_STATE</type>
<position>270,-700</position>
<input>
<ID>ENABLE_0</ID>2779 </input>
<input>
<ID>IN_0</ID>2780 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3887</ID>
<type>AE_DFF_LOW</type>
<position>251,-692.5</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2780 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3888</ID>
<type>AA_AND2</type>
<position>294.5,-700</position>
<input>
<ID>IN_0</ID>2782 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3889</ID>
<type>BA_TRI_STATE</type>
<position>301.5,-700</position>
<input>
<ID>ENABLE_0</ID>2781 </input>
<input>
<ID>IN_0</ID>2782 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3890</ID>
<type>AE_DFF_LOW</type>
<position>282,-692.5</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2782 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3891</ID>
<type>AA_AND2</type>
<position>325,-700</position>
<input>
<ID>IN_0</ID>2784 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3892</ID>
<type>BA_TRI_STATE</type>
<position>332,-700</position>
<input>
<ID>ENABLE_0</ID>2783 </input>
<input>
<ID>IN_0</ID>2784 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3893</ID>
<type>AE_DFF_LOW</type>
<position>313,-692.5</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2784 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3894</ID>
<type>AA_AND2</type>
<position>356.5,-700</position>
<input>
<ID>IN_0</ID>2786 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2785 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3895</ID>
<type>BA_TRI_STATE</type>
<position>363.5,-700</position>
<input>
<ID>ENABLE_0</ID>2785 </input>
<input>
<ID>IN_0</ID>2786 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3896</ID>
<type>AE_DFF_LOW</type>
<position>344,-692.5</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2786 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3897</ID>
<type>AA_AND2</type>
<position>386,-700</position>
<input>
<ID>IN_0</ID>2788 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2787 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3898</ID>
<type>BA_TRI_STATE</type>
<position>393,-700</position>
<input>
<ID>ENABLE_0</ID>2787 </input>
<input>
<ID>IN_0</ID>2788 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3899</ID>
<type>AE_DFF_LOW</type>
<position>374,-692.5</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2788 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3900</ID>
<type>AA_AND2</type>
<position>417.5,-700</position>
<input>
<ID>IN_0</ID>2790 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2789 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3901</ID>
<type>BA_TRI_STATE</type>
<position>424.5,-700</position>
<input>
<ID>ENABLE_0</ID>2789 </input>
<input>
<ID>IN_0</ID>2790 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3902</ID>
<type>AE_DFF_LOW</type>
<position>405,-692.5</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2790 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3903</ID>
<type>AA_AND2</type>
<position>448,-700</position>
<input>
<ID>IN_0</ID>2792 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2791 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3904</ID>
<type>BA_TRI_STATE</type>
<position>455,-700</position>
<input>
<ID>ENABLE_0</ID>2791 </input>
<input>
<ID>IN_0</ID>2792 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3905</ID>
<type>AE_DFF_LOW</type>
<position>436,-692.5</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2792 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3906</ID>
<type>AA_AND2</type>
<position>479.5,-700</position>
<input>
<ID>IN_0</ID>2794 </input>
<input>
<ID>IN_1</ID>2828 </input>
<output>
<ID>OUT</ID>2793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3907</ID>
<type>BA_TRI_STATE</type>
<position>486.5,-700</position>
<input>
<ID>ENABLE_0</ID>2793 </input>
<input>
<ID>IN_0</ID>2794 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3908</ID>
<type>AE_DFF_LOW</type>
<position>467,-692.5</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2794 </output>
<input>
<ID>clock</ID>2827 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3909</ID>
<type>AA_AND2</type>
<position>263.5,-684</position>
<input>
<ID>IN_0</ID>2796 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2795 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3910</ID>
<type>BA_TRI_STATE</type>
<position>270.5,-684</position>
<input>
<ID>ENABLE_0</ID>2795 </input>
<input>
<ID>IN_0</ID>2796 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3911</ID>
<type>AE_DFF_LOW</type>
<position>251.5,-676.5</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2796 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3912</ID>
<type>AA_AND2</type>
<position>295,-684</position>
<input>
<ID>IN_0</ID>2798 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2797 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3913</ID>
<type>BA_TRI_STATE</type>
<position>302,-684</position>
<input>
<ID>ENABLE_0</ID>2797 </input>
<input>
<ID>IN_0</ID>2798 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3914</ID>
<type>AE_DFF_LOW</type>
<position>282.5,-676.5</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2798 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3915</ID>
<type>AA_AND2</type>
<position>325.5,-684</position>
<input>
<ID>IN_0</ID>2800 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2799 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3916</ID>
<type>BA_TRI_STATE</type>
<position>332.5,-684</position>
<input>
<ID>ENABLE_0</ID>2799 </input>
<input>
<ID>IN_0</ID>2800 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3917</ID>
<type>AE_DFF_LOW</type>
<position>313.5,-676.5</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2800 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3918</ID>
<type>AA_AND2</type>
<position>357,-684</position>
<input>
<ID>IN_0</ID>2802 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2801 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3919</ID>
<type>BA_TRI_STATE</type>
<position>364,-684</position>
<input>
<ID>ENABLE_0</ID>2801 </input>
<input>
<ID>IN_0</ID>2802 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3920</ID>
<type>AE_DFF_LOW</type>
<position>344.5,-676.5</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2802 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3921</ID>
<type>AA_AND2</type>
<position>386.5,-684</position>
<input>
<ID>IN_0</ID>2804 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2803 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3922</ID>
<type>BA_TRI_STATE</type>
<position>393.5,-684</position>
<input>
<ID>ENABLE_0</ID>2803 </input>
<input>
<ID>IN_0</ID>2804 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3923</ID>
<type>AE_DFF_LOW</type>
<position>374.5,-676.5</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2804 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3924</ID>
<type>AA_AND2</type>
<position>418,-684</position>
<input>
<ID>IN_0</ID>2806 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2805 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3925</ID>
<type>BA_TRI_STATE</type>
<position>425,-684</position>
<input>
<ID>ENABLE_0</ID>2805 </input>
<input>
<ID>IN_0</ID>2806 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3926</ID>
<type>AE_DFF_LOW</type>
<position>405.5,-676.5</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2806 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3927</ID>
<type>AA_AND2</type>
<position>448.5,-684</position>
<input>
<ID>IN_0</ID>2808 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2807 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3928</ID>
<type>BA_TRI_STATE</type>
<position>455.5,-684</position>
<input>
<ID>ENABLE_0</ID>2807 </input>
<input>
<ID>IN_0</ID>2808 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3929</ID>
<type>AE_DFF_LOW</type>
<position>436.5,-676.5</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2808 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3930</ID>
<type>AA_AND2</type>
<position>480,-684</position>
<input>
<ID>IN_0</ID>2810 </input>
<input>
<ID>IN_1</ID>2764 </input>
<output>
<ID>OUT</ID>2809 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3931</ID>
<type>BA_TRI_STATE</type>
<position>487,-684</position>
<input>
<ID>ENABLE_0</ID>2809 </input>
<input>
<ID>IN_0</ID>2810 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3932</ID>
<type>AE_DFF_LOW</type>
<position>467.5,-676.5</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2810 </output>
<input>
<ID>clock</ID>2763 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3933</ID>
<type>AA_AND2</type>
<position>264,-668.5</position>
<input>
<ID>IN_0</ID>2812 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2811 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3934</ID>
<type>BA_TRI_STATE</type>
<position>271,-668.5</position>
<input>
<ID>ENABLE_0</ID>2811 </input>
<input>
<ID>IN_0</ID>2812 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3935</ID>
<type>AE_DFF_LOW</type>
<position>252,-661</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2812 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3936</ID>
<type>AA_AND2</type>
<position>295.5,-668.5</position>
<input>
<ID>IN_0</ID>2814 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2813 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3937</ID>
<type>BA_TRI_STATE</type>
<position>302.5,-668.5</position>
<input>
<ID>ENABLE_0</ID>2813 </input>
<input>
<ID>IN_0</ID>2814 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3938</ID>
<type>AE_DFF_LOW</type>
<position>283,-661</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2814 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3939</ID>
<type>AA_AND2</type>
<position>326,-668.5</position>
<input>
<ID>IN_0</ID>2816 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2815 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3940</ID>
<type>BA_TRI_STATE</type>
<position>333,-668.5</position>
<input>
<ID>ENABLE_0</ID>2815 </input>
<input>
<ID>IN_0</ID>2816 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3941</ID>
<type>AE_DFF_LOW</type>
<position>314,-661</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2816 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3942</ID>
<type>AA_AND2</type>
<position>357.5,-668.5</position>
<input>
<ID>IN_0</ID>2818 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3943</ID>
<type>BA_TRI_STATE</type>
<position>364.5,-668.5</position>
<input>
<ID>ENABLE_0</ID>2817 </input>
<input>
<ID>IN_0</ID>2818 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3944</ID>
<type>AE_DFF_LOW</type>
<position>345,-661</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2818 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3945</ID>
<type>AA_AND2</type>
<position>387,-668.5</position>
<input>
<ID>IN_0</ID>2820 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3946</ID>
<type>BA_TRI_STATE</type>
<position>394,-668.5</position>
<input>
<ID>ENABLE_0</ID>2819 </input>
<input>
<ID>IN_0</ID>2820 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3947</ID>
<type>AE_DFF_LOW</type>
<position>375,-661</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2820 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3948</ID>
<type>AA_AND2</type>
<position>418.5,-668.5</position>
<input>
<ID>IN_0</ID>2822 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2821 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3949</ID>
<type>BA_TRI_STATE</type>
<position>425.5,-668.5</position>
<input>
<ID>ENABLE_0</ID>2821 </input>
<input>
<ID>IN_0</ID>2822 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3950</ID>
<type>AE_DFF_LOW</type>
<position>406,-661</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2822 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3951</ID>
<type>AA_AND2</type>
<position>449,-668.5</position>
<input>
<ID>IN_0</ID>2824 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2823 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3952</ID>
<type>BA_TRI_STATE</type>
<position>456,-668.5</position>
<input>
<ID>ENABLE_0</ID>2823 </input>
<input>
<ID>IN_0</ID>2824 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3953</ID>
<type>AE_DFF_LOW</type>
<position>437,-661</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2824 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3954</ID>
<type>AA_AND2</type>
<position>480.5,-668.5</position>
<input>
<ID>IN_0</ID>2826 </input>
<input>
<ID>IN_1</ID>2762 </input>
<output>
<ID>OUT</ID>2825 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3955</ID>
<type>BA_TRI_STATE</type>
<position>487.5,-668.5</position>
<input>
<ID>ENABLE_0</ID>2825 </input>
<input>
<ID>IN_0</ID>2826 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3956</ID>
<type>AE_DFF_LOW</type>
<position>468,-661</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2826 </output>
<input>
<ID>clock</ID>2761 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3957</ID>
<type>HA_JUNC_2</type>
<position>340.5,-586.5</position>
<input>
<ID>N_in0</ID>2833 </input>
<input>
<ID>N_in1</ID>4184 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3958</ID>
<type>HA_JUNC_2</type>
<position>371.5,-587</position>
<input>
<ID>N_in0</ID>2834 </input>
<input>
<ID>N_in1</ID>4186 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3959</ID>
<type>HA_JUNC_2</type>
<position>401.5,-586.5</position>
<input>
<ID>N_in0</ID>2835 </input>
<input>
<ID>N_in1</ID>4188 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3960</ID>
<type>HA_JUNC_2</type>
<position>432.5,-586.5</position>
<input>
<ID>N_in0</ID>2836 </input>
<input>
<ID>N_in1</ID>4190 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3961</ID>
<type>HA_JUNC_2</type>
<position>463.5,-587</position>
<input>
<ID>N_in0</ID>2837 </input>
<input>
<ID>N_in1</ID>4192 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3962</ID>
<type>HA_JUNC_2</type>
<position>275.5,-579.5</position>
<input>
<ID>N_in0</ID>2838 </input>
<input>
<ID>N_in1</ID>4179 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3963</ID>
<type>HA_JUNC_2</type>
<position>275.5,-736.5</position>
<input>
<ID>N_in0</ID>4207 </input>
<input>
<ID>N_in1</ID>2838 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3964</ID>
<type>HA_JUNC_2</type>
<position>338.5,-735.5</position>
<input>
<ID>N_in0</ID>4203 </input>
<input>
<ID>N_in1</ID>2840 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3965</ID>
<type>HA_JUNC_2</type>
<position>369,-735</position>
<input>
<ID>N_in0</ID>4201 </input>
<input>
<ID>N_in1</ID>2841 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3966</ID>
<type>HA_JUNC_2</type>
<position>399.5,-735</position>
<input>
<ID>N_in0</ID>4199 </input>
<input>
<ID>N_in1</ID>2842 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3967</ID>
<type>HA_JUNC_2</type>
<position>430.5,-735</position>
<input>
<ID>N_in0</ID>4197 </input>
<input>
<ID>N_in1</ID>2843 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3968</ID>
<type>HA_JUNC_2</type>
<position>461.5,-735.5</position>
<input>
<ID>N_in0</ID>4195 </input>
<input>
<ID>N_in1</ID>2844 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3969</ID>
<type>HA_JUNC_2</type>
<position>492,-735</position>
<input>
<ID>N_in0</ID>4194 </input>
<input>
<ID>N_in1</ID>2845 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3970</ID>
<type>HA_JUNC_2</type>
<position>492,-578</position>
<input>
<ID>N_in0</ID>2845 </input>
<input>
<ID>N_in1</ID>4193 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3971</ID>
<type>HA_JUNC_2</type>
<position>461.5,-578.5</position>
<input>
<ID>N_in0</ID>2844 </input>
<input>
<ID>N_in1</ID>4191 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3972</ID>
<type>HA_JUNC_2</type>
<position>430.5,-579.5</position>
<input>
<ID>N_in0</ID>2843 </input>
<input>
<ID>N_in1</ID>4189 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3973</ID>
<type>HA_JUNC_2</type>
<position>399.5,-579.5</position>
<input>
<ID>N_in0</ID>2842 </input>
<input>
<ID>N_in1</ID>4187 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3974</ID>
<type>HA_JUNC_2</type>
<position>369,-579.5</position>
<input>
<ID>N_in0</ID>2841 </input>
<input>
<ID>N_in1</ID>4185 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3975</ID>
<type>HA_JUNC_2</type>
<position>338.5,-579.5</position>
<input>
<ID>N_in0</ID>2840 </input>
<input>
<ID>N_in1</ID>4183 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3976</ID>
<type>HA_JUNC_2</type>
<position>306.5,-579.5</position>
<input>
<ID>N_in0</ID>2839 </input>
<input>
<ID>N_in1</ID>4181 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>3977</ID>
<type>BE_DECODER_3x8</type>
<position>196.5,-652</position>
<input>
<ID>ENABLE</ID>73 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>2853 </output>
<output>
<ID>OUT_1</ID>2852 </output>
<output>
<ID>OUT_2</ID>2851 </output>
<output>
<ID>OUT_3</ID>2850 </output>
<output>
<ID>OUT_4</ID>2849 </output>
<output>
<ID>OUT_5</ID>2848 </output>
<output>
<ID>OUT_6</ID>2847 </output>
<output>
<ID>OUT_7</ID>2846 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>3978</ID>
<type>BA_TRI_STATE</type>
<position>238.5,-666.5</position>
<input>
<ID>ENABLE_0</ID>2850 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2762 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3979</ID>
<type>AA_AND2</type>
<position>232.5,-662</position>
<input>
<ID>IN_0</ID>2850 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2761 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3980</ID>
<type>BA_TRI_STATE</type>
<position>238.5,-682.5</position>
<input>
<ID>ENABLE_0</ID>2851 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2764 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3981</ID>
<type>AA_AND2</type>
<position>232.5,-677.5</position>
<input>
<ID>IN_0</ID>2851 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2763 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3982</ID>
<type>BA_TRI_STATE</type>
<position>238.5,-698.5</position>
<input>
<ID>ENABLE_0</ID>2852 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2828 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3983</ID>
<type>AA_AND2</type>
<position>232.5,-693.5</position>
<input>
<ID>IN_0</ID>2852 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2827 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3984</ID>
<type>BA_TRI_STATE</type>
<position>238.5,-715.5</position>
<input>
<ID>ENABLE_0</ID>2853 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2830 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3985</ID>
<type>AA_AND2</type>
<position>232.5,-710.5</position>
<input>
<ID>IN_0</ID>2853 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2829 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3986</ID>
<type>AA_AND2</type>
<position>263.5,-652</position>
<input>
<ID>IN_0</ID>2855 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2854 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3987</ID>
<type>BA_TRI_STATE</type>
<position>270.5,-652</position>
<input>
<ID>ENABLE_0</ID>2854 </input>
<input>
<ID>IN_0</ID>2855 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3988</ID>
<type>AE_DFF_LOW</type>
<position>251.5,-644.5</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2855 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3989</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-601.5</position>
<input>
<ID>ENABLE_0</ID>2846 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2919 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3990</ID>
<type>AA_AND2</type>
<position>233,-597</position>
<input>
<ID>IN_0</ID>2846 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2920 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3991</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-617.5</position>
<input>
<ID>ENABLE_0</ID>2847 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2755 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3992</ID>
<type>AA_AND2</type>
<position>295,-652</position>
<input>
<ID>IN_0</ID>2857 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2856 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3993</ID>
<type>AA_AND2</type>
<position>232.5,-612.5</position>
<input>
<ID>IN_0</ID>2847 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2756 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3994</ID>
<type>BA_TRI_STATE</type>
<position>302,-652</position>
<input>
<ID>ENABLE_0</ID>2856 </input>
<input>
<ID>IN_0</ID>2857 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3995</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-633.5</position>
<input>
<ID>ENABLE_0</ID>2848 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2757 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3996</ID>
<type>AE_DFF_LOW</type>
<position>282.5,-644.5</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2857 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3997</ID>
<type>AA_AND2</type>
<position>232.5,-628.5</position>
<input>
<ID>IN_0</ID>2848 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2758 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3998</ID>
<type>AA_AND2</type>
<position>325.5,-652</position>
<input>
<ID>IN_0</ID>2859 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2858 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3999</ID>
<type>BA_TRI_STATE</type>
<position>239.5,-650.5</position>
<input>
<ID>ENABLE_0</ID>2849 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2760 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4000</ID>
<type>BA_TRI_STATE</type>
<position>332.5,-652</position>
<input>
<ID>ENABLE_0</ID>2858 </input>
<input>
<ID>IN_0</ID>2859 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4001</ID>
<type>AA_AND2</type>
<position>232.5,-645.5</position>
<input>
<ID>IN_0</ID>2849 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2759 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4002</ID>
<type>AE_DFF_LOW</type>
<position>313.5,-644.5</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2859 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4003</ID>
<type>AA_AND2</type>
<position>357,-652</position>
<input>
<ID>IN_0</ID>2861 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2860 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4004</ID>
<type>BA_TRI_STATE</type>
<position>364,-652</position>
<input>
<ID>ENABLE_0</ID>2860 </input>
<input>
<ID>IN_0</ID>2861 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4005</ID>
<type>AE_DFF_LOW</type>
<position>344.5,-644.5</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2861 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4006</ID>
<type>AA_AND2</type>
<position>386.5,-652</position>
<input>
<ID>IN_0</ID>2863 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2862 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4007</ID>
<type>BA_TRI_STATE</type>
<position>393.5,-652</position>
<input>
<ID>ENABLE_0</ID>2862 </input>
<input>
<ID>IN_0</ID>2863 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4008</ID>
<type>AE_DFF_LOW</type>
<position>374.5,-644.5</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2863 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4009</ID>
<type>AA_AND2</type>
<position>418,-652</position>
<input>
<ID>IN_0</ID>2865 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2864 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4010</ID>
<type>BA_TRI_STATE</type>
<position>425,-652</position>
<input>
<ID>ENABLE_0</ID>2864 </input>
<input>
<ID>IN_0</ID>2865 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4011</ID>
<type>AE_DFF_LOW</type>
<position>405.5,-644.5</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2865 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4012</ID>
<type>AA_AND2</type>
<position>448.5,-652</position>
<input>
<ID>IN_0</ID>2867 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2866 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4013</ID>
<type>BA_TRI_STATE</type>
<position>455.5,-652</position>
<input>
<ID>ENABLE_0</ID>2866 </input>
<input>
<ID>IN_0</ID>2867 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4014</ID>
<type>AE_DFF_LOW</type>
<position>436.5,-644.5</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2867 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4015</ID>
<type>AA_AND2</type>
<position>480,-652</position>
<input>
<ID>IN_0</ID>2869 </input>
<input>
<ID>IN_1</ID>2760 </input>
<output>
<ID>OUT</ID>2868 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4016</ID>
<type>BA_TRI_STATE</type>
<position>487,-652</position>
<input>
<ID>ENABLE_0</ID>2868 </input>
<input>
<ID>IN_0</ID>2869 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4017</ID>
<type>AE_DFF_LOW</type>
<position>467.5,-644.5</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2869 </output>
<input>
<ID>clock</ID>2759 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4018</ID>
<type>AA_AND2</type>
<position>264,-635</position>
<input>
<ID>IN_0</ID>2871 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2870 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4019</ID>
<type>BA_TRI_STATE</type>
<position>271,-635</position>
<input>
<ID>ENABLE_0</ID>2870 </input>
<input>
<ID>IN_0</ID>2871 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4020</ID>
<type>AE_DFF_LOW</type>
<position>252,-627.5</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2871 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4021</ID>
<type>AA_AND2</type>
<position>295.5,-635</position>
<input>
<ID>IN_0</ID>2873 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2872 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4022</ID>
<type>BA_TRI_STATE</type>
<position>302.5,-635</position>
<input>
<ID>ENABLE_0</ID>2872 </input>
<input>
<ID>IN_0</ID>2873 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4023</ID>
<type>AE_DFF_LOW</type>
<position>283,-627.5</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2873 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4024</ID>
<type>AA_AND2</type>
<position>326,-635</position>
<input>
<ID>IN_0</ID>2875 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2874 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4025</ID>
<type>BA_TRI_STATE</type>
<position>333,-635</position>
<input>
<ID>ENABLE_0</ID>2874 </input>
<input>
<ID>IN_0</ID>2875 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4026</ID>
<type>AE_DFF_LOW</type>
<position>314,-627.5</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2875 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4027</ID>
<type>AA_AND2</type>
<position>357.5,-635</position>
<input>
<ID>IN_0</ID>2877 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2876 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4028</ID>
<type>BA_TRI_STATE</type>
<position>364.5,-635</position>
<input>
<ID>ENABLE_0</ID>2876 </input>
<input>
<ID>IN_0</ID>2877 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4029</ID>
<type>AE_DFF_LOW</type>
<position>345,-627.5</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2877 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4030</ID>
<type>AA_AND2</type>
<position>387,-635</position>
<input>
<ID>IN_0</ID>2879 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2878 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4031</ID>
<type>BA_TRI_STATE</type>
<position>394,-635</position>
<input>
<ID>ENABLE_0</ID>2878 </input>
<input>
<ID>IN_0</ID>2879 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4032</ID>
<type>AE_DFF_LOW</type>
<position>375,-627.5</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2879 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4033</ID>
<type>AA_AND2</type>
<position>418.5,-635</position>
<input>
<ID>IN_0</ID>2881 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2880 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4034</ID>
<type>BA_TRI_STATE</type>
<position>425.5,-635</position>
<input>
<ID>ENABLE_0</ID>2880 </input>
<input>
<ID>IN_0</ID>2881 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4035</ID>
<type>AE_DFF_LOW</type>
<position>406,-627.5</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2881 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4036</ID>
<type>AA_AND2</type>
<position>449,-635</position>
<input>
<ID>IN_0</ID>2883 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2882 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4037</ID>
<type>BA_TRI_STATE</type>
<position>456,-635</position>
<input>
<ID>ENABLE_0</ID>2882 </input>
<input>
<ID>IN_0</ID>2883 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4038</ID>
<type>AE_DFF_LOW</type>
<position>437,-627.5</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2883 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4039</ID>
<type>AA_AND2</type>
<position>480.5,-635</position>
<input>
<ID>IN_0</ID>2885 </input>
<input>
<ID>IN_1</ID>2757 </input>
<output>
<ID>OUT</ID>2884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4040</ID>
<type>BA_TRI_STATE</type>
<position>487.5,-635</position>
<input>
<ID>ENABLE_0</ID>2884 </input>
<input>
<ID>IN_0</ID>2885 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4041</ID>
<type>AE_DFF_LOW</type>
<position>468,-627.5</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2885 </output>
<input>
<ID>clock</ID>2758 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4042</ID>
<type>AA_AND2</type>
<position>264.5,-619</position>
<input>
<ID>IN_0</ID>2887 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2886 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4043</ID>
<type>BA_TRI_STATE</type>
<position>271.5,-619</position>
<input>
<ID>ENABLE_0</ID>2886 </input>
<input>
<ID>IN_0</ID>2887 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4044</ID>
<type>AE_DFF_LOW</type>
<position>252.5,-611.5</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2887 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4045</ID>
<type>AA_AND2</type>
<position>296,-619</position>
<input>
<ID>IN_0</ID>2889 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2888 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4046</ID>
<type>BA_TRI_STATE</type>
<position>303,-619</position>
<input>
<ID>ENABLE_0</ID>2888 </input>
<input>
<ID>IN_0</ID>2889 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4047</ID>
<type>AE_DFF_LOW</type>
<position>283.5,-611.5</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2889 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4048</ID>
<type>AA_AND2</type>
<position>326.5,-619</position>
<input>
<ID>IN_0</ID>2891 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2890 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4049</ID>
<type>BA_TRI_STATE</type>
<position>333.5,-619</position>
<input>
<ID>ENABLE_0</ID>2890 </input>
<input>
<ID>IN_0</ID>2891 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4050</ID>
<type>AE_DFF_LOW</type>
<position>314.5,-611.5</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2891 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4051</ID>
<type>AA_AND2</type>
<position>358,-619</position>
<input>
<ID>IN_0</ID>2893 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2892 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4052</ID>
<type>BA_TRI_STATE</type>
<position>365,-619</position>
<input>
<ID>ENABLE_0</ID>2892 </input>
<input>
<ID>IN_0</ID>2893 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4053</ID>
<type>AE_DFF_LOW</type>
<position>345.5,-611.5</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2893 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4054</ID>
<type>AA_AND2</type>
<position>387.5,-619</position>
<input>
<ID>IN_0</ID>2895 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2894 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4055</ID>
<type>BA_TRI_STATE</type>
<position>394.5,-619</position>
<input>
<ID>ENABLE_0</ID>2894 </input>
<input>
<ID>IN_0</ID>2895 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4056</ID>
<type>AE_DFF_LOW</type>
<position>375.5,-611.5</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2895 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4057</ID>
<type>AA_AND2</type>
<position>419,-619</position>
<input>
<ID>IN_0</ID>2897 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2896 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4058</ID>
<type>BA_TRI_STATE</type>
<position>426,-619</position>
<input>
<ID>ENABLE_0</ID>2896 </input>
<input>
<ID>IN_0</ID>2897 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4059</ID>
<type>AE_DFF_LOW</type>
<position>406.5,-611.5</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2897 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4060</ID>
<type>AA_AND2</type>
<position>449.5,-619</position>
<input>
<ID>IN_0</ID>2899 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2898 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4061</ID>
<type>BA_TRI_STATE</type>
<position>456.5,-619</position>
<input>
<ID>ENABLE_0</ID>2898 </input>
<input>
<ID>IN_0</ID>2899 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4062</ID>
<type>AE_DFF_LOW</type>
<position>437.5,-611.5</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2899 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4063</ID>
<type>AA_AND2</type>
<position>481,-619</position>
<input>
<ID>IN_0</ID>2901 </input>
<input>
<ID>IN_1</ID>2755 </input>
<output>
<ID>OUT</ID>2900 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4064</ID>
<type>BA_TRI_STATE</type>
<position>488,-619</position>
<input>
<ID>ENABLE_0</ID>2900 </input>
<input>
<ID>IN_0</ID>2901 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4065</ID>
<type>AE_DFF_LOW</type>
<position>468.5,-611.5</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2901 </output>
<input>
<ID>clock</ID>2756 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4066</ID>
<type>AA_AND2</type>
<position>265,-603.5</position>
<input>
<ID>IN_0</ID>2903 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2902 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4067</ID>
<type>BA_TRI_STATE</type>
<position>272,-603.5</position>
<input>
<ID>ENABLE_0</ID>2902 </input>
<input>
<ID>IN_0</ID>2903 </input>
<output>
<ID>OUT_0</ID>2838 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4068</ID>
<type>AE_DFF_LOW</type>
<position>253,-596</position>
<input>
<ID>IN_0</ID>2918 </input>
<output>
<ID>OUT_0</ID>2903 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4069</ID>
<type>AA_AND2</type>
<position>296.5,-603.5</position>
<input>
<ID>IN_0</ID>2905 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2904 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4070</ID>
<type>BA_TRI_STATE</type>
<position>303.5,-603.5</position>
<input>
<ID>ENABLE_0</ID>2904 </input>
<input>
<ID>IN_0</ID>2905 </input>
<output>
<ID>OUT_0</ID>2839 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4071</ID>
<type>AE_DFF_LOW</type>
<position>284,-596</position>
<input>
<ID>IN_0</ID>2831 </input>
<output>
<ID>OUT_0</ID>2905 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4072</ID>
<type>AA_AND2</type>
<position>327,-603.5</position>
<input>
<ID>IN_0</ID>2907 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2906 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4073</ID>
<type>BA_TRI_STATE</type>
<position>334,-603.5</position>
<input>
<ID>ENABLE_0</ID>2906 </input>
<input>
<ID>IN_0</ID>2907 </input>
<output>
<ID>OUT_0</ID>2840 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4074</ID>
<type>AE_DFF_LOW</type>
<position>315,-596</position>
<input>
<ID>IN_0</ID>2832 </input>
<output>
<ID>OUT_0</ID>2907 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4075</ID>
<type>AA_AND2</type>
<position>358.5,-603.5</position>
<input>
<ID>IN_0</ID>2909 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2908 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4076</ID>
<type>BA_TRI_STATE</type>
<position>365.5,-603.5</position>
<input>
<ID>ENABLE_0</ID>2908 </input>
<input>
<ID>IN_0</ID>2909 </input>
<output>
<ID>OUT_0</ID>2841 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4077</ID>
<type>AE_DFF_LOW</type>
<position>346,-596</position>
<input>
<ID>IN_0</ID>2833 </input>
<output>
<ID>OUT_0</ID>2909 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4078</ID>
<type>AA_AND2</type>
<position>388,-603.5</position>
<input>
<ID>IN_0</ID>2911 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2910 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4079</ID>
<type>BA_TRI_STATE</type>
<position>395,-603.5</position>
<input>
<ID>ENABLE_0</ID>2910 </input>
<input>
<ID>IN_0</ID>2911 </input>
<output>
<ID>OUT_0</ID>2842 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4080</ID>
<type>AE_DFF_LOW</type>
<position>376,-596</position>
<input>
<ID>IN_0</ID>2834 </input>
<output>
<ID>OUT_0</ID>2911 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4081</ID>
<type>AA_AND2</type>
<position>419.5,-603.5</position>
<input>
<ID>IN_0</ID>2913 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2912 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4082</ID>
<type>BA_TRI_STATE</type>
<position>426.5,-603.5</position>
<input>
<ID>ENABLE_0</ID>2912 </input>
<input>
<ID>IN_0</ID>2913 </input>
<output>
<ID>OUT_0</ID>2843 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4083</ID>
<type>AE_DFF_LOW</type>
<position>407,-596</position>
<input>
<ID>IN_0</ID>2835 </input>
<output>
<ID>OUT_0</ID>2913 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4084</ID>
<type>AA_AND2</type>
<position>450,-603.5</position>
<input>
<ID>IN_0</ID>2915 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2914 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4085</ID>
<type>BA_TRI_STATE</type>
<position>457,-603.5</position>
<input>
<ID>ENABLE_0</ID>2914 </input>
<input>
<ID>IN_0</ID>2915 </input>
<output>
<ID>OUT_0</ID>2844 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4086</ID>
<type>AE_DFF_LOW</type>
<position>438,-596</position>
<input>
<ID>IN_0</ID>2836 </input>
<output>
<ID>OUT_0</ID>2915 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4087</ID>
<type>AA_AND2</type>
<position>481.5,-603.5</position>
<input>
<ID>IN_0</ID>2917 </input>
<input>
<ID>IN_1</ID>2919 </input>
<output>
<ID>OUT</ID>2916 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4088</ID>
<type>BA_TRI_STATE</type>
<position>488.5,-603.5</position>
<input>
<ID>ENABLE_0</ID>2916 </input>
<input>
<ID>IN_0</ID>2917 </input>
<output>
<ID>OUT_0</ID>2845 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4089</ID>
<type>AE_DFF_LOW</type>
<position>469,-596</position>
<input>
<ID>IN_0</ID>2837 </input>
<output>
<ID>OUT_0</ID>2917 </output>
<input>
<ID>clock</ID>2920 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4090</ID>
<type>AA_AND2</type>
<position>266.5,22</position>
<input>
<ID>IN_0</ID>2922 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2921 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4091</ID>
<type>BA_TRI_STATE</type>
<position>273.5,22</position>
<input>
<ID>ENABLE_0</ID>2921 </input>
<input>
<ID>IN_0</ID>2922 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4092</ID>
<type>AE_DFF_LOW</type>
<position>254.5,29.5</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>2922 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4093</ID>
<type>HA_JUNC_2</type>
<position>250.5,11</position>
<input>
<ID>N_in0</ID>4130 </input>
<input>
<ID>N_in1</ID>3086 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4094</ID>
<type>HA_JUNC_2</type>
<position>281.5,10.5</position>
<input>
<ID>N_in0</ID>4132 </input>
<input>
<ID>N_in1</ID>2999 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4095</ID>
<type>HA_JUNC_2</type>
<position>313.5,10.5</position>
<input>
<ID>N_in0</ID>4134 </input>
<input>
<ID>N_in1</ID>3000 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4096</ID>
<type>HA_JUNC_2</type>
<position>344.5,11.5</position>
<input>
<ID>N_in0</ID>4136 </input>
<input>
<ID>N_in1</ID>3001 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4097</ID>
<type>HA_JUNC_2</type>
<position>374.5,12.5</position>
<input>
<ID>N_in0</ID>4138 </input>
<input>
<ID>N_in1</ID>3002 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4098</ID>
<type>HA_JUNC_2</type>
<position>405.5,13</position>
<input>
<ID>N_in0</ID>4140 </input>
<input>
<ID>N_in1</ID>3003 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4099</ID>
<type>HA_JUNC_2</type>
<position>467.5,12</position>
<input>
<ID>N_in0</ID>4144 </input>
<input>
<ID>N_in1</ID>3005 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4100</ID>
<type>HA_JUNC_2</type>
<position>436.5,14</position>
<input>
<ID>N_in0</ID>4142 </input>
<input>
<ID>N_in1</ID>3004 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4101</ID>
<type>HA_JUNC_2</type>
<position>250.5,152.5</position>
<input>
<ID>N_in0</ID>3086 </input>
<input>
<ID>N_in1</ID>4128 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4102</ID>
<type>HA_JUNC_2</type>
<position>281.5,152.5</position>
<input>
<ID>N_in0</ID>2999 </input>
<input>
<ID>N_in1</ID>4127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4103</ID>
<type>HA_JUNC_2</type>
<position>313.5,152.5</position>
<input>
<ID>N_in0</ID>3000 </input>
<input>
<ID>N_in1</ID>4125 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4104</ID>
<type>AA_AND2</type>
<position>298,22</position>
<input>
<ID>IN_0</ID>2934 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2933 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4105</ID>
<type>BA_TRI_STATE</type>
<position>305,22</position>
<input>
<ID>ENABLE_0</ID>2933 </input>
<input>
<ID>IN_0</ID>2934 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4106</ID>
<type>AE_DFF_LOW</type>
<position>285.5,29.5</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>2934 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4107</ID>
<type>AA_AND2</type>
<position>328.5,22</position>
<input>
<ID>IN_0</ID>2936 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2935 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4108</ID>
<type>BA_TRI_STATE</type>
<position>335.5,22</position>
<input>
<ID>ENABLE_0</ID>2935 </input>
<input>
<ID>IN_0</ID>2936 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4109</ID>
<type>AE_DFF_LOW</type>
<position>316.5,29.5</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>2936 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4110</ID>
<type>AA_AND2</type>
<position>360,22</position>
<input>
<ID>IN_0</ID>2938 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2937 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4111</ID>
<type>BA_TRI_STATE</type>
<position>367,22</position>
<input>
<ID>ENABLE_0</ID>2937 </input>
<input>
<ID>IN_0</ID>2938 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4112</ID>
<type>AE_DFF_LOW</type>
<position>347.5,29.5</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>2938 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4113</ID>
<type>AA_AND2</type>
<position>389.5,22</position>
<input>
<ID>IN_0</ID>2940 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2939 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4114</ID>
<type>BA_TRI_STATE</type>
<position>396.5,22</position>
<input>
<ID>ENABLE_0</ID>2939 </input>
<input>
<ID>IN_0</ID>2940 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4115</ID>
<type>AE_DFF_LOW</type>
<position>377.5,29.5</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>2940 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4116</ID>
<type>AA_AND2</type>
<position>421,22</position>
<input>
<ID>IN_0</ID>2942 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2941 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4117</ID>
<type>BA_TRI_STATE</type>
<position>428,22</position>
<input>
<ID>ENABLE_0</ID>2941 </input>
<input>
<ID>IN_0</ID>2942 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4118</ID>
<type>AE_DFF_LOW</type>
<position>408.5,29.5</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>2942 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4119</ID>
<type>AA_AND2</type>
<position>451.5,22</position>
<input>
<ID>IN_0</ID>2944 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2943 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4120</ID>
<type>BA_TRI_STATE</type>
<position>458.5,22</position>
<input>
<ID>ENABLE_0</ID>2943 </input>
<input>
<ID>IN_0</ID>2944 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4121</ID>
<type>AE_DFF_LOW</type>
<position>439.5,29.5</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>2944 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4122</ID>
<type>AA_AND2</type>
<position>483,22</position>
<input>
<ID>IN_0</ID>2946 </input>
<input>
<ID>IN_1</ID>2998 </input>
<output>
<ID>OUT</ID>2945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4123</ID>
<type>BA_TRI_STATE</type>
<position>490,22</position>
<input>
<ID>ENABLE_0</ID>2945 </input>
<input>
<ID>IN_0</ID>2946 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4124</ID>
<type>AE_DFF_LOW</type>
<position>470.5,29.5</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>2946 </output>
<input>
<ID>clock</ID>2997 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4125</ID>
<type>AA_AND2</type>
<position>267,39</position>
<input>
<ID>IN_0</ID>2948 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2947 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4126</ID>
<type>BA_TRI_STATE</type>
<position>274,39</position>
<input>
<ID>ENABLE_0</ID>2947 </input>
<input>
<ID>IN_0</ID>2948 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4127</ID>
<type>AE_DFF_LOW</type>
<position>255,46.5</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>2948 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4128</ID>
<type>AA_AND2</type>
<position>298.5,39</position>
<input>
<ID>IN_0</ID>2950 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2949 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4129</ID>
<type>BA_TRI_STATE</type>
<position>305.5,39</position>
<input>
<ID>ENABLE_0</ID>2949 </input>
<input>
<ID>IN_0</ID>2950 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4130</ID>
<type>AE_DFF_LOW</type>
<position>286,46.5</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>2950 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4131</ID>
<type>AA_AND2</type>
<position>329,39</position>
<input>
<ID>IN_0</ID>2952 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2951 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4132</ID>
<type>BA_TRI_STATE</type>
<position>336,39</position>
<input>
<ID>ENABLE_0</ID>2951 </input>
<input>
<ID>IN_0</ID>2952 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4133</ID>
<type>AE_DFF_LOW</type>
<position>317,46.5</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>2952 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4134</ID>
<type>AA_AND2</type>
<position>360.5,39</position>
<input>
<ID>IN_0</ID>2954 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2953 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4135</ID>
<type>BA_TRI_STATE</type>
<position>367.5,39</position>
<input>
<ID>ENABLE_0</ID>2953 </input>
<input>
<ID>IN_0</ID>2954 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4136</ID>
<type>AE_DFF_LOW</type>
<position>348,46.5</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>2954 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4137</ID>
<type>AA_AND2</type>
<position>390,39</position>
<input>
<ID>IN_0</ID>2956 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2955 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4138</ID>
<type>BA_TRI_STATE</type>
<position>397,39</position>
<input>
<ID>ENABLE_0</ID>2955 </input>
<input>
<ID>IN_0</ID>2956 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4139</ID>
<type>AE_DFF_LOW</type>
<position>378,46.5</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>2956 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4140</ID>
<type>AA_AND2</type>
<position>421.5,39</position>
<input>
<ID>IN_0</ID>2958 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2957 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4141</ID>
<type>BA_TRI_STATE</type>
<position>428.5,39</position>
<input>
<ID>ENABLE_0</ID>2957 </input>
<input>
<ID>IN_0</ID>2958 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4142</ID>
<type>AE_DFF_LOW</type>
<position>409,46.5</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>2958 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4143</ID>
<type>AA_AND2</type>
<position>452,39</position>
<input>
<ID>IN_0</ID>2960 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2959 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4144</ID>
<type>BA_TRI_STATE</type>
<position>459,39</position>
<input>
<ID>ENABLE_0</ID>2959 </input>
<input>
<ID>IN_0</ID>2960 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4145</ID>
<type>AE_DFF_LOW</type>
<position>440,46.5</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>2960 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4146</ID>
<type>AA_AND2</type>
<position>483.5,39</position>
<input>
<ID>IN_0</ID>2962 </input>
<input>
<ID>IN_1</ID>2996 </input>
<output>
<ID>OUT</ID>2961 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4147</ID>
<type>BA_TRI_STATE</type>
<position>490.5,39</position>
<input>
<ID>ENABLE_0</ID>2961 </input>
<input>
<ID>IN_0</ID>2962 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4148</ID>
<type>AE_DFF_LOW</type>
<position>471,46.5</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>2962 </output>
<input>
<ID>clock</ID>2995 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4149</ID>
<type>AA_AND2</type>
<position>267.5,55</position>
<input>
<ID>IN_0</ID>2964 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2963 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4150</ID>
<type>BA_TRI_STATE</type>
<position>274.5,55</position>
<input>
<ID>ENABLE_0</ID>2963 </input>
<input>
<ID>IN_0</ID>2964 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4151</ID>
<type>AE_DFF_LOW</type>
<position>255.5,62.5</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>2964 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4152</ID>
<type>AA_AND2</type>
<position>299,55</position>
<input>
<ID>IN_0</ID>2966 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2965 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4153</ID>
<type>BA_TRI_STATE</type>
<position>306,55</position>
<input>
<ID>ENABLE_0</ID>2965 </input>
<input>
<ID>IN_0</ID>2966 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4154</ID>
<type>AE_DFF_LOW</type>
<position>286.5,62.5</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>2966 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4155</ID>
<type>AA_AND2</type>
<position>329.5,55</position>
<input>
<ID>IN_0</ID>2968 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2967 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4156</ID>
<type>BA_TRI_STATE</type>
<position>336.5,55</position>
<input>
<ID>ENABLE_0</ID>2967 </input>
<input>
<ID>IN_0</ID>2968 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4157</ID>
<type>AE_DFF_LOW</type>
<position>317.5,62.5</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>2968 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4158</ID>
<type>AA_AND2</type>
<position>361,55</position>
<input>
<ID>IN_0</ID>2970 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2969 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4159</ID>
<type>BA_TRI_STATE</type>
<position>368,55</position>
<input>
<ID>ENABLE_0</ID>2969 </input>
<input>
<ID>IN_0</ID>2970 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4160</ID>
<type>AE_DFF_LOW</type>
<position>348.5,62.5</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>2970 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4161</ID>
<type>AA_AND2</type>
<position>390.5,55</position>
<input>
<ID>IN_0</ID>2972 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2971 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4162</ID>
<type>BA_TRI_STATE</type>
<position>397.5,55</position>
<input>
<ID>ENABLE_0</ID>2971 </input>
<input>
<ID>IN_0</ID>2972 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4163</ID>
<type>AE_DFF_LOW</type>
<position>378.5,62.5</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>2972 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4164</ID>
<type>AA_AND2</type>
<position>422,55</position>
<input>
<ID>IN_0</ID>2974 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2973 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4165</ID>
<type>BA_TRI_STATE</type>
<position>429,55</position>
<input>
<ID>ENABLE_0</ID>2973 </input>
<input>
<ID>IN_0</ID>2974 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4166</ID>
<type>AE_DFF_LOW</type>
<position>409.5,62.5</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>2974 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4167</ID>
<type>AA_AND2</type>
<position>452.5,55</position>
<input>
<ID>IN_0</ID>2976 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2975 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4168</ID>
<type>BA_TRI_STATE</type>
<position>459.5,55</position>
<input>
<ID>ENABLE_0</ID>2975 </input>
<input>
<ID>IN_0</ID>2976 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4169</ID>
<type>AE_DFF_LOW</type>
<position>440.5,62.5</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>2976 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4170</ID>
<type>AA_AND2</type>
<position>484,55</position>
<input>
<ID>IN_0</ID>2978 </input>
<input>
<ID>IN_1</ID>2932 </input>
<output>
<ID>OUT</ID>2977 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4171</ID>
<type>BA_TRI_STATE</type>
<position>491,55</position>
<input>
<ID>ENABLE_0</ID>2977 </input>
<input>
<ID>IN_0</ID>2978 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4172</ID>
<type>AE_DFF_LOW</type>
<position>471.5,62.5</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>2978 </output>
<input>
<ID>clock</ID>2931 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4173</ID>
<type>AA_AND2</type>
<position>268,70.5</position>
<input>
<ID>IN_0</ID>2980 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2979 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4174</ID>
<type>BA_TRI_STATE</type>
<position>275,70.5</position>
<input>
<ID>ENABLE_0</ID>2979 </input>
<input>
<ID>IN_0</ID>2980 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4175</ID>
<type>AE_DFF_LOW</type>
<position>256,78</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>2980 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4176</ID>
<type>AA_AND2</type>
<position>299.5,70.5</position>
<input>
<ID>IN_0</ID>2982 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2981 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4177</ID>
<type>BA_TRI_STATE</type>
<position>306.5,70.5</position>
<input>
<ID>ENABLE_0</ID>2981 </input>
<input>
<ID>IN_0</ID>2982 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4178</ID>
<type>AE_DFF_LOW</type>
<position>287,78</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>2982 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4179</ID>
<type>AA_AND2</type>
<position>330,70.5</position>
<input>
<ID>IN_0</ID>2984 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2983 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4180</ID>
<type>BA_TRI_STATE</type>
<position>337,70.5</position>
<input>
<ID>ENABLE_0</ID>2983 </input>
<input>
<ID>IN_0</ID>2984 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4181</ID>
<type>AE_DFF_LOW</type>
<position>318,78</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>2984 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4182</ID>
<type>AA_AND2</type>
<position>361.5,70.5</position>
<input>
<ID>IN_0</ID>2986 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2985 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4183</ID>
<type>BA_TRI_STATE</type>
<position>368.5,70.5</position>
<input>
<ID>ENABLE_0</ID>2985 </input>
<input>
<ID>IN_0</ID>2986 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4184</ID>
<type>AE_DFF_LOW</type>
<position>349,78</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>2986 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4185</ID>
<type>AA_AND2</type>
<position>391,70.5</position>
<input>
<ID>IN_0</ID>2988 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2987 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4186</ID>
<type>BA_TRI_STATE</type>
<position>398,70.5</position>
<input>
<ID>ENABLE_0</ID>2987 </input>
<input>
<ID>IN_0</ID>2988 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4187</ID>
<type>AE_DFF_LOW</type>
<position>379,78</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>2988 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4188</ID>
<type>AA_AND2</type>
<position>422.5,70.5</position>
<input>
<ID>IN_0</ID>2990 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2989 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4189</ID>
<type>BA_TRI_STATE</type>
<position>429.5,70.5</position>
<input>
<ID>ENABLE_0</ID>2989 </input>
<input>
<ID>IN_0</ID>2990 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4190</ID>
<type>AE_DFF_LOW</type>
<position>410,78</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>2990 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4191</ID>
<type>AA_AND2</type>
<position>453,70.5</position>
<input>
<ID>IN_0</ID>2992 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2991 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4192</ID>
<type>BA_TRI_STATE</type>
<position>460,70.5</position>
<input>
<ID>ENABLE_0</ID>2991 </input>
<input>
<ID>IN_0</ID>2992 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4193</ID>
<type>AE_DFF_LOW</type>
<position>441,78</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>2992 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4194</ID>
<type>AA_AND2</type>
<position>484.5,70.5</position>
<input>
<ID>IN_0</ID>2994 </input>
<input>
<ID>IN_1</ID>2930 </input>
<output>
<ID>OUT</ID>2993 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4195</ID>
<type>BA_TRI_STATE</type>
<position>491.5,70.5</position>
<input>
<ID>ENABLE_0</ID>2993 </input>
<input>
<ID>IN_0</ID>2994 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4196</ID>
<type>AE_DFF_LOW</type>
<position>472,78</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>2994 </output>
<input>
<ID>clock</ID>2929 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4197</ID>
<type>HA_JUNC_2</type>
<position>344.5,152.5</position>
<input>
<ID>N_in0</ID>3001 </input>
<input>
<ID>N_in1</ID>4124 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4198</ID>
<type>HA_JUNC_2</type>
<position>375.5,152</position>
<input>
<ID>N_in0</ID>3002 </input>
<input>
<ID>N_in1</ID>4122 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4199</ID>
<type>HA_JUNC_2</type>
<position>405.5,152.5</position>
<input>
<ID>N_in0</ID>3003 </input>
<input>
<ID>N_in1</ID>4120 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4200</ID>
<type>HA_JUNC_2</type>
<position>436.5,152.5</position>
<input>
<ID>N_in0</ID>3004 </input>
<input>
<ID>N_in1</ID>4117 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4201</ID>
<type>HA_JUNC_2</type>
<position>467.5,152</position>
<input>
<ID>N_in0</ID>3005 </input>
<input>
<ID>N_in1</ID>4115 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4202</ID>
<type>HA_JUNC_2</type>
<position>279.5,159.5</position>
<input>
<ID>N_in0</ID>3006 </input>
<input>
<ID>N_in1</ID>4126 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4203</ID>
<type>HA_JUNC_2</type>
<position>279.5,2.5</position>
<input>
<ID>N_in0</ID>4131 </input>
<input>
<ID>N_in1</ID>3006 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4204</ID>
<type>HA_JUNC_2</type>
<position>342.5,3.5</position>
<input>
<ID>N_in0</ID>4135 </input>
<input>
<ID>N_in1</ID>3008 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4205</ID>
<type>HA_JUNC_2</type>
<position>373,4</position>
<input>
<ID>N_in0</ID>4137 </input>
<input>
<ID>N_in1</ID>3009 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4206</ID>
<type>HA_JUNC_2</type>
<position>403.5,4</position>
<input>
<ID>N_in0</ID>4139 </input>
<input>
<ID>N_in1</ID>3010 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4207</ID>
<type>HA_JUNC_2</type>
<position>434.5,4</position>
<input>
<ID>N_in0</ID>4141 </input>
<input>
<ID>N_in1</ID>3011 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4208</ID>
<type>HA_JUNC_2</type>
<position>465.5,3.5</position>
<input>
<ID>N_in0</ID>4143 </input>
<input>
<ID>N_in1</ID>3012 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4209</ID>
<type>HA_JUNC_2</type>
<position>496,4</position>
<input>
<ID>N_in0</ID>4145 </input>
<input>
<ID>N_in1</ID>3013 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4210</ID>
<type>HA_JUNC_2</type>
<position>496,161</position>
<input>
<ID>N_in0</ID>3013 </input>
<input>
<ID>N_in1</ID>4114 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4211</ID>
<type>HA_JUNC_2</type>
<position>465.5,160.5</position>
<input>
<ID>N_in0</ID>3012 </input>
<input>
<ID>N_in1</ID>4116 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4212</ID>
<type>HA_JUNC_2</type>
<position>434.5,159.5</position>
<input>
<ID>N_in0</ID>3011 </input>
<input>
<ID>N_in1</ID>4118 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4213</ID>
<type>HA_JUNC_2</type>
<position>403.5,159.5</position>
<input>
<ID>N_in0</ID>3010 </input>
<input>
<ID>N_in1</ID>4119 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4214</ID>
<type>HA_JUNC_2</type>
<position>373,159.5</position>
<input>
<ID>N_in0</ID>3009 </input>
<input>
<ID>N_in1</ID>4121 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4215</ID>
<type>HA_JUNC_2</type>
<position>342.5,159.5</position>
<input>
<ID>N_in0</ID>3008 </input>
<input>
<ID>N_in1</ID>4123 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4216</ID>
<type>HA_JUNC_2</type>
<position>310.5,159.5</position>
<input>
<ID>N_in0</ID>3007 </input>
<input>
<ID>N_in1</ID>4129 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4217</ID>
<type>BE_DECODER_3x8</type>
<position>200.5,87</position>
<input>
<ID>ENABLE</ID>68 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>3021 </output>
<output>
<ID>OUT_1</ID>3020 </output>
<output>
<ID>OUT_2</ID>3019 </output>
<output>
<ID>OUT_3</ID>3018 </output>
<output>
<ID>OUT_4</ID>3017 </output>
<output>
<ID>OUT_5</ID>3016 </output>
<output>
<ID>OUT_6</ID>3015 </output>
<output>
<ID>OUT_7</ID>3014 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4218</ID>
<type>BA_TRI_STATE</type>
<position>242.5,72.5</position>
<input>
<ID>ENABLE_0</ID>3018 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2930 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4219</ID>
<type>AA_AND2</type>
<position>236.5,77</position>
<input>
<ID>IN_0</ID>3018 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2929 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4220</ID>
<type>BA_TRI_STATE</type>
<position>242.5,56.5</position>
<input>
<ID>ENABLE_0</ID>3019 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2932 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4221</ID>
<type>AA_AND2</type>
<position>236.5,61.5</position>
<input>
<ID>IN_0</ID>3019 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2931 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4222</ID>
<type>BA_TRI_STATE</type>
<position>242.5,40.5</position>
<input>
<ID>ENABLE_0</ID>3020 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2996 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4223</ID>
<type>AA_AND2</type>
<position>236.5,45.5</position>
<input>
<ID>IN_0</ID>3020 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2995 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4224</ID>
<type>BA_TRI_STATE</type>
<position>242.5,23.5</position>
<input>
<ID>ENABLE_0</ID>3021 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2998 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4225</ID>
<type>AA_AND2</type>
<position>236.5,28.5</position>
<input>
<ID>IN_0</ID>3021 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2997 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4226</ID>
<type>AA_AND2</type>
<position>267.5,87</position>
<input>
<ID>IN_0</ID>3023 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3022 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4227</ID>
<type>BA_TRI_STATE</type>
<position>274.5,87</position>
<input>
<ID>ENABLE_0</ID>3022 </input>
<input>
<ID>IN_0</ID>3023 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4228</ID>
<type>AE_DFF_LOW</type>
<position>255.5,94.5</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>3023 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4229</ID>
<type>BA_TRI_STATE</type>
<position>243.5,137.5</position>
<input>
<ID>ENABLE_0</ID>3014 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3087 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4230</ID>
<type>AA_AND2</type>
<position>237,142</position>
<input>
<ID>IN_0</ID>3014 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3088 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4231</ID>
<type>BA_TRI_STATE</type>
<position>243.5,121.5</position>
<input>
<ID>ENABLE_0</ID>3015 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2923 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4232</ID>
<type>AA_AND2</type>
<position>299,87</position>
<input>
<ID>IN_0</ID>3025 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3024 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4233</ID>
<type>AA_AND2</type>
<position>236.5,126.5</position>
<input>
<ID>IN_0</ID>3015 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2924 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4234</ID>
<type>BA_TRI_STATE</type>
<position>306,87</position>
<input>
<ID>ENABLE_0</ID>3024 </input>
<input>
<ID>IN_0</ID>3025 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4235</ID>
<type>BA_TRI_STATE</type>
<position>243.5,105.5</position>
<input>
<ID>ENABLE_0</ID>3016 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2925 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4236</ID>
<type>AE_DFF_LOW</type>
<position>286.5,94.5</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>3025 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4237</ID>
<type>AA_AND2</type>
<position>236.5,110.5</position>
<input>
<ID>IN_0</ID>3016 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2926 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4238</ID>
<type>AA_AND2</type>
<position>329.5,87</position>
<input>
<ID>IN_0</ID>3027 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3026 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4239</ID>
<type>BA_TRI_STATE</type>
<position>243.5,88.5</position>
<input>
<ID>ENABLE_0</ID>3017 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>2928 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4240</ID>
<type>BA_TRI_STATE</type>
<position>336.5,87</position>
<input>
<ID>ENABLE_0</ID>3026 </input>
<input>
<ID>IN_0</ID>3027 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4241</ID>
<type>AA_AND2</type>
<position>236.5,93.5</position>
<input>
<ID>IN_0</ID>3017 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>2927 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4242</ID>
<type>AE_DFF_LOW</type>
<position>317.5,94.5</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>3027 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4243</ID>
<type>AA_AND2</type>
<position>361,87</position>
<input>
<ID>IN_0</ID>3029 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3028 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4244</ID>
<type>BA_TRI_STATE</type>
<position>368,87</position>
<input>
<ID>ENABLE_0</ID>3028 </input>
<input>
<ID>IN_0</ID>3029 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4245</ID>
<type>AE_DFF_LOW</type>
<position>348.5,94.5</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>3029 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4246</ID>
<type>AA_AND2</type>
<position>390.5,87</position>
<input>
<ID>IN_0</ID>3031 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4247</ID>
<type>BA_TRI_STATE</type>
<position>397.5,87</position>
<input>
<ID>ENABLE_0</ID>3030 </input>
<input>
<ID>IN_0</ID>3031 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4248</ID>
<type>AE_DFF_LOW</type>
<position>378.5,94.5</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>3031 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4249</ID>
<type>AA_AND2</type>
<position>422,87</position>
<input>
<ID>IN_0</ID>3033 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3032 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4250</ID>
<type>BA_TRI_STATE</type>
<position>429,87</position>
<input>
<ID>ENABLE_0</ID>3032 </input>
<input>
<ID>IN_0</ID>3033 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4251</ID>
<type>AE_DFF_LOW</type>
<position>409.5,94.5</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>3033 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4252</ID>
<type>AA_AND2</type>
<position>452.5,87</position>
<input>
<ID>IN_0</ID>3035 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3034 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4253</ID>
<type>BA_TRI_STATE</type>
<position>459.5,87</position>
<input>
<ID>ENABLE_0</ID>3034 </input>
<input>
<ID>IN_0</ID>3035 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4254</ID>
<type>AE_DFF_LOW</type>
<position>440.5,94.5</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>3035 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4255</ID>
<type>AA_AND2</type>
<position>484,87</position>
<input>
<ID>IN_0</ID>3037 </input>
<input>
<ID>IN_1</ID>2928 </input>
<output>
<ID>OUT</ID>3036 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4256</ID>
<type>BA_TRI_STATE</type>
<position>491,87</position>
<input>
<ID>ENABLE_0</ID>3036 </input>
<input>
<ID>IN_0</ID>3037 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4257</ID>
<type>AE_DFF_LOW</type>
<position>471.5,94.5</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>3037 </output>
<input>
<ID>clock</ID>2927 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4258</ID>
<type>AA_AND2</type>
<position>268,104</position>
<input>
<ID>IN_0</ID>3039 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3038 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4259</ID>
<type>BA_TRI_STATE</type>
<position>275,104</position>
<input>
<ID>ENABLE_0</ID>3038 </input>
<input>
<ID>IN_0</ID>3039 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4260</ID>
<type>AE_DFF_LOW</type>
<position>256,111.5</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>3039 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4261</ID>
<type>AA_AND2</type>
<position>299.5,104</position>
<input>
<ID>IN_0</ID>3041 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3040 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4262</ID>
<type>BA_TRI_STATE</type>
<position>306.5,104</position>
<input>
<ID>ENABLE_0</ID>3040 </input>
<input>
<ID>IN_0</ID>3041 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4263</ID>
<type>AE_DFF_LOW</type>
<position>287,111.5</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>3041 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4264</ID>
<type>AA_AND2</type>
<position>330,104</position>
<input>
<ID>IN_0</ID>3043 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3042 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4265</ID>
<type>BA_TRI_STATE</type>
<position>337,104</position>
<input>
<ID>ENABLE_0</ID>3042 </input>
<input>
<ID>IN_0</ID>3043 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4266</ID>
<type>AE_DFF_LOW</type>
<position>318,111.5</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>3043 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4267</ID>
<type>AA_AND2</type>
<position>361.5,104</position>
<input>
<ID>IN_0</ID>3045 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3044 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4268</ID>
<type>BA_TRI_STATE</type>
<position>368.5,104</position>
<input>
<ID>ENABLE_0</ID>3044 </input>
<input>
<ID>IN_0</ID>3045 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4269</ID>
<type>AE_DFF_LOW</type>
<position>349,111.5</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>3045 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4270</ID>
<type>AA_AND2</type>
<position>391,104</position>
<input>
<ID>IN_0</ID>3047 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3046 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4271</ID>
<type>BA_TRI_STATE</type>
<position>398,104</position>
<input>
<ID>ENABLE_0</ID>3046 </input>
<input>
<ID>IN_0</ID>3047 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4272</ID>
<type>AE_DFF_LOW</type>
<position>379,111.5</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>3047 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4273</ID>
<type>AA_AND2</type>
<position>422.5,104</position>
<input>
<ID>IN_0</ID>3049 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3048 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4274</ID>
<type>BA_TRI_STATE</type>
<position>429.5,104</position>
<input>
<ID>ENABLE_0</ID>3048 </input>
<input>
<ID>IN_0</ID>3049 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4275</ID>
<type>AE_DFF_LOW</type>
<position>410,111.5</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>3049 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4276</ID>
<type>AA_AND2</type>
<position>453,104</position>
<input>
<ID>IN_0</ID>3051 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3050 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4277</ID>
<type>BA_TRI_STATE</type>
<position>460,104</position>
<input>
<ID>ENABLE_0</ID>3050 </input>
<input>
<ID>IN_0</ID>3051 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4278</ID>
<type>AE_DFF_LOW</type>
<position>441,111.5</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>3051 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4279</ID>
<type>AA_AND2</type>
<position>484.5,104</position>
<input>
<ID>IN_0</ID>3053 </input>
<input>
<ID>IN_1</ID>2925 </input>
<output>
<ID>OUT</ID>3052 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4280</ID>
<type>BA_TRI_STATE</type>
<position>491.5,104</position>
<input>
<ID>ENABLE_0</ID>3052 </input>
<input>
<ID>IN_0</ID>3053 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4281</ID>
<type>AE_DFF_LOW</type>
<position>472,111.5</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>3053 </output>
<input>
<ID>clock</ID>2926 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4282</ID>
<type>AA_AND2</type>
<position>268.5,120</position>
<input>
<ID>IN_0</ID>3055 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3054 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4283</ID>
<type>BA_TRI_STATE</type>
<position>275.5,120</position>
<input>
<ID>ENABLE_0</ID>3054 </input>
<input>
<ID>IN_0</ID>3055 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4284</ID>
<type>AE_DFF_LOW</type>
<position>256.5,127.5</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>3055 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4285</ID>
<type>AA_AND2</type>
<position>300,120</position>
<input>
<ID>IN_0</ID>3057 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3056 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4286</ID>
<type>BA_TRI_STATE</type>
<position>307,120</position>
<input>
<ID>ENABLE_0</ID>3056 </input>
<input>
<ID>IN_0</ID>3057 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4287</ID>
<type>AE_DFF_LOW</type>
<position>287.5,127.5</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>3057 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4288</ID>
<type>AA_AND2</type>
<position>330.5,120</position>
<input>
<ID>IN_0</ID>3059 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3058 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4289</ID>
<type>BA_TRI_STATE</type>
<position>337.5,120</position>
<input>
<ID>ENABLE_0</ID>3058 </input>
<input>
<ID>IN_0</ID>3059 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4290</ID>
<type>AE_DFF_LOW</type>
<position>318.5,127.5</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>3059 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4291</ID>
<type>AA_AND2</type>
<position>362,120</position>
<input>
<ID>IN_0</ID>3061 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4292</ID>
<type>BA_TRI_STATE</type>
<position>369,120</position>
<input>
<ID>ENABLE_0</ID>3060 </input>
<input>
<ID>IN_0</ID>3061 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4293</ID>
<type>AE_DFF_LOW</type>
<position>349.5,127.5</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>3061 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4294</ID>
<type>AA_AND2</type>
<position>391.5,120</position>
<input>
<ID>IN_0</ID>3063 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3062 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4295</ID>
<type>BA_TRI_STATE</type>
<position>398.5,120</position>
<input>
<ID>ENABLE_0</ID>3062 </input>
<input>
<ID>IN_0</ID>3063 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4296</ID>
<type>AE_DFF_LOW</type>
<position>379.5,127.5</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>3063 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4297</ID>
<type>AA_AND2</type>
<position>423,120</position>
<input>
<ID>IN_0</ID>3065 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4298</ID>
<type>BA_TRI_STATE</type>
<position>430,120</position>
<input>
<ID>ENABLE_0</ID>3064 </input>
<input>
<ID>IN_0</ID>3065 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4299</ID>
<type>AE_DFF_LOW</type>
<position>410.5,127.5</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>3065 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4300</ID>
<type>AA_AND2</type>
<position>453.5,120</position>
<input>
<ID>IN_0</ID>3067 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3066 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4301</ID>
<type>BA_TRI_STATE</type>
<position>460.5,120</position>
<input>
<ID>ENABLE_0</ID>3066 </input>
<input>
<ID>IN_0</ID>3067 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4302</ID>
<type>AE_DFF_LOW</type>
<position>441.5,127.5</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>3067 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4303</ID>
<type>AA_AND2</type>
<position>485,120</position>
<input>
<ID>IN_0</ID>3069 </input>
<input>
<ID>IN_1</ID>2923 </input>
<output>
<ID>OUT</ID>3068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4304</ID>
<type>BA_TRI_STATE</type>
<position>492,120</position>
<input>
<ID>ENABLE_0</ID>3068 </input>
<input>
<ID>IN_0</ID>3069 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4305</ID>
<type>AE_DFF_LOW</type>
<position>472.5,127.5</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>3069 </output>
<input>
<ID>clock</ID>2924 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4306</ID>
<type>AA_AND2</type>
<position>269,135.5</position>
<input>
<ID>IN_0</ID>3071 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4307</ID>
<type>BA_TRI_STATE</type>
<position>276,135.5</position>
<input>
<ID>ENABLE_0</ID>3070 </input>
<input>
<ID>IN_0</ID>3071 </input>
<output>
<ID>OUT_0</ID>3006 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4308</ID>
<type>AE_DFF_LOW</type>
<position>257,143</position>
<input>
<ID>IN_0</ID>3086 </input>
<output>
<ID>OUT_0</ID>3071 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4309</ID>
<type>AA_AND2</type>
<position>300.5,135.5</position>
<input>
<ID>IN_0</ID>3073 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3072 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4310</ID>
<type>BA_TRI_STATE</type>
<position>307.5,135.5</position>
<input>
<ID>ENABLE_0</ID>3072 </input>
<input>
<ID>IN_0</ID>3073 </input>
<output>
<ID>OUT_0</ID>3007 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4311</ID>
<type>AE_DFF_LOW</type>
<position>288,143</position>
<input>
<ID>IN_0</ID>2999 </input>
<output>
<ID>OUT_0</ID>3073 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4312</ID>
<type>AA_AND2</type>
<position>331,135.5</position>
<input>
<ID>IN_0</ID>3075 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4313</ID>
<type>BA_TRI_STATE</type>
<position>338,135.5</position>
<input>
<ID>ENABLE_0</ID>3074 </input>
<input>
<ID>IN_0</ID>3075 </input>
<output>
<ID>OUT_0</ID>3008 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4314</ID>
<type>AE_DFF_LOW</type>
<position>319,143</position>
<input>
<ID>IN_0</ID>3000 </input>
<output>
<ID>OUT_0</ID>3075 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4315</ID>
<type>AA_AND2</type>
<position>362.5,135.5</position>
<input>
<ID>IN_0</ID>3077 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3076 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4316</ID>
<type>BA_TRI_STATE</type>
<position>369.5,135.5</position>
<input>
<ID>ENABLE_0</ID>3076 </input>
<input>
<ID>IN_0</ID>3077 </input>
<output>
<ID>OUT_0</ID>3009 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4317</ID>
<type>AE_DFF_LOW</type>
<position>350,143</position>
<input>
<ID>IN_0</ID>3001 </input>
<output>
<ID>OUT_0</ID>3077 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4318</ID>
<type>AA_AND2</type>
<position>392,135.5</position>
<input>
<ID>IN_0</ID>3079 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3078 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4319</ID>
<type>BA_TRI_STATE</type>
<position>399,135.5</position>
<input>
<ID>ENABLE_0</ID>3078 </input>
<input>
<ID>IN_0</ID>3079 </input>
<output>
<ID>OUT_0</ID>3010 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4320</ID>
<type>AE_DFF_LOW</type>
<position>380,143</position>
<input>
<ID>IN_0</ID>3002 </input>
<output>
<ID>OUT_0</ID>3079 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4321</ID>
<type>AA_AND2</type>
<position>423.5,135.5</position>
<input>
<ID>IN_0</ID>3081 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4322</ID>
<type>BA_TRI_STATE</type>
<position>430.5,135.5</position>
<input>
<ID>ENABLE_0</ID>3080 </input>
<input>
<ID>IN_0</ID>3081 </input>
<output>
<ID>OUT_0</ID>3011 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4323</ID>
<type>AE_DFF_LOW</type>
<position>411,143</position>
<input>
<ID>IN_0</ID>3003 </input>
<output>
<ID>OUT_0</ID>3081 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4324</ID>
<type>AA_AND2</type>
<position>454,135.5</position>
<input>
<ID>IN_0</ID>3083 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3082 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4325</ID>
<type>BA_TRI_STATE</type>
<position>461,135.5</position>
<input>
<ID>ENABLE_0</ID>3082 </input>
<input>
<ID>IN_0</ID>3083 </input>
<output>
<ID>OUT_0</ID>3012 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4326</ID>
<type>AE_DFF_LOW</type>
<position>442,143</position>
<input>
<ID>IN_0</ID>3004 </input>
<output>
<ID>OUT_0</ID>3083 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4327</ID>
<type>AA_AND2</type>
<position>485.5,135.5</position>
<input>
<ID>IN_0</ID>3085 </input>
<input>
<ID>IN_1</ID>3087 </input>
<output>
<ID>OUT</ID>3084 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4328</ID>
<type>BA_TRI_STATE</type>
<position>492.5,135.5</position>
<input>
<ID>ENABLE_0</ID>3084 </input>
<input>
<ID>IN_0</ID>3085 </input>
<output>
<ID>OUT_0</ID>3013 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4329</ID>
<type>AE_DFF_LOW</type>
<position>473,143</position>
<input>
<ID>IN_0</ID>3005 </input>
<output>
<ID>OUT_0</ID>3085 </output>
<input>
<ID>clock</ID>3088 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4810</ID>
<type>AA_AND2</type>
<position>261.5,203</position>
<input>
<ID>IN_0</ID>3426 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3425 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4811</ID>
<type>BA_TRI_STATE</type>
<position>268.5,203</position>
<input>
<ID>ENABLE_0</ID>3425 </input>
<input>
<ID>IN_0</ID>3426 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4812</ID>
<type>AE_DFF_LOW</type>
<position>249.5,210.5</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3426 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4813</ID>
<type>HA_JUNC_2</type>
<position>245.5,192</position>
<input>
<ID>N_in0</ID>4128 </input>
<input>
<ID>N_in1</ID>3590 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4814</ID>
<type>HA_JUNC_2</type>
<position>276.5,191.5</position>
<input>
<ID>N_in0</ID>4127 </input>
<input>
<ID>N_in1</ID>3503 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4815</ID>
<type>HA_JUNC_2</type>
<position>308.5,191.5</position>
<input>
<ID>N_in0</ID>4125 </input>
<input>
<ID>N_in1</ID>3504 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4816</ID>
<type>HA_JUNC_2</type>
<position>339.5,192.5</position>
<input>
<ID>N_in0</ID>4124 </input>
<input>
<ID>N_in1</ID>3505 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4817</ID>
<type>HA_JUNC_2</type>
<position>369.5,193.5</position>
<input>
<ID>N_in0</ID>4122 </input>
<input>
<ID>N_in1</ID>3506 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4818</ID>
<type>HA_JUNC_2</type>
<position>400.5,194</position>
<input>
<ID>N_in0</ID>4120 </input>
<input>
<ID>N_in1</ID>3507 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4819</ID>
<type>HA_JUNC_2</type>
<position>462.5,193</position>
<input>
<ID>N_in0</ID>4115 </input>
<input>
<ID>N_in1</ID>3509 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4820</ID>
<type>HA_JUNC_2</type>
<position>431.5,195</position>
<input>
<ID>N_in0</ID>4117 </input>
<input>
<ID>N_in1</ID>3508 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4821</ID>
<type>HA_JUNC_2</type>
<position>245.5,333.5</position>
<input>
<ID>N_in0</ID>3590 </input>
<input>
<ID>N_in1</ID>4097 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4822</ID>
<type>HA_JUNC_2</type>
<position>276.5,333.5</position>
<input>
<ID>N_in0</ID>3503 </input>
<input>
<ID>N_in1</ID>4099 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4823</ID>
<type>HA_JUNC_2</type>
<position>308.5,333.5</position>
<input>
<ID>N_in0</ID>3504 </input>
<input>
<ID>N_in1</ID>4102 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4824</ID>
<type>AA_AND2</type>
<position>293,203</position>
<input>
<ID>IN_0</ID>3438 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4825</ID>
<type>BA_TRI_STATE</type>
<position>300,203</position>
<input>
<ID>ENABLE_0</ID>3437 </input>
<input>
<ID>IN_0</ID>3438 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4826</ID>
<type>AE_DFF_LOW</type>
<position>280.5,210.5</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3438 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4827</ID>
<type>AA_AND2</type>
<position>323.5,203</position>
<input>
<ID>IN_0</ID>3440 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4828</ID>
<type>BA_TRI_STATE</type>
<position>330.5,203</position>
<input>
<ID>ENABLE_0</ID>3439 </input>
<input>
<ID>IN_0</ID>3440 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4829</ID>
<type>AE_DFF_LOW</type>
<position>311.5,210.5</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3440 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4830</ID>
<type>AA_AND2</type>
<position>355,203</position>
<input>
<ID>IN_0</ID>3442 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3441 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4831</ID>
<type>BA_TRI_STATE</type>
<position>362,203</position>
<input>
<ID>ENABLE_0</ID>3441 </input>
<input>
<ID>IN_0</ID>3442 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4832</ID>
<type>AE_DFF_LOW</type>
<position>342.5,210.5</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3442 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4833</ID>
<type>AA_AND2</type>
<position>384.5,203</position>
<input>
<ID>IN_0</ID>3444 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3443 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4834</ID>
<type>BA_TRI_STATE</type>
<position>391.5,203</position>
<input>
<ID>ENABLE_0</ID>3443 </input>
<input>
<ID>IN_0</ID>3444 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4835</ID>
<type>AE_DFF_LOW</type>
<position>372.5,210.5</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3444 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4836</ID>
<type>AA_AND2</type>
<position>416,203</position>
<input>
<ID>IN_0</ID>3446 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4837</ID>
<type>BA_TRI_STATE</type>
<position>423,203</position>
<input>
<ID>ENABLE_0</ID>3445 </input>
<input>
<ID>IN_0</ID>3446 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4838</ID>
<type>AE_DFF_LOW</type>
<position>403.5,210.5</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3446 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4839</ID>
<type>AA_AND2</type>
<position>446.5,203</position>
<input>
<ID>IN_0</ID>3448 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3447 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4840</ID>
<type>BA_TRI_STATE</type>
<position>453.5,203</position>
<input>
<ID>ENABLE_0</ID>3447 </input>
<input>
<ID>IN_0</ID>3448 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4841</ID>
<type>AE_DFF_LOW</type>
<position>434.5,210.5</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3448 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4842</ID>
<type>AA_AND2</type>
<position>478,203</position>
<input>
<ID>IN_0</ID>3450 </input>
<input>
<ID>IN_1</ID>3502 </input>
<output>
<ID>OUT</ID>3449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4843</ID>
<type>BA_TRI_STATE</type>
<position>485,203</position>
<input>
<ID>ENABLE_0</ID>3449 </input>
<input>
<ID>IN_0</ID>3450 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4844</ID>
<type>AE_DFF_LOW</type>
<position>465.5,210.5</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3450 </output>
<input>
<ID>clock</ID>3501 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4845</ID>
<type>AA_AND2</type>
<position>262,220</position>
<input>
<ID>IN_0</ID>3452 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4846</ID>
<type>BA_TRI_STATE</type>
<position>269,220</position>
<input>
<ID>ENABLE_0</ID>3451 </input>
<input>
<ID>IN_0</ID>3452 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4847</ID>
<type>AE_DFF_LOW</type>
<position>250,227.5</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3452 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4848</ID>
<type>AA_AND2</type>
<position>293.5,220</position>
<input>
<ID>IN_0</ID>3454 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4849</ID>
<type>BA_TRI_STATE</type>
<position>300.5,220</position>
<input>
<ID>ENABLE_0</ID>3453 </input>
<input>
<ID>IN_0</ID>3454 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4850</ID>
<type>AE_DFF_LOW</type>
<position>281,227.5</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3454 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4851</ID>
<type>AA_AND2</type>
<position>324,220</position>
<input>
<ID>IN_0</ID>3456 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3455 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4852</ID>
<type>BA_TRI_STATE</type>
<position>331,220</position>
<input>
<ID>ENABLE_0</ID>3455 </input>
<input>
<ID>IN_0</ID>3456 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4853</ID>
<type>AE_DFF_LOW</type>
<position>312,227.5</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3456 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4854</ID>
<type>AA_AND2</type>
<position>355.5,220</position>
<input>
<ID>IN_0</ID>3458 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3457 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4855</ID>
<type>BA_TRI_STATE</type>
<position>362.5,220</position>
<input>
<ID>ENABLE_0</ID>3457 </input>
<input>
<ID>IN_0</ID>3458 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4856</ID>
<type>AE_DFF_LOW</type>
<position>343,227.5</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3458 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4857</ID>
<type>AA_AND2</type>
<position>385,220</position>
<input>
<ID>IN_0</ID>3460 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3459 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4858</ID>
<type>BA_TRI_STATE</type>
<position>392,220</position>
<input>
<ID>ENABLE_0</ID>3459 </input>
<input>
<ID>IN_0</ID>3460 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4859</ID>
<type>AE_DFF_LOW</type>
<position>373,227.5</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3460 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4860</ID>
<type>AA_AND2</type>
<position>416.5,220</position>
<input>
<ID>IN_0</ID>3462 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3461 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4861</ID>
<type>BA_TRI_STATE</type>
<position>423.5,220</position>
<input>
<ID>ENABLE_0</ID>3461 </input>
<input>
<ID>IN_0</ID>3462 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4862</ID>
<type>AE_DFF_LOW</type>
<position>404,227.5</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3462 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4863</ID>
<type>AA_AND2</type>
<position>447,220</position>
<input>
<ID>IN_0</ID>3464 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3463 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4864</ID>
<type>BA_TRI_STATE</type>
<position>454,220</position>
<input>
<ID>ENABLE_0</ID>3463 </input>
<input>
<ID>IN_0</ID>3464 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4865</ID>
<type>AE_DFF_LOW</type>
<position>435,227.5</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3464 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4866</ID>
<type>AA_AND2</type>
<position>478.5,220</position>
<input>
<ID>IN_0</ID>3466 </input>
<input>
<ID>IN_1</ID>3500 </input>
<output>
<ID>OUT</ID>3465 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4867</ID>
<type>BA_TRI_STATE</type>
<position>485.5,220</position>
<input>
<ID>ENABLE_0</ID>3465 </input>
<input>
<ID>IN_0</ID>3466 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4868</ID>
<type>AE_DFF_LOW</type>
<position>466,227.5</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3466 </output>
<input>
<ID>clock</ID>3499 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4869</ID>
<type>AA_AND2</type>
<position>262.5,236</position>
<input>
<ID>IN_0</ID>3468 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3467 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4870</ID>
<type>BA_TRI_STATE</type>
<position>269.5,236</position>
<input>
<ID>ENABLE_0</ID>3467 </input>
<input>
<ID>IN_0</ID>3468 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4871</ID>
<type>AE_DFF_LOW</type>
<position>250.5,243.5</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3468 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4872</ID>
<type>AA_AND2</type>
<position>294,236</position>
<input>
<ID>IN_0</ID>3470 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3469 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4873</ID>
<type>BA_TRI_STATE</type>
<position>301,236</position>
<input>
<ID>ENABLE_0</ID>3469 </input>
<input>
<ID>IN_0</ID>3470 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4874</ID>
<type>AE_DFF_LOW</type>
<position>281.5,243.5</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3470 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4875</ID>
<type>AA_AND2</type>
<position>324.5,236</position>
<input>
<ID>IN_0</ID>3472 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3471 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4876</ID>
<type>BA_TRI_STATE</type>
<position>331.5,236</position>
<input>
<ID>ENABLE_0</ID>3471 </input>
<input>
<ID>IN_0</ID>3472 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4877</ID>
<type>AE_DFF_LOW</type>
<position>312.5,243.5</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3472 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4878</ID>
<type>AA_AND2</type>
<position>356,236</position>
<input>
<ID>IN_0</ID>3474 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3473 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4879</ID>
<type>BA_TRI_STATE</type>
<position>363,236</position>
<input>
<ID>ENABLE_0</ID>3473 </input>
<input>
<ID>IN_0</ID>3474 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4880</ID>
<type>AE_DFF_LOW</type>
<position>343.5,243.5</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3474 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4881</ID>
<type>AA_AND2</type>
<position>385.5,236</position>
<input>
<ID>IN_0</ID>3476 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3475 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4882</ID>
<type>BA_TRI_STATE</type>
<position>392.5,236</position>
<input>
<ID>ENABLE_0</ID>3475 </input>
<input>
<ID>IN_0</ID>3476 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4883</ID>
<type>AE_DFF_LOW</type>
<position>373.5,243.5</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3476 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4884</ID>
<type>AA_AND2</type>
<position>417,236</position>
<input>
<ID>IN_0</ID>3478 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3477 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4885</ID>
<type>BA_TRI_STATE</type>
<position>424,236</position>
<input>
<ID>ENABLE_0</ID>3477 </input>
<input>
<ID>IN_0</ID>3478 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4886</ID>
<type>AE_DFF_LOW</type>
<position>404.5,243.5</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3478 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4887</ID>
<type>AA_AND2</type>
<position>447.5,236</position>
<input>
<ID>IN_0</ID>3480 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4888</ID>
<type>BA_TRI_STATE</type>
<position>454.5,236</position>
<input>
<ID>ENABLE_0</ID>3479 </input>
<input>
<ID>IN_0</ID>3480 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4889</ID>
<type>AE_DFF_LOW</type>
<position>435.5,243.5</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3480 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4890</ID>
<type>AA_AND2</type>
<position>479,236</position>
<input>
<ID>IN_0</ID>3482 </input>
<input>
<ID>IN_1</ID>3436 </input>
<output>
<ID>OUT</ID>3481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4891</ID>
<type>BA_TRI_STATE</type>
<position>486,236</position>
<input>
<ID>ENABLE_0</ID>3481 </input>
<input>
<ID>IN_0</ID>3482 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4892</ID>
<type>AE_DFF_LOW</type>
<position>466.5,243.5</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3482 </output>
<input>
<ID>clock</ID>3435 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4893</ID>
<type>AA_AND2</type>
<position>263,251.5</position>
<input>
<ID>IN_0</ID>3484 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4894</ID>
<type>BA_TRI_STATE</type>
<position>270,251.5</position>
<input>
<ID>ENABLE_0</ID>3483 </input>
<input>
<ID>IN_0</ID>3484 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4895</ID>
<type>AE_DFF_LOW</type>
<position>251,259</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3484 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4896</ID>
<type>AA_AND2</type>
<position>294.5,251.5</position>
<input>
<ID>IN_0</ID>3486 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4897</ID>
<type>BA_TRI_STATE</type>
<position>301.5,251.5</position>
<input>
<ID>ENABLE_0</ID>3485 </input>
<input>
<ID>IN_0</ID>3486 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4898</ID>
<type>AE_DFF_LOW</type>
<position>282,259</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3486 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4899</ID>
<type>AA_AND2</type>
<position>325,251.5</position>
<input>
<ID>IN_0</ID>3488 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4900</ID>
<type>BA_TRI_STATE</type>
<position>332,251.5</position>
<input>
<ID>ENABLE_0</ID>3487 </input>
<input>
<ID>IN_0</ID>3488 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4901</ID>
<type>AE_DFF_LOW</type>
<position>313,259</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3488 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4902</ID>
<type>AA_AND2</type>
<position>356.5,251.5</position>
<input>
<ID>IN_0</ID>3490 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3489 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4903</ID>
<type>BA_TRI_STATE</type>
<position>363.5,251.5</position>
<input>
<ID>ENABLE_0</ID>3489 </input>
<input>
<ID>IN_0</ID>3490 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4904</ID>
<type>AE_DFF_LOW</type>
<position>344,259</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3490 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4905</ID>
<type>AA_AND2</type>
<position>386,251.5</position>
<input>
<ID>IN_0</ID>3492 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3491 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4906</ID>
<type>BA_TRI_STATE</type>
<position>393,251.5</position>
<input>
<ID>ENABLE_0</ID>3491 </input>
<input>
<ID>IN_0</ID>3492 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4907</ID>
<type>AE_DFF_LOW</type>
<position>374,259</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3492 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4908</ID>
<type>AA_AND2</type>
<position>417.5,251.5</position>
<input>
<ID>IN_0</ID>3494 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3493 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4909</ID>
<type>BA_TRI_STATE</type>
<position>424.5,251.5</position>
<input>
<ID>ENABLE_0</ID>3493 </input>
<input>
<ID>IN_0</ID>3494 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4910</ID>
<type>AE_DFF_LOW</type>
<position>405,259</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3494 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4911</ID>
<type>AA_AND2</type>
<position>448,251.5</position>
<input>
<ID>IN_0</ID>3496 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4912</ID>
<type>BA_TRI_STATE</type>
<position>455,251.5</position>
<input>
<ID>ENABLE_0</ID>3495 </input>
<input>
<ID>IN_0</ID>3496 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4913</ID>
<type>AE_DFF_LOW</type>
<position>436,259</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3496 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4914</ID>
<type>AA_AND2</type>
<position>479.5,251.5</position>
<input>
<ID>IN_0</ID>3498 </input>
<input>
<ID>IN_1</ID>3434 </input>
<output>
<ID>OUT</ID>3497 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4915</ID>
<type>BA_TRI_STATE</type>
<position>486.5,251.5</position>
<input>
<ID>ENABLE_0</ID>3497 </input>
<input>
<ID>IN_0</ID>3498 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4916</ID>
<type>AE_DFF_LOW</type>
<position>467,259</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3498 </output>
<input>
<ID>clock</ID>3433 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4917</ID>
<type>HA_JUNC_2</type>
<position>339.5,333.5</position>
<input>
<ID>N_in0</ID>3505 </input>
<input>
<ID>N_in1</ID>4104 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4918</ID>
<type>HA_JUNC_2</type>
<position>370.5,333</position>
<input>
<ID>N_in0</ID>3506 </input>
<input>
<ID>N_in1</ID>4106 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4919</ID>
<type>HA_JUNC_2</type>
<position>400.5,333.5</position>
<input>
<ID>N_in0</ID>3507 </input>
<input>
<ID>N_in1</ID>4108 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4920</ID>
<type>HA_JUNC_2</type>
<position>431.5,333.5</position>
<input>
<ID>N_in0</ID>3508 </input>
<input>
<ID>N_in1</ID>4110 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4921</ID>
<type>HA_JUNC_2</type>
<position>462.5,333</position>
<input>
<ID>N_in0</ID>3509 </input>
<input>
<ID>N_in1</ID>4112 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4922</ID>
<type>HA_JUNC_2</type>
<position>274.5,340.5</position>
<input>
<ID>N_in0</ID>3510 </input>
<input>
<ID>N_in1</ID>4098 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4923</ID>
<type>HA_JUNC_2</type>
<position>274.5,183.5</position>
<input>
<ID>N_in0</ID>4126 </input>
<input>
<ID>N_in1</ID>3510 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4924</ID>
<type>HA_JUNC_2</type>
<position>337.5,184.5</position>
<input>
<ID>N_in0</ID>4123 </input>
<input>
<ID>N_in1</ID>3512 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4925</ID>
<type>HA_JUNC_2</type>
<position>368,185</position>
<input>
<ID>N_in0</ID>4121 </input>
<input>
<ID>N_in1</ID>3513 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4926</ID>
<type>HA_JUNC_2</type>
<position>398.5,185</position>
<input>
<ID>N_in0</ID>4119 </input>
<input>
<ID>N_in1</ID>3514 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4927</ID>
<type>HA_JUNC_2</type>
<position>429.5,185</position>
<input>
<ID>N_in0</ID>4118 </input>
<input>
<ID>N_in1</ID>3515 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4928</ID>
<type>HA_JUNC_2</type>
<position>460.5,184.5</position>
<input>
<ID>N_in0</ID>4116 </input>
<input>
<ID>N_in1</ID>3516 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4929</ID>
<type>HA_JUNC_2</type>
<position>491,185</position>
<input>
<ID>N_in0</ID>4114 </input>
<input>
<ID>N_in1</ID>3517 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4930</ID>
<type>HA_JUNC_2</type>
<position>491,342</position>
<input>
<ID>N_in0</ID>3517 </input>
<input>
<ID>N_in1</ID>4113 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4931</ID>
<type>HA_JUNC_2</type>
<position>460.5,341.5</position>
<input>
<ID>N_in0</ID>3516 </input>
<input>
<ID>N_in1</ID>4111 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4932</ID>
<type>HA_JUNC_2</type>
<position>429.5,340.5</position>
<input>
<ID>N_in0</ID>3515 </input>
<input>
<ID>N_in1</ID>4109 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4933</ID>
<type>HA_JUNC_2</type>
<position>398.5,340.5</position>
<input>
<ID>N_in0</ID>3514 </input>
<input>
<ID>N_in1</ID>4107 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4934</ID>
<type>HA_JUNC_2</type>
<position>368,340.5</position>
<input>
<ID>N_in0</ID>3513 </input>
<input>
<ID>N_in1</ID>4105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4935</ID>
<type>HA_JUNC_2</type>
<position>337.5,340.5</position>
<input>
<ID>N_in0</ID>3512 </input>
<input>
<ID>N_in1</ID>4103 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4936</ID>
<type>HA_JUNC_2</type>
<position>305.5,340.5</position>
<input>
<ID>N_in0</ID>3511 </input>
<input>
<ID>N_in1</ID>4101 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>4937</ID>
<type>BE_DECODER_3x8</type>
<position>195.5,268</position>
<input>
<ID>ENABLE</ID>67 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>3525 </output>
<output>
<ID>OUT_1</ID>3524 </output>
<output>
<ID>OUT_2</ID>3523 </output>
<output>
<ID>OUT_3</ID>3522 </output>
<output>
<ID>OUT_4</ID>3521 </output>
<output>
<ID>OUT_5</ID>3520 </output>
<output>
<ID>OUT_6</ID>3519 </output>
<output>
<ID>OUT_7</ID>3518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4938</ID>
<type>BA_TRI_STATE</type>
<position>237.5,253.5</position>
<input>
<ID>ENABLE_0</ID>3522 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4939</ID>
<type>AA_AND2</type>
<position>231.5,258</position>
<input>
<ID>IN_0</ID>3522 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4940</ID>
<type>BA_TRI_STATE</type>
<position>237.5,237.5</position>
<input>
<ID>ENABLE_0</ID>3523 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3436 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4941</ID>
<type>AA_AND2</type>
<position>231.5,242.5</position>
<input>
<ID>IN_0</ID>3523 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4942</ID>
<type>BA_TRI_STATE</type>
<position>237.5,221.5</position>
<input>
<ID>ENABLE_0</ID>3524 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3500 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4943</ID>
<type>AA_AND2</type>
<position>231.5,226.5</position>
<input>
<ID>IN_0</ID>3524 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3499 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4944</ID>
<type>BA_TRI_STATE</type>
<position>237.5,204.5</position>
<input>
<ID>ENABLE_0</ID>3525 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3502 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4945</ID>
<type>AA_AND2</type>
<position>231.5,209.5</position>
<input>
<ID>IN_0</ID>3525 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3501 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4946</ID>
<type>AA_AND2</type>
<position>262.5,268</position>
<input>
<ID>IN_0</ID>3527 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3526 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4947</ID>
<type>BA_TRI_STATE</type>
<position>269.5,268</position>
<input>
<ID>ENABLE_0</ID>3526 </input>
<input>
<ID>IN_0</ID>3527 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4948</ID>
<type>AE_DFF_LOW</type>
<position>250.5,275.5</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3527 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4949</ID>
<type>BA_TRI_STATE</type>
<position>238.5,318.5</position>
<input>
<ID>ENABLE_0</ID>3518 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4950</ID>
<type>AA_AND2</type>
<position>232,323</position>
<input>
<ID>IN_0</ID>3518 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3592 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4951</ID>
<type>BA_TRI_STATE</type>
<position>238.5,302.5</position>
<input>
<ID>ENABLE_0</ID>3519 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3427 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4952</ID>
<type>AA_AND2</type>
<position>294,268</position>
<input>
<ID>IN_0</ID>3529 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4953</ID>
<type>AA_AND2</type>
<position>231.5,307.5</position>
<input>
<ID>IN_0</ID>3519 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4954</ID>
<type>BA_TRI_STATE</type>
<position>301,268</position>
<input>
<ID>ENABLE_0</ID>3528 </input>
<input>
<ID>IN_0</ID>3529 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4955</ID>
<type>BA_TRI_STATE</type>
<position>238.5,286.5</position>
<input>
<ID>ENABLE_0</ID>3520 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3429 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4956</ID>
<type>AE_DFF_LOW</type>
<position>281.5,275.5</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3529 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4957</ID>
<type>AA_AND2</type>
<position>231.5,291.5</position>
<input>
<ID>IN_0</ID>3520 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4958</ID>
<type>AA_AND2</type>
<position>324.5,268</position>
<input>
<ID>IN_0</ID>3531 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3530 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4959</ID>
<type>BA_TRI_STATE</type>
<position>238.5,269.5</position>
<input>
<ID>ENABLE_0</ID>3521 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4960</ID>
<type>BA_TRI_STATE</type>
<position>331.5,268</position>
<input>
<ID>ENABLE_0</ID>3530 </input>
<input>
<ID>IN_0</ID>3531 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4961</ID>
<type>AA_AND2</type>
<position>231.5,274.5</position>
<input>
<ID>IN_0</ID>3521 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4962</ID>
<type>AE_DFF_LOW</type>
<position>312.5,275.5</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3531 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4963</ID>
<type>AA_AND2</type>
<position>356,268</position>
<input>
<ID>IN_0</ID>3533 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4964</ID>
<type>BA_TRI_STATE</type>
<position>363,268</position>
<input>
<ID>ENABLE_0</ID>3532 </input>
<input>
<ID>IN_0</ID>3533 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4965</ID>
<type>AE_DFF_LOW</type>
<position>343.5,275.5</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3533 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4966</ID>
<type>AA_AND2</type>
<position>385.5,268</position>
<input>
<ID>IN_0</ID>3535 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3534 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4967</ID>
<type>BA_TRI_STATE</type>
<position>392.5,268</position>
<input>
<ID>ENABLE_0</ID>3534 </input>
<input>
<ID>IN_0</ID>3535 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4968</ID>
<type>AE_DFF_LOW</type>
<position>373.5,275.5</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3535 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4969</ID>
<type>AA_AND2</type>
<position>417,268</position>
<input>
<ID>IN_0</ID>3537 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3536 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4970</ID>
<type>BA_TRI_STATE</type>
<position>424,268</position>
<input>
<ID>ENABLE_0</ID>3536 </input>
<input>
<ID>IN_0</ID>3537 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4971</ID>
<type>AE_DFF_LOW</type>
<position>404.5,275.5</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3537 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4972</ID>
<type>AA_AND2</type>
<position>447.5,268</position>
<input>
<ID>IN_0</ID>3539 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3538 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4973</ID>
<type>BA_TRI_STATE</type>
<position>454.5,268</position>
<input>
<ID>ENABLE_0</ID>3538 </input>
<input>
<ID>IN_0</ID>3539 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4974</ID>
<type>AE_DFF_LOW</type>
<position>435.5,275.5</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3539 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4975</ID>
<type>AA_AND2</type>
<position>479,268</position>
<input>
<ID>IN_0</ID>3541 </input>
<input>
<ID>IN_1</ID>3432 </input>
<output>
<ID>OUT</ID>3540 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4976</ID>
<type>BA_TRI_STATE</type>
<position>486,268</position>
<input>
<ID>ENABLE_0</ID>3540 </input>
<input>
<ID>IN_0</ID>3541 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4977</ID>
<type>AE_DFF_LOW</type>
<position>466.5,275.5</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3541 </output>
<input>
<ID>clock</ID>3431 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4978</ID>
<type>AA_AND2</type>
<position>263,285</position>
<input>
<ID>IN_0</ID>3543 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3542 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4979</ID>
<type>BA_TRI_STATE</type>
<position>270,285</position>
<input>
<ID>ENABLE_0</ID>3542 </input>
<input>
<ID>IN_0</ID>3543 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4980</ID>
<type>AE_DFF_LOW</type>
<position>251,292.5</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3543 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4981</ID>
<type>AA_AND2</type>
<position>294.5,285</position>
<input>
<ID>IN_0</ID>3545 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3544 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4982</ID>
<type>BA_TRI_STATE</type>
<position>301.5,285</position>
<input>
<ID>ENABLE_0</ID>3544 </input>
<input>
<ID>IN_0</ID>3545 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4983</ID>
<type>AE_DFF_LOW</type>
<position>282,292.5</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3545 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4984</ID>
<type>AA_AND2</type>
<position>325,285</position>
<input>
<ID>IN_0</ID>3547 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4985</ID>
<type>BA_TRI_STATE</type>
<position>332,285</position>
<input>
<ID>ENABLE_0</ID>3546 </input>
<input>
<ID>IN_0</ID>3547 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4986</ID>
<type>AE_DFF_LOW</type>
<position>313,292.5</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3547 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4987</ID>
<type>AA_AND2</type>
<position>356.5,285</position>
<input>
<ID>IN_0</ID>3549 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3548 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4988</ID>
<type>BA_TRI_STATE</type>
<position>363.5,285</position>
<input>
<ID>ENABLE_0</ID>3548 </input>
<input>
<ID>IN_0</ID>3549 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4989</ID>
<type>AE_DFF_LOW</type>
<position>344,292.5</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3549 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4990</ID>
<type>AA_AND2</type>
<position>386,285</position>
<input>
<ID>IN_0</ID>3551 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3550 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4991</ID>
<type>BA_TRI_STATE</type>
<position>393,285</position>
<input>
<ID>ENABLE_0</ID>3550 </input>
<input>
<ID>IN_0</ID>3551 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4992</ID>
<type>AE_DFF_LOW</type>
<position>374,292.5</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3551 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4993</ID>
<type>AA_AND2</type>
<position>417.5,285</position>
<input>
<ID>IN_0</ID>3553 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3552 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4994</ID>
<type>BA_TRI_STATE</type>
<position>424.5,285</position>
<input>
<ID>ENABLE_0</ID>3552 </input>
<input>
<ID>IN_0</ID>3553 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4995</ID>
<type>AE_DFF_LOW</type>
<position>405,292.5</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3553 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4996</ID>
<type>AA_AND2</type>
<position>448,285</position>
<input>
<ID>IN_0</ID>3555 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3554 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4997</ID>
<type>BA_TRI_STATE</type>
<position>455,285</position>
<input>
<ID>ENABLE_0</ID>3554 </input>
<input>
<ID>IN_0</ID>3555 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4998</ID>
<type>AE_DFF_LOW</type>
<position>436,292.5</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3555 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4999</ID>
<type>AA_AND2</type>
<position>479.5,285</position>
<input>
<ID>IN_0</ID>3557 </input>
<input>
<ID>IN_1</ID>3429 </input>
<output>
<ID>OUT</ID>3556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5000</ID>
<type>BA_TRI_STATE</type>
<position>486.5,285</position>
<input>
<ID>ENABLE_0</ID>3556 </input>
<input>
<ID>IN_0</ID>3557 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5001</ID>
<type>AE_DFF_LOW</type>
<position>467,292.5</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3557 </output>
<input>
<ID>clock</ID>3430 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5002</ID>
<type>AA_AND2</type>
<position>263.5,301</position>
<input>
<ID>IN_0</ID>3559 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3558 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5003</ID>
<type>BA_TRI_STATE</type>
<position>270.5,301</position>
<input>
<ID>ENABLE_0</ID>3558 </input>
<input>
<ID>IN_0</ID>3559 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5004</ID>
<type>AE_DFF_LOW</type>
<position>251.5,308.5</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3559 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5005</ID>
<type>AA_AND2</type>
<position>295,301</position>
<input>
<ID>IN_0</ID>3561 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3560 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5006</ID>
<type>BA_TRI_STATE</type>
<position>302,301</position>
<input>
<ID>ENABLE_0</ID>3560 </input>
<input>
<ID>IN_0</ID>3561 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5007</ID>
<type>AE_DFF_LOW</type>
<position>282.5,308.5</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3561 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5008</ID>
<type>AA_AND2</type>
<position>325.5,301</position>
<input>
<ID>IN_0</ID>3563 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3562 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5009</ID>
<type>BA_TRI_STATE</type>
<position>332.5,301</position>
<input>
<ID>ENABLE_0</ID>3562 </input>
<input>
<ID>IN_0</ID>3563 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5010</ID>
<type>AE_DFF_LOW</type>
<position>313.5,308.5</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3563 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5011</ID>
<type>AA_AND2</type>
<position>357,301</position>
<input>
<ID>IN_0</ID>3565 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5012</ID>
<type>BA_TRI_STATE</type>
<position>364,301</position>
<input>
<ID>ENABLE_0</ID>3564 </input>
<input>
<ID>IN_0</ID>3565 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5013</ID>
<type>AE_DFF_LOW</type>
<position>344.5,308.5</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3565 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5014</ID>
<type>AA_AND2</type>
<position>386.5,301</position>
<input>
<ID>IN_0</ID>3567 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3566 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5015</ID>
<type>BA_TRI_STATE</type>
<position>393.5,301</position>
<input>
<ID>ENABLE_0</ID>3566 </input>
<input>
<ID>IN_0</ID>3567 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5016</ID>
<type>AE_DFF_LOW</type>
<position>374.5,308.5</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3567 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5017</ID>
<type>AA_AND2</type>
<position>418,301</position>
<input>
<ID>IN_0</ID>3569 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3568 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5018</ID>
<type>BA_TRI_STATE</type>
<position>425,301</position>
<input>
<ID>ENABLE_0</ID>3568 </input>
<input>
<ID>IN_0</ID>3569 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5019</ID>
<type>AE_DFF_LOW</type>
<position>405.5,308.5</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3569 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5020</ID>
<type>AA_AND2</type>
<position>448.5,301</position>
<input>
<ID>IN_0</ID>3571 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3570 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5021</ID>
<type>BA_TRI_STATE</type>
<position>455.5,301</position>
<input>
<ID>ENABLE_0</ID>3570 </input>
<input>
<ID>IN_0</ID>3571 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5022</ID>
<type>AE_DFF_LOW</type>
<position>436.5,308.5</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3571 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5023</ID>
<type>AA_AND2</type>
<position>480,301</position>
<input>
<ID>IN_0</ID>3573 </input>
<input>
<ID>IN_1</ID>3427 </input>
<output>
<ID>OUT</ID>3572 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5024</ID>
<type>BA_TRI_STATE</type>
<position>487,301</position>
<input>
<ID>ENABLE_0</ID>3572 </input>
<input>
<ID>IN_0</ID>3573 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5025</ID>
<type>AE_DFF_LOW</type>
<position>467.5,308.5</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3573 </output>
<input>
<ID>clock</ID>3428 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5026</ID>
<type>AA_AND2</type>
<position>264,316.5</position>
<input>
<ID>IN_0</ID>3575 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3574 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5027</ID>
<type>BA_TRI_STATE</type>
<position>271,316.5</position>
<input>
<ID>ENABLE_0</ID>3574 </input>
<input>
<ID>IN_0</ID>3575 </input>
<output>
<ID>OUT_0</ID>3510 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5028</ID>
<type>AE_DFF_LOW</type>
<position>252,324</position>
<input>
<ID>IN_0</ID>3590 </input>
<output>
<ID>OUT_0</ID>3575 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5029</ID>
<type>AA_AND2</type>
<position>295.5,316.5</position>
<input>
<ID>IN_0</ID>3577 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3576 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5030</ID>
<type>BA_TRI_STATE</type>
<position>302.5,316.5</position>
<input>
<ID>ENABLE_0</ID>3576 </input>
<input>
<ID>IN_0</ID>3577 </input>
<output>
<ID>OUT_0</ID>3511 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5031</ID>
<type>AE_DFF_LOW</type>
<position>283,324</position>
<input>
<ID>IN_0</ID>3503 </input>
<output>
<ID>OUT_0</ID>3577 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5032</ID>
<type>AA_AND2</type>
<position>326,316.5</position>
<input>
<ID>IN_0</ID>3579 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3578 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5033</ID>
<type>BA_TRI_STATE</type>
<position>333,316.5</position>
<input>
<ID>ENABLE_0</ID>3578 </input>
<input>
<ID>IN_0</ID>3579 </input>
<output>
<ID>OUT_0</ID>3512 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5034</ID>
<type>AE_DFF_LOW</type>
<position>314,324</position>
<input>
<ID>IN_0</ID>3504 </input>
<output>
<ID>OUT_0</ID>3579 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5035</ID>
<type>AA_AND2</type>
<position>357.5,316.5</position>
<input>
<ID>IN_0</ID>3581 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5036</ID>
<type>BA_TRI_STATE</type>
<position>364.5,316.5</position>
<input>
<ID>ENABLE_0</ID>3580 </input>
<input>
<ID>IN_0</ID>3581 </input>
<output>
<ID>OUT_0</ID>3513 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5037</ID>
<type>AE_DFF_LOW</type>
<position>345,324</position>
<input>
<ID>IN_0</ID>3505 </input>
<output>
<ID>OUT_0</ID>3581 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5038</ID>
<type>AA_AND2</type>
<position>387,316.5</position>
<input>
<ID>IN_0</ID>3583 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3582 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5039</ID>
<type>BA_TRI_STATE</type>
<position>394,316.5</position>
<input>
<ID>ENABLE_0</ID>3582 </input>
<input>
<ID>IN_0</ID>3583 </input>
<output>
<ID>OUT_0</ID>3514 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5040</ID>
<type>AE_DFF_LOW</type>
<position>375,324</position>
<input>
<ID>IN_0</ID>3506 </input>
<output>
<ID>OUT_0</ID>3583 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5041</ID>
<type>AA_AND2</type>
<position>418.5,316.5</position>
<input>
<ID>IN_0</ID>3585 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5042</ID>
<type>BA_TRI_STATE</type>
<position>425.5,316.5</position>
<input>
<ID>ENABLE_0</ID>3584 </input>
<input>
<ID>IN_0</ID>3585 </input>
<output>
<ID>OUT_0</ID>3515 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5043</ID>
<type>AE_DFF_LOW</type>
<position>406,324</position>
<input>
<ID>IN_0</ID>3507 </input>
<output>
<ID>OUT_0</ID>3585 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5044</ID>
<type>AA_AND2</type>
<position>449,316.5</position>
<input>
<ID>IN_0</ID>3587 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5045</ID>
<type>BA_TRI_STATE</type>
<position>456,316.5</position>
<input>
<ID>ENABLE_0</ID>3586 </input>
<input>
<ID>IN_0</ID>3587 </input>
<output>
<ID>OUT_0</ID>3516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5046</ID>
<type>AE_DFF_LOW</type>
<position>437,324</position>
<input>
<ID>IN_0</ID>3508 </input>
<output>
<ID>OUT_0</ID>3587 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5047</ID>
<type>AA_AND2</type>
<position>480.5,316.5</position>
<input>
<ID>IN_0</ID>3589 </input>
<input>
<ID>IN_1</ID>3591 </input>
<output>
<ID>OUT</ID>3588 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5048</ID>
<type>BA_TRI_STATE</type>
<position>487.5,316.5</position>
<input>
<ID>ENABLE_0</ID>3588 </input>
<input>
<ID>IN_0</ID>3589 </input>
<output>
<ID>OUT_0</ID>3517 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5049</ID>
<type>AE_DFF_LOW</type>
<position>468,324</position>
<input>
<ID>IN_0</ID>3509 </input>
<output>
<ID>OUT_0</ID>3589 </output>
<input>
<ID>clock</ID>3592 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2170</ID>
<type>AA_AND2</type>
<position>265.5,-182</position>
<input>
<ID>IN_0</ID>1578 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1577 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2171</ID>
<type>BA_TRI_STATE</type>
<position>272.5,-182</position>
<input>
<ID>ENABLE_0</ID>1577 </input>
<input>
<ID>IN_0</ID>1578 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2172</ID>
<type>AE_DFF_LOW</type>
<position>253.5,-174.5</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1578 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2173</ID>
<type>HA_JUNC_2</type>
<position>249.5,-193</position>
<input>
<ID>N_in0</ID>4161 </input>
<input>
<ID>N_in1</ID>1742 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2174</ID>
<type>HA_JUNC_2</type>
<position>280.5,-193.5</position>
<input>
<ID>N_in0</ID>4160 </input>
<input>
<ID>N_in1</ID>1655 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2175</ID>
<type>HA_JUNC_2</type>
<position>312.5,-193.5</position>
<input>
<ID>N_in0</ID>4158 </input>
<input>
<ID>N_in1</ID>1656 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2176</ID>
<type>HA_JUNC_2</type>
<position>343.5,-192.5</position>
<input>
<ID>N_in0</ID>4156 </input>
<input>
<ID>N_in1</ID>1657 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2177</ID>
<type>HA_JUNC_2</type>
<position>373.5,-191.5</position>
<input>
<ID>N_in0</ID>4154 </input>
<input>
<ID>N_in1</ID>1658 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2178</ID>
<type>HA_JUNC_2</type>
<position>404.5,-191</position>
<input>
<ID>N_in0</ID>4151 </input>
<input>
<ID>N_in1</ID>1659 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2179</ID>
<type>HA_JUNC_2</type>
<position>466.5,-192</position>
<input>
<ID>N_in0</ID>4147 </input>
<input>
<ID>N_in1</ID>1661 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2180</ID>
<type>HA_JUNC_2</type>
<position>435.5,-190</position>
<input>
<ID>N_in0</ID>4149 </input>
<input>
<ID>N_in1</ID>1660 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2181</ID>
<type>HA_JUNC_2</type>
<position>249.5,-51.5</position>
<input>
<ID>N_in0</ID>1742 </input>
<input>
<ID>N_in1</ID>4130 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2182</ID>
<type>HA_JUNC_2</type>
<position>280.5,-51.5</position>
<input>
<ID>N_in0</ID>1655 </input>
<input>
<ID>N_in1</ID>4132 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2183</ID>
<type>HA_JUNC_2</type>
<position>312.5,-51.5</position>
<input>
<ID>N_in0</ID>1656 </input>
<input>
<ID>N_in1</ID>4134 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2184</ID>
<type>AA_AND2</type>
<position>297,-182</position>
<input>
<ID>IN_0</ID>1590 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1589 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2185</ID>
<type>BA_TRI_STATE</type>
<position>304,-182</position>
<input>
<ID>ENABLE_0</ID>1589 </input>
<input>
<ID>IN_0</ID>1590 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2186</ID>
<type>AE_DFF_LOW</type>
<position>284.5,-174.5</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1590 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2187</ID>
<type>AA_AND2</type>
<position>327.5,-182</position>
<input>
<ID>IN_0</ID>1592 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2188</ID>
<type>BA_TRI_STATE</type>
<position>334.5,-182</position>
<input>
<ID>ENABLE_0</ID>1591 </input>
<input>
<ID>IN_0</ID>1592 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2189</ID>
<type>AE_DFF_LOW</type>
<position>315.5,-174.5</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1592 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2190</ID>
<type>AA_AND2</type>
<position>359,-182</position>
<input>
<ID>IN_0</ID>1594 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2191</ID>
<type>BA_TRI_STATE</type>
<position>366,-182</position>
<input>
<ID>ENABLE_0</ID>1593 </input>
<input>
<ID>IN_0</ID>1594 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2192</ID>
<type>AE_DFF_LOW</type>
<position>346.5,-174.5</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1594 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2193</ID>
<type>AA_AND2</type>
<position>388.5,-182</position>
<input>
<ID>IN_0</ID>1596 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2194</ID>
<type>BA_TRI_STATE</type>
<position>395.5,-182</position>
<input>
<ID>ENABLE_0</ID>1595 </input>
<input>
<ID>IN_0</ID>1596 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2195</ID>
<type>AE_DFF_LOW</type>
<position>376.5,-174.5</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1596 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2196</ID>
<type>AA_AND2</type>
<position>420,-182</position>
<input>
<ID>IN_0</ID>1598 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2197</ID>
<type>BA_TRI_STATE</type>
<position>427,-182</position>
<input>
<ID>ENABLE_0</ID>1597 </input>
<input>
<ID>IN_0</ID>1598 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2198</ID>
<type>AE_DFF_LOW</type>
<position>407.5,-174.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1598 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2199</ID>
<type>AA_AND2</type>
<position>450.5,-182</position>
<input>
<ID>IN_0</ID>1600 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2200</ID>
<type>BA_TRI_STATE</type>
<position>457.5,-182</position>
<input>
<ID>ENABLE_0</ID>1599 </input>
<input>
<ID>IN_0</ID>1600 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2201</ID>
<type>AE_DFF_LOW</type>
<position>438.5,-174.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1600 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2202</ID>
<type>AA_AND2</type>
<position>482,-182</position>
<input>
<ID>IN_0</ID>1602 </input>
<input>
<ID>IN_1</ID>1654 </input>
<output>
<ID>OUT</ID>1601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2203</ID>
<type>BA_TRI_STATE</type>
<position>489,-182</position>
<input>
<ID>ENABLE_0</ID>1601 </input>
<input>
<ID>IN_0</ID>1602 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2204</ID>
<type>AE_DFF_LOW</type>
<position>469.5,-174.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1602 </output>
<input>
<ID>clock</ID>1653 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2205</ID>
<type>AA_AND2</type>
<position>266,-165</position>
<input>
<ID>IN_0</ID>1604 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1603 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2206</ID>
<type>BA_TRI_STATE</type>
<position>273,-165</position>
<input>
<ID>ENABLE_0</ID>1603 </input>
<input>
<ID>IN_0</ID>1604 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2207</ID>
<type>AE_DFF_LOW</type>
<position>254,-157.5</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1604 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2208</ID>
<type>AA_AND2</type>
<position>297.5,-165</position>
<input>
<ID>IN_0</ID>1606 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1605 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2209</ID>
<type>BA_TRI_STATE</type>
<position>304.5,-165</position>
<input>
<ID>ENABLE_0</ID>1605 </input>
<input>
<ID>IN_0</ID>1606 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2210</ID>
<type>AE_DFF_LOW</type>
<position>285,-157.5</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1606 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2211</ID>
<type>AA_AND2</type>
<position>328,-165</position>
<input>
<ID>IN_0</ID>1608 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1607 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5290</ID>
<type>AA_AND2</type>
<position>257.5,-891</position>
<input>
<ID>IN_0</ID>3762 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3761 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2212</ID>
<type>BA_TRI_STATE</type>
<position>335,-165</position>
<input>
<ID>ENABLE_0</ID>1607 </input>
<input>
<ID>IN_0</ID>1608 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5291</ID>
<type>BA_TRI_STATE</type>
<position>264.5,-891</position>
<input>
<ID>ENABLE_0</ID>3761 </input>
<input>
<ID>IN_0</ID>3762 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2213</ID>
<type>AE_DFF_LOW</type>
<position>316,-157.5</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1608 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5292</ID>
<type>AE_DFF_LOW</type>
<position>245.5,-883.5</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3762 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2214</ID>
<type>AA_AND2</type>
<position>359.5,-165</position>
<input>
<ID>IN_0</ID>1610 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1609 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5293</ID>
<type>HA_JUNC_2</type>
<position>241.5,-902</position>
<input>
<ID>N_in0</ID>20 </input>
<input>
<ID>N_in1</ID>3926 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2215</ID>
<type>BA_TRI_STATE</type>
<position>366.5,-165</position>
<input>
<ID>ENABLE_0</ID>1609 </input>
<input>
<ID>IN_0</ID>1610 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5294</ID>
<type>HA_JUNC_2</type>
<position>272.5,-902.5</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>3839 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2216</ID>
<type>AE_DFF_LOW</type>
<position>347,-157.5</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1610 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5295</ID>
<type>HA_JUNC_2</type>
<position>304.5,-902.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>3840 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2217</ID>
<type>AA_AND2</type>
<position>389,-165</position>
<input>
<ID>IN_0</ID>1612 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5296</ID>
<type>HA_JUNC_2</type>
<position>335.5,-901.5</position>
<input>
<ID>N_in0</ID>23 </input>
<input>
<ID>N_in1</ID>3841 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2218</ID>
<type>BA_TRI_STATE</type>
<position>396,-165</position>
<input>
<ID>ENABLE_0</ID>1611 </input>
<input>
<ID>IN_0</ID>1612 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5297</ID>
<type>HA_JUNC_2</type>
<position>365.5,-900.5</position>
<input>
<ID>N_in0</ID>24 </input>
<input>
<ID>N_in1</ID>3842 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2219</ID>
<type>AE_DFF_LOW</type>
<position>377,-157.5</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1612 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5298</ID>
<type>HA_JUNC_2</type>
<position>396.5,-900</position>
<input>
<ID>N_in0</ID>25 </input>
<input>
<ID>N_in1</ID>3843 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2220</ID>
<type>AA_AND2</type>
<position>420.5,-165</position>
<input>
<ID>IN_0</ID>1614 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1613 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5299</ID>
<type>HA_JUNC_2</type>
<position>458.5,-901</position>
<input>
<ID>N_in0</ID>27 </input>
<input>
<ID>N_in1</ID>3845 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2221</ID>
<type>BA_TRI_STATE</type>
<position>427.5,-165</position>
<input>
<ID>ENABLE_0</ID>1613 </input>
<input>
<ID>IN_0</ID>1614 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5300</ID>
<type>HA_JUNC_2</type>
<position>427.5,-899</position>
<input>
<ID>N_in0</ID>26 </input>
<input>
<ID>N_in1</ID>3844 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2222</ID>
<type>AE_DFF_LOW</type>
<position>408,-157.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1614 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5301</ID>
<type>HA_JUNC_2</type>
<position>241.5,-760.5</position>
<input>
<ID>N_in0</ID>3926 </input>
<input>
<ID>N_in1</ID>4209 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2223</ID>
<type>AA_AND2</type>
<position>451,-165</position>
<input>
<ID>IN_0</ID>1616 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1615 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5302</ID>
<type>HA_JUNC_2</type>
<position>272.5,-760.5</position>
<input>
<ID>N_in0</ID>3839 </input>
<input>
<ID>N_in1</ID>4208 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2224</ID>
<type>BA_TRI_STATE</type>
<position>458,-165</position>
<input>
<ID>ENABLE_0</ID>1615 </input>
<input>
<ID>IN_0</ID>1616 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5303</ID>
<type>HA_JUNC_2</type>
<position>304.5,-760.5</position>
<input>
<ID>N_in0</ID>3840 </input>
<input>
<ID>N_in1</ID>4205 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2225</ID>
<type>AE_DFF_LOW</type>
<position>439,-157.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1616 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5304</ID>
<type>AA_AND2</type>
<position>289,-891</position>
<input>
<ID>IN_0</ID>3774 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3773 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2226</ID>
<type>AA_AND2</type>
<position>482.5,-165</position>
<input>
<ID>IN_0</ID>1618 </input>
<input>
<ID>IN_1</ID>1652 </input>
<output>
<ID>OUT</ID>1617 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5305</ID>
<type>BA_TRI_STATE</type>
<position>296,-891</position>
<input>
<ID>ENABLE_0</ID>3773 </input>
<input>
<ID>IN_0</ID>3774 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2227</ID>
<type>BA_TRI_STATE</type>
<position>489.5,-165</position>
<input>
<ID>ENABLE_0</ID>1617 </input>
<input>
<ID>IN_0</ID>1618 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5306</ID>
<type>AE_DFF_LOW</type>
<position>276.5,-883.5</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3774 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2228</ID>
<type>AE_DFF_LOW</type>
<position>470,-157.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1618 </output>
<input>
<ID>clock</ID>1651 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5307</ID>
<type>AA_AND2</type>
<position>319.5,-891</position>
<input>
<ID>IN_0</ID>3776 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2229</ID>
<type>AA_AND2</type>
<position>266.5,-149</position>
<input>
<ID>IN_0</ID>1620 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1619 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5308</ID>
<type>BA_TRI_STATE</type>
<position>326.5,-891</position>
<input>
<ID>ENABLE_0</ID>3775 </input>
<input>
<ID>IN_0</ID>3776 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2230</ID>
<type>BA_TRI_STATE</type>
<position>273.5,-149</position>
<input>
<ID>ENABLE_0</ID>1619 </input>
<input>
<ID>IN_0</ID>1620 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5309</ID>
<type>AE_DFF_LOW</type>
<position>307.5,-883.5</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3776 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2231</ID>
<type>AE_DFF_LOW</type>
<position>254.5,-141.5</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1620 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5310</ID>
<type>AA_AND2</type>
<position>351,-891</position>
<input>
<ID>IN_0</ID>3778 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3777 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2232</ID>
<type>AA_AND2</type>
<position>298,-149</position>
<input>
<ID>IN_0</ID>1622 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1621 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5311</ID>
<type>BA_TRI_STATE</type>
<position>358,-891</position>
<input>
<ID>ENABLE_0</ID>3777 </input>
<input>
<ID>IN_0</ID>3778 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2233</ID>
<type>BA_TRI_STATE</type>
<position>305,-149</position>
<input>
<ID>ENABLE_0</ID>1621 </input>
<input>
<ID>IN_0</ID>1622 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5312</ID>
<type>AE_DFF_LOW</type>
<position>338.5,-883.5</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3778 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2234</ID>
<type>AE_DFF_LOW</type>
<position>285.5,-141.5</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1622 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5313</ID>
<type>AA_AND2</type>
<position>380.5,-891</position>
<input>
<ID>IN_0</ID>3780 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3779 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2235</ID>
<type>AA_AND2</type>
<position>328.5,-149</position>
<input>
<ID>IN_0</ID>1624 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1623 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5314</ID>
<type>BA_TRI_STATE</type>
<position>387.5,-891</position>
<input>
<ID>ENABLE_0</ID>3779 </input>
<input>
<ID>IN_0</ID>3780 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2236</ID>
<type>BA_TRI_STATE</type>
<position>335.5,-149</position>
<input>
<ID>ENABLE_0</ID>1623 </input>
<input>
<ID>IN_0</ID>1624 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5315</ID>
<type>AE_DFF_LOW</type>
<position>368.5,-883.5</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3780 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2237</ID>
<type>AE_DFF_LOW</type>
<position>316.5,-141.5</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1624 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5316</ID>
<type>AA_AND2</type>
<position>412,-891</position>
<input>
<ID>IN_0</ID>3782 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2238</ID>
<type>AA_AND2</type>
<position>360,-149</position>
<input>
<ID>IN_0</ID>1626 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5317</ID>
<type>BA_TRI_STATE</type>
<position>419,-891</position>
<input>
<ID>ENABLE_0</ID>3781 </input>
<input>
<ID>IN_0</ID>3782 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2239</ID>
<type>BA_TRI_STATE</type>
<position>367,-149</position>
<input>
<ID>ENABLE_0</ID>1625 </input>
<input>
<ID>IN_0</ID>1626 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5318</ID>
<type>AE_DFF_LOW</type>
<position>399.5,-883.5</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3782 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2240</ID>
<type>AE_DFF_LOW</type>
<position>347.5,-141.5</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1626 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5319</ID>
<type>AA_AND2</type>
<position>442.5,-891</position>
<input>
<ID>IN_0</ID>3784 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2241</ID>
<type>AA_AND2</type>
<position>389.5,-149</position>
<input>
<ID>IN_0</ID>1628 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5320</ID>
<type>BA_TRI_STATE</type>
<position>449.5,-891</position>
<input>
<ID>ENABLE_0</ID>3783 </input>
<input>
<ID>IN_0</ID>3784 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2242</ID>
<type>BA_TRI_STATE</type>
<position>396.5,-149</position>
<input>
<ID>ENABLE_0</ID>1627 </input>
<input>
<ID>IN_0</ID>1628 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5321</ID>
<type>AE_DFF_LOW</type>
<position>430.5,-883.5</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3784 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2243</ID>
<type>AE_DFF_LOW</type>
<position>377.5,-141.5</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1628 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5322</ID>
<type>AA_AND2</type>
<position>474,-891</position>
<input>
<ID>IN_0</ID>3786 </input>
<input>
<ID>IN_1</ID>3838 </input>
<output>
<ID>OUT</ID>3785 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2244</ID>
<type>AA_AND2</type>
<position>421,-149</position>
<input>
<ID>IN_0</ID>1630 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1629 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5323</ID>
<type>BA_TRI_STATE</type>
<position>481,-891</position>
<input>
<ID>ENABLE_0</ID>3785 </input>
<input>
<ID>IN_0</ID>3786 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2245</ID>
<type>BA_TRI_STATE</type>
<position>428,-149</position>
<input>
<ID>ENABLE_0</ID>1629 </input>
<input>
<ID>IN_0</ID>1630 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5324</ID>
<type>AE_DFF_LOW</type>
<position>461.5,-883.5</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3786 </output>
<input>
<ID>clock</ID>3837 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2246</ID>
<type>AE_DFF_LOW</type>
<position>408.5,-141.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1630 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5325</ID>
<type>AA_AND2</type>
<position>258,-874</position>
<input>
<ID>IN_0</ID>3788 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3787 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2247</ID>
<type>AA_AND2</type>
<position>451.5,-149</position>
<input>
<ID>IN_0</ID>1632 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1631 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5326</ID>
<type>BA_TRI_STATE</type>
<position>265,-874</position>
<input>
<ID>ENABLE_0</ID>3787 </input>
<input>
<ID>IN_0</ID>3788 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2248</ID>
<type>BA_TRI_STATE</type>
<position>458.5,-149</position>
<input>
<ID>ENABLE_0</ID>1631 </input>
<input>
<ID>IN_0</ID>1632 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5327</ID>
<type>AE_DFF_LOW</type>
<position>246,-866.5</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3788 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2249</ID>
<type>AE_DFF_LOW</type>
<position>439.5,-141.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1632 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5328</ID>
<type>AA_AND2</type>
<position>289.5,-874</position>
<input>
<ID>IN_0</ID>3790 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3789 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2250</ID>
<type>AA_AND2</type>
<position>483,-149</position>
<input>
<ID>IN_0</ID>1634 </input>
<input>
<ID>IN_1</ID>1588 </input>
<output>
<ID>OUT</ID>1633 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5329</ID>
<type>BA_TRI_STATE</type>
<position>296.5,-874</position>
<input>
<ID>ENABLE_0</ID>3789 </input>
<input>
<ID>IN_0</ID>3790 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2251</ID>
<type>BA_TRI_STATE</type>
<position>490,-149</position>
<input>
<ID>ENABLE_0</ID>1633 </input>
<input>
<ID>IN_0</ID>1634 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5330</ID>
<type>AE_DFF_LOW</type>
<position>277,-866.5</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3790 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2252</ID>
<type>AE_DFF_LOW</type>
<position>470.5,-141.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1634 </output>
<input>
<ID>clock</ID>1587 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5331</ID>
<type>AA_AND2</type>
<position>320,-874</position>
<input>
<ID>IN_0</ID>3792 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3791 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2253</ID>
<type>AA_AND2</type>
<position>267,-133.5</position>
<input>
<ID>IN_0</ID>1636 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1635 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5332</ID>
<type>BA_TRI_STATE</type>
<position>327,-874</position>
<input>
<ID>ENABLE_0</ID>3791 </input>
<input>
<ID>IN_0</ID>3792 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2254</ID>
<type>BA_TRI_STATE</type>
<position>274,-133.5</position>
<input>
<ID>ENABLE_0</ID>1635 </input>
<input>
<ID>IN_0</ID>1636 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5333</ID>
<type>AE_DFF_LOW</type>
<position>308,-866.5</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3792 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2255</ID>
<type>AE_DFF_LOW</type>
<position>255,-126</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1636 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5334</ID>
<type>AA_AND2</type>
<position>351.5,-874</position>
<input>
<ID>IN_0</ID>3794 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2256</ID>
<type>AA_AND2</type>
<position>298.5,-133.5</position>
<input>
<ID>IN_0</ID>1638 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1637 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5335</ID>
<type>BA_TRI_STATE</type>
<position>358.5,-874</position>
<input>
<ID>ENABLE_0</ID>3793 </input>
<input>
<ID>IN_0</ID>3794 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2257</ID>
<type>BA_TRI_STATE</type>
<position>305.5,-133.5</position>
<input>
<ID>ENABLE_0</ID>1637 </input>
<input>
<ID>IN_0</ID>1638 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5336</ID>
<type>AE_DFF_LOW</type>
<position>339,-866.5</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3794 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2258</ID>
<type>AE_DFF_LOW</type>
<position>286,-126</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1638 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5337</ID>
<type>AA_AND2</type>
<position>381,-874</position>
<input>
<ID>IN_0</ID>3796 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3795 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2259</ID>
<type>AA_AND2</type>
<position>329,-133.5</position>
<input>
<ID>IN_0</ID>1640 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1639 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5338</ID>
<type>BA_TRI_STATE</type>
<position>388,-874</position>
<input>
<ID>ENABLE_0</ID>3795 </input>
<input>
<ID>IN_0</ID>3796 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2260</ID>
<type>BA_TRI_STATE</type>
<position>336,-133.5</position>
<input>
<ID>ENABLE_0</ID>1639 </input>
<input>
<ID>IN_0</ID>1640 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5339</ID>
<type>AE_DFF_LOW</type>
<position>369,-866.5</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3796 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2261</ID>
<type>AE_DFF_LOW</type>
<position>317,-126</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1640 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5340</ID>
<type>AA_AND2</type>
<position>412.5,-874</position>
<input>
<ID>IN_0</ID>3798 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3797 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2262</ID>
<type>AA_AND2</type>
<position>360.5,-133.5</position>
<input>
<ID>IN_0</ID>1642 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5341</ID>
<type>BA_TRI_STATE</type>
<position>419.5,-874</position>
<input>
<ID>ENABLE_0</ID>3797 </input>
<input>
<ID>IN_0</ID>3798 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2263</ID>
<type>BA_TRI_STATE</type>
<position>367.5,-133.5</position>
<input>
<ID>ENABLE_0</ID>1641 </input>
<input>
<ID>IN_0</ID>1642 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5342</ID>
<type>AE_DFF_LOW</type>
<position>400,-866.5</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3798 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2264</ID>
<type>AE_DFF_LOW</type>
<position>348,-126</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1642 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5343</ID>
<type>AA_AND2</type>
<position>443,-874</position>
<input>
<ID>IN_0</ID>3800 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3799 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2265</ID>
<type>AA_AND2</type>
<position>390,-133.5</position>
<input>
<ID>IN_0</ID>1644 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1643 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5344</ID>
<type>BA_TRI_STATE</type>
<position>450,-874</position>
<input>
<ID>ENABLE_0</ID>3799 </input>
<input>
<ID>IN_0</ID>3800 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2266</ID>
<type>BA_TRI_STATE</type>
<position>397,-133.5</position>
<input>
<ID>ENABLE_0</ID>1643 </input>
<input>
<ID>IN_0</ID>1644 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5345</ID>
<type>AE_DFF_LOW</type>
<position>431,-866.5</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3800 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2267</ID>
<type>AE_DFF_LOW</type>
<position>378,-126</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1644 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5346</ID>
<type>AA_AND2</type>
<position>474.5,-874</position>
<input>
<ID>IN_0</ID>3802 </input>
<input>
<ID>IN_1</ID>3836 </input>
<output>
<ID>OUT</ID>3801 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2268</ID>
<type>AA_AND2</type>
<position>421.5,-133.5</position>
<input>
<ID>IN_0</ID>1646 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5347</ID>
<type>BA_TRI_STATE</type>
<position>481.5,-874</position>
<input>
<ID>ENABLE_0</ID>3801 </input>
<input>
<ID>IN_0</ID>3802 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2269</ID>
<type>BA_TRI_STATE</type>
<position>428.5,-133.5</position>
<input>
<ID>ENABLE_0</ID>1645 </input>
<input>
<ID>IN_0</ID>1646 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5348</ID>
<type>AE_DFF_LOW</type>
<position>462,-866.5</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3802 </output>
<input>
<ID>clock</ID>3835 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2270</ID>
<type>AE_DFF_LOW</type>
<position>409,-126</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1646 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5349</ID>
<type>AA_AND2</type>
<position>258.5,-858</position>
<input>
<ID>IN_0</ID>3804 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3803 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2271</ID>
<type>AA_AND2</type>
<position>452,-133.5</position>
<input>
<ID>IN_0</ID>1648 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1647 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5350</ID>
<type>BA_TRI_STATE</type>
<position>265.5,-858</position>
<input>
<ID>ENABLE_0</ID>3803 </input>
<input>
<ID>IN_0</ID>3804 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2272</ID>
<type>BA_TRI_STATE</type>
<position>459,-133.5</position>
<input>
<ID>ENABLE_0</ID>1647 </input>
<input>
<ID>IN_0</ID>1648 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5351</ID>
<type>AE_DFF_LOW</type>
<position>246.5,-850.5</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3804 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2273</ID>
<type>AE_DFF_LOW</type>
<position>440,-126</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1648 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5352</ID>
<type>AA_AND2</type>
<position>290,-858</position>
<input>
<ID>IN_0</ID>3806 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3805 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2274</ID>
<type>AA_AND2</type>
<position>483.5,-133.5</position>
<input>
<ID>IN_0</ID>1650 </input>
<input>
<ID>IN_1</ID>1586 </input>
<output>
<ID>OUT</ID>1649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5353</ID>
<type>BA_TRI_STATE</type>
<position>297,-858</position>
<input>
<ID>ENABLE_0</ID>3805 </input>
<input>
<ID>IN_0</ID>3806 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2275</ID>
<type>BA_TRI_STATE</type>
<position>490.5,-133.5</position>
<input>
<ID>ENABLE_0</ID>1649 </input>
<input>
<ID>IN_0</ID>1650 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5354</ID>
<type>AE_DFF_LOW</type>
<position>277.5,-850.5</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3806 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2276</ID>
<type>AE_DFF_LOW</type>
<position>471,-126</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1650 </output>
<input>
<ID>clock</ID>1585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5355</ID>
<type>AA_AND2</type>
<position>320.5,-858</position>
<input>
<ID>IN_0</ID>3808 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3807 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2277</ID>
<type>HA_JUNC_2</type>
<position>343.5,-51.5</position>
<input>
<ID>N_in0</ID>1657 </input>
<input>
<ID>N_in1</ID>4136 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5356</ID>
<type>BA_TRI_STATE</type>
<position>327.5,-858</position>
<input>
<ID>ENABLE_0</ID>3807 </input>
<input>
<ID>IN_0</ID>3808 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2278</ID>
<type>HA_JUNC_2</type>
<position>374.5,-52</position>
<input>
<ID>N_in0</ID>1658 </input>
<input>
<ID>N_in1</ID>4138 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5357</ID>
<type>AE_DFF_LOW</type>
<position>308.5,-850.5</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3808 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2279</ID>
<type>HA_JUNC_2</type>
<position>404.5,-51.5</position>
<input>
<ID>N_in0</ID>1659 </input>
<input>
<ID>N_in1</ID>4140 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5358</ID>
<type>AA_AND2</type>
<position>352,-858</position>
<input>
<ID>IN_0</ID>3810 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3809 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2280</ID>
<type>HA_JUNC_2</type>
<position>435.5,-51.5</position>
<input>
<ID>N_in0</ID>1660 </input>
<input>
<ID>N_in1</ID>4142 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5359</ID>
<type>BA_TRI_STATE</type>
<position>359,-858</position>
<input>
<ID>ENABLE_0</ID>3809 </input>
<input>
<ID>IN_0</ID>3810 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2281</ID>
<type>HA_JUNC_2</type>
<position>466.5,-52</position>
<input>
<ID>N_in0</ID>1661 </input>
<input>
<ID>N_in1</ID>4144 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5360</ID>
<type>AE_DFF_LOW</type>
<position>339.5,-850.5</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3810 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2282</ID>
<type>HA_JUNC_2</type>
<position>278.5,-44.5</position>
<input>
<ID>N_in0</ID>1662 </input>
<input>
<ID>N_in1</ID>4131 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5361</ID>
<type>AA_AND2</type>
<position>381.5,-858</position>
<input>
<ID>IN_0</ID>3812 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3811 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2283</ID>
<type>HA_JUNC_2</type>
<position>278.5,-201.5</position>
<input>
<ID>N_in0</ID>4159 </input>
<input>
<ID>N_in1</ID>1662 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5362</ID>
<type>BA_TRI_STATE</type>
<position>388.5,-858</position>
<input>
<ID>ENABLE_0</ID>3811 </input>
<input>
<ID>IN_0</ID>3812 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2284</ID>
<type>HA_JUNC_2</type>
<position>341.5,-200.5</position>
<input>
<ID>N_in0</ID>4155 </input>
<input>
<ID>N_in1</ID>1664 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5363</ID>
<type>AE_DFF_LOW</type>
<position>369.5,-850.5</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3812 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2285</ID>
<type>HA_JUNC_2</type>
<position>372,-200</position>
<input>
<ID>N_in0</ID>4153 </input>
<input>
<ID>N_in1</ID>1665 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5364</ID>
<type>AA_AND2</type>
<position>413,-858</position>
<input>
<ID>IN_0</ID>3814 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3813 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2286</ID>
<type>HA_JUNC_2</type>
<position>402.5,-200</position>
<input>
<ID>N_in0</ID>4152 </input>
<input>
<ID>N_in1</ID>1666 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5365</ID>
<type>BA_TRI_STATE</type>
<position>420,-858</position>
<input>
<ID>ENABLE_0</ID>3813 </input>
<input>
<ID>IN_0</ID>3814 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2287</ID>
<type>HA_JUNC_2</type>
<position>433.5,-200</position>
<input>
<ID>N_in0</ID>4150 </input>
<input>
<ID>N_in1</ID>1667 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5366</ID>
<type>AE_DFF_LOW</type>
<position>400.5,-850.5</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3814 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2288</ID>
<type>HA_JUNC_2</type>
<position>464.5,-200.5</position>
<input>
<ID>N_in0</ID>4148 </input>
<input>
<ID>N_in1</ID>1668 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5367</ID>
<type>AA_AND2</type>
<position>443.5,-858</position>
<input>
<ID>IN_0</ID>3816 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3815 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2289</ID>
<type>HA_JUNC_2</type>
<position>495,-200</position>
<input>
<ID>N_in0</ID>4146 </input>
<input>
<ID>N_in1</ID>1669 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5368</ID>
<type>BA_TRI_STATE</type>
<position>450.5,-858</position>
<input>
<ID>ENABLE_0</ID>3815 </input>
<input>
<ID>IN_0</ID>3816 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2290</ID>
<type>HA_JUNC_2</type>
<position>495,-43</position>
<input>
<ID>N_in0</ID>1669 </input>
<input>
<ID>N_in1</ID>4145 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5369</ID>
<type>AE_DFF_LOW</type>
<position>431.5,-850.5</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3816 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2291</ID>
<type>HA_JUNC_2</type>
<position>464.5,-43.5</position>
<input>
<ID>N_in0</ID>1668 </input>
<input>
<ID>N_in1</ID>4143 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5370</ID>
<type>AA_AND2</type>
<position>475,-858</position>
<input>
<ID>IN_0</ID>3818 </input>
<input>
<ID>IN_1</ID>3772 </input>
<output>
<ID>OUT</ID>3817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2292</ID>
<type>HA_JUNC_2</type>
<position>433.5,-44.5</position>
<input>
<ID>N_in0</ID>1667 </input>
<input>
<ID>N_in1</ID>4141 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5371</ID>
<type>BA_TRI_STATE</type>
<position>482,-858</position>
<input>
<ID>ENABLE_0</ID>3817 </input>
<input>
<ID>IN_0</ID>3818 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2293</ID>
<type>HA_JUNC_2</type>
<position>402.5,-44.5</position>
<input>
<ID>N_in0</ID>1666 </input>
<input>
<ID>N_in1</ID>4139 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5372</ID>
<type>AE_DFF_LOW</type>
<position>462.5,-850.5</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3818 </output>
<input>
<ID>clock</ID>3771 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2294</ID>
<type>HA_JUNC_2</type>
<position>372,-44.5</position>
<input>
<ID>N_in0</ID>1665 </input>
<input>
<ID>N_in1</ID>4137 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5373</ID>
<type>AA_AND2</type>
<position>259,-842.5</position>
<input>
<ID>IN_0</ID>3820 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2295</ID>
<type>HA_JUNC_2</type>
<position>341.5,-44.5</position>
<input>
<ID>N_in0</ID>1664 </input>
<input>
<ID>N_in1</ID>4135 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5374</ID>
<type>BA_TRI_STATE</type>
<position>266,-842.5</position>
<input>
<ID>ENABLE_0</ID>3819 </input>
<input>
<ID>IN_0</ID>3820 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2296</ID>
<type>HA_JUNC_2</type>
<position>309.5,-44.5</position>
<input>
<ID>N_in0</ID>1663 </input>
<input>
<ID>N_in1</ID>4133 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5375</ID>
<type>AE_DFF_LOW</type>
<position>247,-835</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3820 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2297</ID>
<type>BE_DECODER_3x8</type>
<position>199.5,-117</position>
<input>
<ID>ENABLE</ID>69 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>1677 </output>
<output>
<ID>OUT_1</ID>1676 </output>
<output>
<ID>OUT_2</ID>1675 </output>
<output>
<ID>OUT_3</ID>1674 </output>
<output>
<ID>OUT_4</ID>1673 </output>
<output>
<ID>OUT_5</ID>1672 </output>
<output>
<ID>OUT_6</ID>1671 </output>
<output>
<ID>OUT_7</ID>1670 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>5376</ID>
<type>AA_AND2</type>
<position>290.5,-842.5</position>
<input>
<ID>IN_0</ID>3822 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3821 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2298</ID>
<type>BA_TRI_STATE</type>
<position>241.5,-131.5</position>
<input>
<ID>ENABLE_0</ID>1674 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5377</ID>
<type>BA_TRI_STATE</type>
<position>297.5,-842.5</position>
<input>
<ID>ENABLE_0</ID>3821 </input>
<input>
<ID>IN_0</ID>3822 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2299</ID>
<type>AA_AND2</type>
<position>235.5,-127</position>
<input>
<ID>IN_0</ID>1674 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1585 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5378</ID>
<type>AE_DFF_LOW</type>
<position>278,-835</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3822 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2300</ID>
<type>BA_TRI_STATE</type>
<position>241.5,-147.5</position>
<input>
<ID>ENABLE_0</ID>1675 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1588 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5379</ID>
<type>AA_AND2</type>
<position>321,-842.5</position>
<input>
<ID>IN_0</ID>3824 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3823 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2301</ID>
<type>AA_AND2</type>
<position>235.5,-142.5</position>
<input>
<ID>IN_0</ID>1675 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1587 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5380</ID>
<type>BA_TRI_STATE</type>
<position>328,-842.5</position>
<input>
<ID>ENABLE_0</ID>3823 </input>
<input>
<ID>IN_0</ID>3824 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2302</ID>
<type>BA_TRI_STATE</type>
<position>241.5,-163.5</position>
<input>
<ID>ENABLE_0</ID>1676 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5381</ID>
<type>AE_DFF_LOW</type>
<position>309,-835</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3824 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2303</ID>
<type>AA_AND2</type>
<position>235.5,-158.5</position>
<input>
<ID>IN_0</ID>1676 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5382</ID>
<type>AA_AND2</type>
<position>352.5,-842.5</position>
<input>
<ID>IN_0</ID>3826 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3825 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2304</ID>
<type>BA_TRI_STATE</type>
<position>241.5,-180.5</position>
<input>
<ID>ENABLE_0</ID>1677 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5383</ID>
<type>BA_TRI_STATE</type>
<position>359.5,-842.5</position>
<input>
<ID>ENABLE_0</ID>3825 </input>
<input>
<ID>IN_0</ID>3826 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2305</ID>
<type>AA_AND2</type>
<position>235.5,-175.5</position>
<input>
<ID>IN_0</ID>1677 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1653 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5384</ID>
<type>AE_DFF_LOW</type>
<position>340,-835</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3826 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2306</ID>
<type>AA_AND2</type>
<position>266.5,-117</position>
<input>
<ID>IN_0</ID>1679 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1678 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5385</ID>
<type>AA_AND2</type>
<position>382,-842.5</position>
<input>
<ID>IN_0</ID>3828 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3827 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2307</ID>
<type>BA_TRI_STATE</type>
<position>273.5,-117</position>
<input>
<ID>ENABLE_0</ID>1678 </input>
<input>
<ID>IN_0</ID>1679 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5386</ID>
<type>BA_TRI_STATE</type>
<position>389,-842.5</position>
<input>
<ID>ENABLE_0</ID>3827 </input>
<input>
<ID>IN_0</ID>3828 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2308</ID>
<type>AE_DFF_LOW</type>
<position>254.5,-109.5</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1679 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5387</ID>
<type>AE_DFF_LOW</type>
<position>370,-835</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3828 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2309</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-66.5</position>
<input>
<ID>ENABLE_0</ID>1670 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1743 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5388</ID>
<type>AA_AND2</type>
<position>413.5,-842.5</position>
<input>
<ID>IN_0</ID>3830 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3829 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2310</ID>
<type>AA_AND2</type>
<position>236,-62</position>
<input>
<ID>IN_0</ID>1670 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1744 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5389</ID>
<type>BA_TRI_STATE</type>
<position>420.5,-842.5</position>
<input>
<ID>ENABLE_0</ID>3829 </input>
<input>
<ID>IN_0</ID>3830 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2311</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-82.5</position>
<input>
<ID>ENABLE_0</ID>1671 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1579 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5390</ID>
<type>AE_DFF_LOW</type>
<position>401,-835</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3830 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2312</ID>
<type>AA_AND2</type>
<position>298,-117</position>
<input>
<ID>IN_0</ID>1681 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1680 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5391</ID>
<type>AA_AND2</type>
<position>444,-842.5</position>
<input>
<ID>IN_0</ID>3832 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3831 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2313</ID>
<type>AA_AND2</type>
<position>235.5,-77.5</position>
<input>
<ID>IN_0</ID>1671 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5392</ID>
<type>BA_TRI_STATE</type>
<position>451,-842.5</position>
<input>
<ID>ENABLE_0</ID>3831 </input>
<input>
<ID>IN_0</ID>3832 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2314</ID>
<type>BA_TRI_STATE</type>
<position>305,-117</position>
<input>
<ID>ENABLE_0</ID>1680 </input>
<input>
<ID>IN_0</ID>1681 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5393</ID>
<type>AE_DFF_LOW</type>
<position>432,-835</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3832 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2315</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-98.5</position>
<input>
<ID>ENABLE_0</ID>1672 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1581 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5394</ID>
<type>AA_AND2</type>
<position>475.5,-842.5</position>
<input>
<ID>IN_0</ID>3834 </input>
<input>
<ID>IN_1</ID>3770 </input>
<output>
<ID>OUT</ID>3833 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2316</ID>
<type>AE_DFF_LOW</type>
<position>285.5,-109.5</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1681 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5395</ID>
<type>BA_TRI_STATE</type>
<position>482.5,-842.5</position>
<input>
<ID>ENABLE_0</ID>3833 </input>
<input>
<ID>IN_0</ID>3834 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2317</ID>
<type>AA_AND2</type>
<position>235.5,-93.5</position>
<input>
<ID>IN_0</ID>1672 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1582 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5396</ID>
<type>AE_DFF_LOW</type>
<position>463,-835</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3834 </output>
<input>
<ID>clock</ID>3769 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2318</ID>
<type>AA_AND2</type>
<position>328.5,-117</position>
<input>
<ID>IN_0</ID>1683 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1682 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5397</ID>
<type>HA_JUNC_2</type>
<position>335.5,-760.5</position>
<input>
<ID>N_in0</ID>3841 </input>
<input>
<ID>N_in1</ID>4204 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2319</ID>
<type>BA_TRI_STATE</type>
<position>242.5,-115.5</position>
<input>
<ID>ENABLE_0</ID>1673 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>1584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5398</ID>
<type>HA_JUNC_2</type>
<position>366.5,-761</position>
<input>
<ID>N_in0</ID>3842 </input>
<input>
<ID>N_in1</ID>4202 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2320</ID>
<type>BA_TRI_STATE</type>
<position>335.5,-117</position>
<input>
<ID>ENABLE_0</ID>1682 </input>
<input>
<ID>IN_0</ID>1683 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5399</ID>
<type>HA_JUNC_2</type>
<position>396.5,-760.5</position>
<input>
<ID>N_in0</ID>3843 </input>
<input>
<ID>N_in1</ID>4200 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2321</ID>
<type>AA_AND2</type>
<position>235.5,-110.5</position>
<input>
<ID>IN_0</ID>1673 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>1583 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5400</ID>
<type>HA_JUNC_2</type>
<position>427.5,-760.5</position>
<input>
<ID>N_in0</ID>3844 </input>
<input>
<ID>N_in1</ID>4198 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2322</ID>
<type>AE_DFF_LOW</type>
<position>316.5,-109.5</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1683 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5401</ID>
<type>HA_JUNC_2</type>
<position>458.5,-761</position>
<input>
<ID>N_in0</ID>3845 </input>
<input>
<ID>N_in1</ID>4196 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2323</ID>
<type>AA_AND2</type>
<position>360,-117</position>
<input>
<ID>IN_0</ID>1685 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1684 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5402</ID>
<type>HA_JUNC_2</type>
<position>270.5,-753.5</position>
<input>
<ID>N_in0</ID>3846 </input>
<input>
<ID>N_in1</ID>4207 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2324</ID>
<type>BA_TRI_STATE</type>
<position>367,-117</position>
<input>
<ID>ENABLE_0</ID>1684 </input>
<input>
<ID>IN_0</ID>1685 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2325</ID>
<type>AE_DFF_LOW</type>
<position>347.5,-109.5</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1685 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2326</ID>
<type>AA_AND2</type>
<position>389.5,-117</position>
<input>
<ID>IN_0</ID>1687 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1686 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2327</ID>
<type>BA_TRI_STATE</type>
<position>396.5,-117</position>
<input>
<ID>ENABLE_0</ID>1686 </input>
<input>
<ID>IN_0</ID>1687 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2328</ID>
<type>AE_DFF_LOW</type>
<position>377.5,-109.5</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1687 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2329</ID>
<type>AA_AND2</type>
<position>421,-117</position>
<input>
<ID>IN_0</ID>1689 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1688 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2330</ID>
<type>BA_TRI_STATE</type>
<position>428,-117</position>
<input>
<ID>ENABLE_0</ID>1688 </input>
<input>
<ID>IN_0</ID>1689 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2331</ID>
<type>AE_DFF_LOW</type>
<position>408.5,-109.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1689 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5410</ID>
<type>HA_JUNC_2</type>
<position>487,-752</position>
<input>
<ID>N_in0</ID>3853 </input>
<input>
<ID>N_in1</ID>4194 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2332</ID>
<type>AA_AND2</type>
<position>451.5,-117</position>
<input>
<ID>IN_0</ID>1691 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1690 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5411</ID>
<type>HA_JUNC_2</type>
<position>456.5,-752.5</position>
<input>
<ID>N_in0</ID>3852 </input>
<input>
<ID>N_in1</ID>4195 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2333</ID>
<type>BA_TRI_STATE</type>
<position>458.5,-117</position>
<input>
<ID>ENABLE_0</ID>1690 </input>
<input>
<ID>IN_0</ID>1691 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5412</ID>
<type>HA_JUNC_2</type>
<position>425.5,-753.5</position>
<input>
<ID>N_in0</ID>3851 </input>
<input>
<ID>N_in1</ID>4197 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2334</ID>
<type>AE_DFF_LOW</type>
<position>439.5,-109.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1691 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5413</ID>
<type>HA_JUNC_2</type>
<position>394.5,-753.5</position>
<input>
<ID>N_in0</ID>3850 </input>
<input>
<ID>N_in1</ID>4199 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2335</ID>
<type>AA_AND2</type>
<position>483,-117</position>
<input>
<ID>IN_0</ID>1693 </input>
<input>
<ID>IN_1</ID>1584 </input>
<output>
<ID>OUT</ID>1692 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5414</ID>
<type>HA_JUNC_2</type>
<position>364,-753.5</position>
<input>
<ID>N_in0</ID>3849 </input>
<input>
<ID>N_in1</ID>4201 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2336</ID>
<type>BA_TRI_STATE</type>
<position>490,-117</position>
<input>
<ID>ENABLE_0</ID>1692 </input>
<input>
<ID>IN_0</ID>1693 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5415</ID>
<type>HA_JUNC_2</type>
<position>333.5,-753.5</position>
<input>
<ID>N_in0</ID>3848 </input>
<input>
<ID>N_in1</ID>4203 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2337</ID>
<type>AE_DFF_LOW</type>
<position>470.5,-109.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1693 </output>
<input>
<ID>clock</ID>1583 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5416</ID>
<type>HA_JUNC_2</type>
<position>301.5,-753.5</position>
<input>
<ID>N_in0</ID>3847 </input>
<input>
<ID>N_in1</ID>4206 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>2338</ID>
<type>AA_AND2</type>
<position>267,-100</position>
<input>
<ID>IN_0</ID>1695 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1694 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5417</ID>
<type>BE_DECODER_3x8</type>
<position>191.5,-826</position>
<input>
<ID>ENABLE</ID>74 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>3861 </output>
<output>
<ID>OUT_1</ID>3860 </output>
<output>
<ID>OUT_2</ID>3859 </output>
<output>
<ID>OUT_3</ID>3858 </output>
<output>
<ID>OUT_4</ID>3857 </output>
<output>
<ID>OUT_5</ID>3856 </output>
<output>
<ID>OUT_6</ID>3855 </output>
<output>
<ID>OUT_7</ID>3854 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2339</ID>
<type>BA_TRI_STATE</type>
<position>274,-100</position>
<input>
<ID>ENABLE_0</ID>1694 </input>
<input>
<ID>IN_0</ID>1695 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5418</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-840.5</position>
<input>
<ID>ENABLE_0</ID>3858 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3770 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2340</ID>
<type>AE_DFF_LOW</type>
<position>255,-92.5</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1695 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5419</ID>
<type>AA_AND2</type>
<position>227.5,-836</position>
<input>
<ID>IN_0</ID>3858 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3769 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2341</ID>
<type>AA_AND2</type>
<position>298.5,-100</position>
<input>
<ID>IN_0</ID>1697 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1696 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5420</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-856.5</position>
<input>
<ID>ENABLE_0</ID>3859 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2342</ID>
<type>BA_TRI_STATE</type>
<position>305.5,-100</position>
<input>
<ID>ENABLE_0</ID>1696 </input>
<input>
<ID>IN_0</ID>1697 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5421</ID>
<type>AA_AND2</type>
<position>227.5,-851.5</position>
<input>
<ID>IN_0</ID>3859 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2343</ID>
<type>AE_DFF_LOW</type>
<position>286,-92.5</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1697 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5422</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-872.5</position>
<input>
<ID>ENABLE_0</ID>3860 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3836 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2344</ID>
<type>AA_AND2</type>
<position>329,-100</position>
<input>
<ID>IN_0</ID>1699 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5423</ID>
<type>AA_AND2</type>
<position>227.5,-867.5</position>
<input>
<ID>IN_0</ID>3860 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3835 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2345</ID>
<type>BA_TRI_STATE</type>
<position>336,-100</position>
<input>
<ID>ENABLE_0</ID>1698 </input>
<input>
<ID>IN_0</ID>1699 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5424</ID>
<type>BA_TRI_STATE</type>
<position>233.5,-889.5</position>
<input>
<ID>ENABLE_0</ID>3861 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3838 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2346</ID>
<type>AE_DFF_LOW</type>
<position>317,-92.5</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1699 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5425</ID>
<type>AA_AND2</type>
<position>227.5,-884.5</position>
<input>
<ID>IN_0</ID>3861 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3837 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2347</ID>
<type>AA_AND2</type>
<position>360.5,-100</position>
<input>
<ID>IN_0</ID>1701 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1700 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5426</ID>
<type>AA_AND2</type>
<position>258.5,-826</position>
<input>
<ID>IN_0</ID>3863 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3862 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2348</ID>
<type>BA_TRI_STATE</type>
<position>367.5,-100</position>
<input>
<ID>ENABLE_0</ID>1700 </input>
<input>
<ID>IN_0</ID>1701 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5427</ID>
<type>BA_TRI_STATE</type>
<position>265.5,-826</position>
<input>
<ID>ENABLE_0</ID>3862 </input>
<input>
<ID>IN_0</ID>3863 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2349</ID>
<type>AE_DFF_LOW</type>
<position>348,-92.5</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1701 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5428</ID>
<type>AE_DFF_LOW</type>
<position>246.5,-818.5</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3863 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2350</ID>
<type>AA_AND2</type>
<position>390,-100</position>
<input>
<ID>IN_0</ID>1703 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1702 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5429</ID>
<type>BA_TRI_STATE</type>
<position>234.5,-775.5</position>
<input>
<ID>ENABLE_0</ID>3854 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3927 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2351</ID>
<type>BA_TRI_STATE</type>
<position>397,-100</position>
<input>
<ID>ENABLE_0</ID>1702 </input>
<input>
<ID>IN_0</ID>1703 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5430</ID>
<type>AA_AND2</type>
<position>228,-771</position>
<input>
<ID>IN_0</ID>3854 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3928 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2352</ID>
<type>AE_DFF_LOW</type>
<position>378,-92.5</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1703 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5431</ID>
<type>BA_TRI_STATE</type>
<position>234.5,-791.5</position>
<input>
<ID>ENABLE_0</ID>3855 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3763 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2353</ID>
<type>AA_AND2</type>
<position>421.5,-100</position>
<input>
<ID>IN_0</ID>1705 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1704 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5432</ID>
<type>AA_AND2</type>
<position>290,-826</position>
<input>
<ID>IN_0</ID>3865 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3864 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2354</ID>
<type>BA_TRI_STATE</type>
<position>428.5,-100</position>
<input>
<ID>ENABLE_0</ID>1704 </input>
<input>
<ID>IN_0</ID>1705 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5433</ID>
<type>AA_AND2</type>
<position>227.5,-786.5</position>
<input>
<ID>IN_0</ID>3855 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3764 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2355</ID>
<type>AE_DFF_LOW</type>
<position>409,-92.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1705 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5434</ID>
<type>BA_TRI_STATE</type>
<position>297,-826</position>
<input>
<ID>ENABLE_0</ID>3864 </input>
<input>
<ID>IN_0</ID>3865 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2356</ID>
<type>AA_AND2</type>
<position>452,-100</position>
<input>
<ID>IN_0</ID>1707 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1706 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5435</ID>
<type>BA_TRI_STATE</type>
<position>234.5,-807.5</position>
<input>
<ID>ENABLE_0</ID>3856 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3765 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2357</ID>
<type>BA_TRI_STATE</type>
<position>459,-100</position>
<input>
<ID>ENABLE_0</ID>1706 </input>
<input>
<ID>IN_0</ID>1707 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5436</ID>
<type>AE_DFF_LOW</type>
<position>277.5,-818.5</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3865 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2358</ID>
<type>AE_DFF_LOW</type>
<position>440,-92.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1707 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5437</ID>
<type>AA_AND2</type>
<position>227.5,-802.5</position>
<input>
<ID>IN_0</ID>3856 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2359</ID>
<type>AA_AND2</type>
<position>483.5,-100</position>
<input>
<ID>IN_0</ID>1709 </input>
<input>
<ID>IN_1</ID>1581 </input>
<output>
<ID>OUT</ID>1708 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5438</ID>
<type>AA_AND2</type>
<position>320.5,-826</position>
<input>
<ID>IN_0</ID>3867 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3866 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2360</ID>
<type>BA_TRI_STATE</type>
<position>490.5,-100</position>
<input>
<ID>ENABLE_0</ID>1708 </input>
<input>
<ID>IN_0</ID>1709 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5439</ID>
<type>BA_TRI_STATE</type>
<position>234.5,-824.5</position>
<input>
<ID>ENABLE_0</ID>3857 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3768 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2361</ID>
<type>AE_DFF_LOW</type>
<position>471,-92.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1709 </output>
<input>
<ID>clock</ID>1582 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5440</ID>
<type>BA_TRI_STATE</type>
<position>327.5,-826</position>
<input>
<ID>ENABLE_0</ID>3866 </input>
<input>
<ID>IN_0</ID>3867 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5441</ID>
<type>AA_AND2</type>
<position>227.5,-819.5</position>
<input>
<ID>IN_0</ID>3857 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3767 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2362</ID>
<type>AA_AND2</type>
<position>267.5,-84</position>
<input>
<ID>IN_0</ID>1711 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1710 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5442</ID>
<type>AE_DFF_LOW</type>
<position>308.5,-818.5</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3867 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2363</ID>
<type>BA_TRI_STATE</type>
<position>274.5,-84</position>
<input>
<ID>ENABLE_0</ID>1710 </input>
<input>
<ID>IN_0</ID>1711 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5443</ID>
<type>AA_AND2</type>
<position>352,-826</position>
<input>
<ID>IN_0</ID>3869 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3868 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2364</ID>
<type>AE_DFF_LOW</type>
<position>255.5,-76.5</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1711 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5444</ID>
<type>BA_TRI_STATE</type>
<position>359,-826</position>
<input>
<ID>ENABLE_0</ID>3868 </input>
<input>
<ID>IN_0</ID>3869 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2365</ID>
<type>AA_AND2</type>
<position>299,-84</position>
<input>
<ID>IN_0</ID>1713 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1712 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5445</ID>
<type>AE_DFF_LOW</type>
<position>339.5,-818.5</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3869 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2366</ID>
<type>BA_TRI_STATE</type>
<position>306,-84</position>
<input>
<ID>ENABLE_0</ID>1712 </input>
<input>
<ID>IN_0</ID>1713 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5446</ID>
<type>AA_AND2</type>
<position>381.5,-826</position>
<input>
<ID>IN_0</ID>3871 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3870 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2367</ID>
<type>AE_DFF_LOW</type>
<position>286.5,-76.5</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1713 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5447</ID>
<type>BA_TRI_STATE</type>
<position>388.5,-826</position>
<input>
<ID>ENABLE_0</ID>3870 </input>
<input>
<ID>IN_0</ID>3871 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2368</ID>
<type>AA_AND2</type>
<position>329.5,-84</position>
<input>
<ID>IN_0</ID>1715 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1714 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5448</ID>
<type>AE_DFF_LOW</type>
<position>369.5,-818.5</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3871 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2369</ID>
<type>BA_TRI_STATE</type>
<position>336.5,-84</position>
<input>
<ID>ENABLE_0</ID>1714 </input>
<input>
<ID>IN_0</ID>1715 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5449</ID>
<type>AA_AND2</type>
<position>413,-826</position>
<input>
<ID>IN_0</ID>3873 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3872 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2370</ID>
<type>AE_DFF_LOW</type>
<position>317.5,-76.5</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1715 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5450</ID>
<type>BA_TRI_STATE</type>
<position>420,-826</position>
<input>
<ID>ENABLE_0</ID>3872 </input>
<input>
<ID>IN_0</ID>3873 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2371</ID>
<type>AA_AND2</type>
<position>361,-84</position>
<input>
<ID>IN_0</ID>1717 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1716 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5451</ID>
<type>AE_DFF_LOW</type>
<position>400.5,-818.5</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3873 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2372</ID>
<type>BA_TRI_STATE</type>
<position>368,-84</position>
<input>
<ID>ENABLE_0</ID>1716 </input>
<input>
<ID>IN_0</ID>1717 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5452</ID>
<type>AA_AND2</type>
<position>443.5,-826</position>
<input>
<ID>IN_0</ID>3875 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3874 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2373</ID>
<type>AE_DFF_LOW</type>
<position>348.5,-76.5</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1717 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5453</ID>
<type>BA_TRI_STATE</type>
<position>450.5,-826</position>
<input>
<ID>ENABLE_0</ID>3874 </input>
<input>
<ID>IN_0</ID>3875 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2374</ID>
<type>AA_AND2</type>
<position>390.5,-84</position>
<input>
<ID>IN_0</ID>1719 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1718 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5454</ID>
<type>AE_DFF_LOW</type>
<position>431.5,-818.5</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3875 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2375</ID>
<type>BA_TRI_STATE</type>
<position>397.5,-84</position>
<input>
<ID>ENABLE_0</ID>1718 </input>
<input>
<ID>IN_0</ID>1719 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5455</ID>
<type>AA_AND2</type>
<position>475,-826</position>
<input>
<ID>IN_0</ID>3877 </input>
<input>
<ID>IN_1</ID>3768 </input>
<output>
<ID>OUT</ID>3876 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2376</ID>
<type>AE_DFF_LOW</type>
<position>378.5,-76.5</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1719 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5456</ID>
<type>BA_TRI_STATE</type>
<position>482,-826</position>
<input>
<ID>ENABLE_0</ID>3876 </input>
<input>
<ID>IN_0</ID>3877 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2377</ID>
<type>AA_AND2</type>
<position>422,-84</position>
<input>
<ID>IN_0</ID>1721 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1720 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5457</ID>
<type>AE_DFF_LOW</type>
<position>462.5,-818.5</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3877 </output>
<input>
<ID>clock</ID>3767 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2378</ID>
<type>BA_TRI_STATE</type>
<position>429,-84</position>
<input>
<ID>ENABLE_0</ID>1720 </input>
<input>
<ID>IN_0</ID>1721 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5458</ID>
<type>AA_AND2</type>
<position>259,-809</position>
<input>
<ID>IN_0</ID>3879 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3878 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2379</ID>
<type>AE_DFF_LOW</type>
<position>409.5,-76.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1721 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5459</ID>
<type>BA_TRI_STATE</type>
<position>266,-809</position>
<input>
<ID>ENABLE_0</ID>3878 </input>
<input>
<ID>IN_0</ID>3879 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2380</ID>
<type>AA_AND2</type>
<position>452.5,-84</position>
<input>
<ID>IN_0</ID>1723 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1722 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5460</ID>
<type>AE_DFF_LOW</type>
<position>247,-801.5</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3879 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2381</ID>
<type>BA_TRI_STATE</type>
<position>459.5,-84</position>
<input>
<ID>ENABLE_0</ID>1722 </input>
<input>
<ID>IN_0</ID>1723 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5461</ID>
<type>AA_AND2</type>
<position>290.5,-809</position>
<input>
<ID>IN_0</ID>3881 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3880 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2382</ID>
<type>AE_DFF_LOW</type>
<position>440.5,-76.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1723 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5462</ID>
<type>BA_TRI_STATE</type>
<position>297.5,-809</position>
<input>
<ID>ENABLE_0</ID>3880 </input>
<input>
<ID>IN_0</ID>3881 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2383</ID>
<type>AA_AND2</type>
<position>484,-84</position>
<input>
<ID>IN_0</ID>1725 </input>
<input>
<ID>IN_1</ID>1579 </input>
<output>
<ID>OUT</ID>1724 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5463</ID>
<type>AE_DFF_LOW</type>
<position>278,-801.5</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3881 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2384</ID>
<type>BA_TRI_STATE</type>
<position>491,-84</position>
<input>
<ID>ENABLE_0</ID>1724 </input>
<input>
<ID>IN_0</ID>1725 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5464</ID>
<type>AA_AND2</type>
<position>321,-809</position>
<input>
<ID>IN_0</ID>3883 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3882 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2385</ID>
<type>AE_DFF_LOW</type>
<position>471.5,-76.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1725 </output>
<input>
<ID>clock</ID>1580 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5465</ID>
<type>BA_TRI_STATE</type>
<position>328,-809</position>
<input>
<ID>ENABLE_0</ID>3882 </input>
<input>
<ID>IN_0</ID>3883 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2386</ID>
<type>AA_AND2</type>
<position>268,-68.5</position>
<input>
<ID>IN_0</ID>1727 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1726 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5466</ID>
<type>AE_DFF_LOW</type>
<position>309,-801.5</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3883 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2387</ID>
<type>BA_TRI_STATE</type>
<position>275,-68.5</position>
<input>
<ID>ENABLE_0</ID>1726 </input>
<input>
<ID>IN_0</ID>1727 </input>
<output>
<ID>OUT_0</ID>1662 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5467</ID>
<type>AA_AND2</type>
<position>352.5,-809</position>
<input>
<ID>IN_0</ID>3885 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2388</ID>
<type>AE_DFF_LOW</type>
<position>256,-61</position>
<input>
<ID>IN_0</ID>1742 </input>
<output>
<ID>OUT_0</ID>1727 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5468</ID>
<type>BA_TRI_STATE</type>
<position>359.5,-809</position>
<input>
<ID>ENABLE_0</ID>3884 </input>
<input>
<ID>IN_0</ID>3885 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2389</ID>
<type>AA_AND2</type>
<position>299.5,-68.5</position>
<input>
<ID>IN_0</ID>1729 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1728 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5469</ID>
<type>AE_DFF_LOW</type>
<position>340,-801.5</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3885 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2390</ID>
<type>BA_TRI_STATE</type>
<position>306.5,-68.5</position>
<input>
<ID>ENABLE_0</ID>1728 </input>
<input>
<ID>IN_0</ID>1729 </input>
<output>
<ID>OUT_0</ID>1663 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5470</ID>
<type>AA_AND2</type>
<position>382,-809</position>
<input>
<ID>IN_0</ID>3887 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3886 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2391</ID>
<type>AE_DFF_LOW</type>
<position>287,-61</position>
<input>
<ID>IN_0</ID>1655 </input>
<output>
<ID>OUT_0</ID>1729 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5471</ID>
<type>BA_TRI_STATE</type>
<position>389,-809</position>
<input>
<ID>ENABLE_0</ID>3886 </input>
<input>
<ID>IN_0</ID>3887 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2392</ID>
<type>AA_AND2</type>
<position>330,-68.5</position>
<input>
<ID>IN_0</ID>1731 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1730 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5472</ID>
<type>AE_DFF_LOW</type>
<position>370,-801.5</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3887 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2393</ID>
<type>BA_TRI_STATE</type>
<position>337,-68.5</position>
<input>
<ID>ENABLE_0</ID>1730 </input>
<input>
<ID>IN_0</ID>1731 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5473</ID>
<type>AA_AND2</type>
<position>413.5,-809</position>
<input>
<ID>IN_0</ID>3889 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3888 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2394</ID>
<type>AE_DFF_LOW</type>
<position>318,-61</position>
<input>
<ID>IN_0</ID>1656 </input>
<output>
<ID>OUT_0</ID>1731 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5474</ID>
<type>BA_TRI_STATE</type>
<position>420.5,-809</position>
<input>
<ID>ENABLE_0</ID>3888 </input>
<input>
<ID>IN_0</ID>3889 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2395</ID>
<type>AA_AND2</type>
<position>361.5,-68.5</position>
<input>
<ID>IN_0</ID>1733 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1732 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5475</ID>
<type>AE_DFF_LOW</type>
<position>401,-801.5</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3889 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2396</ID>
<type>BA_TRI_STATE</type>
<position>368.5,-68.5</position>
<input>
<ID>ENABLE_0</ID>1732 </input>
<input>
<ID>IN_0</ID>1733 </input>
<output>
<ID>OUT_0</ID>1665 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5476</ID>
<type>AA_AND2</type>
<position>444,-809</position>
<input>
<ID>IN_0</ID>3891 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3890 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2397</ID>
<type>AE_DFF_LOW</type>
<position>349,-61</position>
<input>
<ID>IN_0</ID>1657 </input>
<output>
<ID>OUT_0</ID>1733 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5477</ID>
<type>BA_TRI_STATE</type>
<position>451,-809</position>
<input>
<ID>ENABLE_0</ID>3890 </input>
<input>
<ID>IN_0</ID>3891 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2398</ID>
<type>AA_AND2</type>
<position>391,-68.5</position>
<input>
<ID>IN_0</ID>1735 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1734 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5478</ID>
<type>AE_DFF_LOW</type>
<position>432,-801.5</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3891 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2399</ID>
<type>BA_TRI_STATE</type>
<position>398,-68.5</position>
<input>
<ID>ENABLE_0</ID>1734 </input>
<input>
<ID>IN_0</ID>1735 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5479</ID>
<type>AA_AND2</type>
<position>475.5,-809</position>
<input>
<ID>IN_0</ID>3893 </input>
<input>
<ID>IN_1</ID>3765 </input>
<output>
<ID>OUT</ID>3892 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2400</ID>
<type>AE_DFF_LOW</type>
<position>379,-61</position>
<input>
<ID>IN_0</ID>1658 </input>
<output>
<ID>OUT_0</ID>1735 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5480</ID>
<type>BA_TRI_STATE</type>
<position>482.5,-809</position>
<input>
<ID>ENABLE_0</ID>3892 </input>
<input>
<ID>IN_0</ID>3893 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2401</ID>
<type>AA_AND2</type>
<position>422.5,-68.5</position>
<input>
<ID>IN_0</ID>1737 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1736 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5481</ID>
<type>AE_DFF_LOW</type>
<position>463,-801.5</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3893 </output>
<input>
<ID>clock</ID>3766 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2402</ID>
<type>BA_TRI_STATE</type>
<position>429.5,-68.5</position>
<input>
<ID>ENABLE_0</ID>1736 </input>
<input>
<ID>IN_0</ID>1737 </input>
<output>
<ID>OUT_0</ID>1667 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5482</ID>
<type>AA_AND2</type>
<position>259.5,-793</position>
<input>
<ID>IN_0</ID>3895 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3894 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2403</ID>
<type>AE_DFF_LOW</type>
<position>410,-61</position>
<input>
<ID>IN_0</ID>1659 </input>
<output>
<ID>OUT_0</ID>1737 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5483</ID>
<type>BA_TRI_STATE</type>
<position>266.5,-793</position>
<input>
<ID>ENABLE_0</ID>3894 </input>
<input>
<ID>IN_0</ID>3895 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2404</ID>
<type>AA_AND2</type>
<position>453,-68.5</position>
<input>
<ID>IN_0</ID>1739 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5484</ID>
<type>AE_DFF_LOW</type>
<position>247.5,-785.5</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3895 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2405</ID>
<type>BA_TRI_STATE</type>
<position>460,-68.5</position>
<input>
<ID>ENABLE_0</ID>1738 </input>
<input>
<ID>IN_0</ID>1739 </input>
<output>
<ID>OUT_0</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5485</ID>
<type>AA_AND2</type>
<position>291,-793</position>
<input>
<ID>IN_0</ID>3897 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3896 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2406</ID>
<type>AE_DFF_LOW</type>
<position>441,-61</position>
<input>
<ID>IN_0</ID>1660 </input>
<output>
<ID>OUT_0</ID>1739 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5486</ID>
<type>BA_TRI_STATE</type>
<position>298,-793</position>
<input>
<ID>ENABLE_0</ID>3896 </input>
<input>
<ID>IN_0</ID>3897 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2407</ID>
<type>AA_AND2</type>
<position>484.5,-68.5</position>
<input>
<ID>IN_0</ID>1741 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1740 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5487</ID>
<type>AE_DFF_LOW</type>
<position>278.5,-785.5</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3897 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2408</ID>
<type>BA_TRI_STATE</type>
<position>491.5,-68.5</position>
<input>
<ID>ENABLE_0</ID>1740 </input>
<input>
<ID>IN_0</ID>1741 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5488</ID>
<type>AA_AND2</type>
<position>321.5,-793</position>
<input>
<ID>IN_0</ID>3899 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3898 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2409</ID>
<type>AE_DFF_LOW</type>
<position>472,-61</position>
<input>
<ID>IN_0</ID>1661 </input>
<output>
<ID>OUT_0</ID>1741 </output>
<input>
<ID>clock</ID>1744 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5489</ID>
<type>BA_TRI_STATE</type>
<position>328.5,-793</position>
<input>
<ID>ENABLE_0</ID>3898 </input>
<input>
<ID>IN_0</ID>3899 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5490</ID>
<type>AE_DFF_LOW</type>
<position>309.5,-785.5</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3899 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5491</ID>
<type>AA_AND2</type>
<position>353,-793</position>
<input>
<ID>IN_0</ID>3901 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3900 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5492</ID>
<type>BA_TRI_STATE</type>
<position>360,-793</position>
<input>
<ID>ENABLE_0</ID>3900 </input>
<input>
<ID>IN_0</ID>3901 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5493</ID>
<type>AE_DFF_LOW</type>
<position>340.5,-785.5</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3901 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5494</ID>
<type>AA_AND2</type>
<position>382.5,-793</position>
<input>
<ID>IN_0</ID>3903 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3902 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5495</ID>
<type>BA_TRI_STATE</type>
<position>389.5,-793</position>
<input>
<ID>ENABLE_0</ID>3902 </input>
<input>
<ID>IN_0</ID>3903 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5496</ID>
<type>AE_DFF_LOW</type>
<position>370.5,-785.5</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3903 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5497</ID>
<type>AA_AND2</type>
<position>414,-793</position>
<input>
<ID>IN_0</ID>3905 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3904 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5498</ID>
<type>BA_TRI_STATE</type>
<position>421,-793</position>
<input>
<ID>ENABLE_0</ID>3904 </input>
<input>
<ID>IN_0</ID>3905 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5499</ID>
<type>AE_DFF_LOW</type>
<position>401.5,-785.5</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3905 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5500</ID>
<type>AA_AND2</type>
<position>444.5,-793</position>
<input>
<ID>IN_0</ID>3907 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3906 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5501</ID>
<type>BA_TRI_STATE</type>
<position>451.5,-793</position>
<input>
<ID>ENABLE_0</ID>3906 </input>
<input>
<ID>IN_0</ID>3907 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5502</ID>
<type>AE_DFF_LOW</type>
<position>432.5,-785.5</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3907 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5503</ID>
<type>AA_AND2</type>
<position>476,-793</position>
<input>
<ID>IN_0</ID>3909 </input>
<input>
<ID>IN_1</ID>3763 </input>
<output>
<ID>OUT</ID>3908 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5504</ID>
<type>BA_TRI_STATE</type>
<position>483,-793</position>
<input>
<ID>ENABLE_0</ID>3908 </input>
<input>
<ID>IN_0</ID>3909 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5505</ID>
<type>AE_DFF_LOW</type>
<position>463.5,-785.5</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3909 </output>
<input>
<ID>clock</ID>3764 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5506</ID>
<type>AA_AND2</type>
<position>260,-777.5</position>
<input>
<ID>IN_0</ID>3911 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3910 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5507</ID>
<type>BA_TRI_STATE</type>
<position>267,-777.5</position>
<input>
<ID>ENABLE_0</ID>3910 </input>
<input>
<ID>IN_0</ID>3911 </input>
<output>
<ID>OUT_0</ID>3846 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5508</ID>
<type>AE_DFF_LOW</type>
<position>248,-770</position>
<input>
<ID>IN_0</ID>3926 </input>
<output>
<ID>OUT_0</ID>3911 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5509</ID>
<type>AA_AND2</type>
<position>291.5,-777.5</position>
<input>
<ID>IN_0</ID>3913 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3912 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5510</ID>
<type>BA_TRI_STATE</type>
<position>298.5,-777.5</position>
<input>
<ID>ENABLE_0</ID>3912 </input>
<input>
<ID>IN_0</ID>3913 </input>
<output>
<ID>OUT_0</ID>3847 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5511</ID>
<type>AE_DFF_LOW</type>
<position>279,-770</position>
<input>
<ID>IN_0</ID>3839 </input>
<output>
<ID>OUT_0</ID>3913 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5512</ID>
<type>AA_AND2</type>
<position>322,-777.5</position>
<input>
<ID>IN_0</ID>3915 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3914 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5513</ID>
<type>BA_TRI_STATE</type>
<position>329,-777.5</position>
<input>
<ID>ENABLE_0</ID>3914 </input>
<input>
<ID>IN_0</ID>3915 </input>
<output>
<ID>OUT_0</ID>3848 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5514</ID>
<type>AE_DFF_LOW</type>
<position>310,-770</position>
<input>
<ID>IN_0</ID>3840 </input>
<output>
<ID>OUT_0</ID>3915 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5515</ID>
<type>AA_AND2</type>
<position>353.5,-777.5</position>
<input>
<ID>IN_0</ID>3917 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3916 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5516</ID>
<type>BA_TRI_STATE</type>
<position>360.5,-777.5</position>
<input>
<ID>ENABLE_0</ID>3916 </input>
<input>
<ID>IN_0</ID>3917 </input>
<output>
<ID>OUT_0</ID>3849 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5517</ID>
<type>AE_DFF_LOW</type>
<position>341,-770</position>
<input>
<ID>IN_0</ID>3841 </input>
<output>
<ID>OUT_0</ID>3917 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5518</ID>
<type>AA_AND2</type>
<position>383,-777.5</position>
<input>
<ID>IN_0</ID>3919 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3918 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5519</ID>
<type>BA_TRI_STATE</type>
<position>390,-777.5</position>
<input>
<ID>ENABLE_0</ID>3918 </input>
<input>
<ID>IN_0</ID>3919 </input>
<output>
<ID>OUT_0</ID>3850 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5520</ID>
<type>AE_DFF_LOW</type>
<position>371,-770</position>
<input>
<ID>IN_0</ID>3842 </input>
<output>
<ID>OUT_0</ID>3919 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5521</ID>
<type>AA_AND2</type>
<position>414.5,-777.5</position>
<input>
<ID>IN_0</ID>3921 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3920 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5522</ID>
<type>BA_TRI_STATE</type>
<position>421.5,-777.5</position>
<input>
<ID>ENABLE_0</ID>3920 </input>
<input>
<ID>IN_0</ID>3921 </input>
<output>
<ID>OUT_0</ID>3851 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5523</ID>
<type>AE_DFF_LOW</type>
<position>402,-770</position>
<input>
<ID>IN_0</ID>3843 </input>
<output>
<ID>OUT_0</ID>3921 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5524</ID>
<type>AA_AND2</type>
<position>445,-777.5</position>
<input>
<ID>IN_0</ID>3923 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3922 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5525</ID>
<type>BA_TRI_STATE</type>
<position>452,-777.5</position>
<input>
<ID>ENABLE_0</ID>3922 </input>
<input>
<ID>IN_0</ID>3923 </input>
<output>
<ID>OUT_0</ID>3852 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5526</ID>
<type>AE_DFF_LOW</type>
<position>433,-770</position>
<input>
<ID>IN_0</ID>3844 </input>
<output>
<ID>OUT_0</ID>3923 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5527</ID>
<type>AA_AND2</type>
<position>476.5,-777.5</position>
<input>
<ID>IN_0</ID>3925 </input>
<input>
<ID>IN_1</ID>3927 </input>
<output>
<ID>OUT</ID>3924 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5528</ID>
<type>BA_TRI_STATE</type>
<position>483.5,-777.5</position>
<input>
<ID>ENABLE_0</ID>3924 </input>
<input>
<ID>IN_0</ID>3925 </input>
<output>
<ID>OUT_0</ID>3853 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5529</ID>
<type>AE_DFF_LOW</type>
<position>464,-770</position>
<input>
<ID>IN_0</ID>3845 </input>
<output>
<ID>OUT_0</ID>3925 </output>
<input>
<ID>clock</ID>3928 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5530</ID>
<type>AA_AND2</type>
<position>263,386.5</position>
<input>
<ID>IN_0</ID>3930 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3929 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5531</ID>
<type>BA_TRI_STATE</type>
<position>270,386.5</position>
<input>
<ID>ENABLE_0</ID>3929 </input>
<input>
<ID>IN_0</ID>3930 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5532</ID>
<type>AE_DFF_LOW</type>
<position>251,394</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>3930 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5533</ID>
<type>HA_JUNC_2</type>
<position>247,375.5</position>
<input>
<ID>N_in0</ID>4097 </input>
<input>
<ID>N_in1</ID>4094 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5534</ID>
<type>HA_JUNC_2</type>
<position>278,375</position>
<input>
<ID>N_in0</ID>4099 </input>
<input>
<ID>N_in1</ID>4007 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5535</ID>
<type>HA_JUNC_2</type>
<position>310,375</position>
<input>
<ID>N_in0</ID>4102 </input>
<input>
<ID>N_in1</ID>4008 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5536</ID>
<type>HA_JUNC_2</type>
<position>341,376</position>
<input>
<ID>N_in0</ID>4104 </input>
<input>
<ID>N_in1</ID>4009 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5537</ID>
<type>HA_JUNC_2</type>
<position>371,377</position>
<input>
<ID>N_in0</ID>4106 </input>
<input>
<ID>N_in1</ID>4010 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5538</ID>
<type>HA_JUNC_2</type>
<position>402,377.5</position>
<input>
<ID>N_in0</ID>4108 </input>
<input>
<ID>N_in1</ID>4011 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5539</ID>
<type>HA_JUNC_2</type>
<position>464,376.5</position>
<input>
<ID>N_in0</ID>4112 </input>
<input>
<ID>N_in1</ID>4013 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5540</ID>
<type>HA_JUNC_2</type>
<position>433,378.5</position>
<input>
<ID>N_in0</ID>4110 </input>
<input>
<ID>N_in1</ID>4012 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5544</ID>
<type>AA_AND2</type>
<position>294.5,386.5</position>
<input>
<ID>IN_0</ID>3942 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3941 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5545</ID>
<type>BA_TRI_STATE</type>
<position>301.5,386.5</position>
<input>
<ID>ENABLE_0</ID>3941 </input>
<input>
<ID>IN_0</ID>3942 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5546</ID>
<type>AE_DFF_LOW</type>
<position>282,394</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>3942 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5547</ID>
<type>AA_AND2</type>
<position>325,386.5</position>
<input>
<ID>IN_0</ID>3944 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3943 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5548</ID>
<type>BA_TRI_STATE</type>
<position>332,386.5</position>
<input>
<ID>ENABLE_0</ID>3943 </input>
<input>
<ID>IN_0</ID>3944 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5549</ID>
<type>AE_DFF_LOW</type>
<position>313,394</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>3944 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5550</ID>
<type>AA_AND2</type>
<position>356.5,386.5</position>
<input>
<ID>IN_0</ID>3946 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5551</ID>
<type>BA_TRI_STATE</type>
<position>363.5,386.5</position>
<input>
<ID>ENABLE_0</ID>3945 </input>
<input>
<ID>IN_0</ID>3946 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5552</ID>
<type>AE_DFF_LOW</type>
<position>344,394</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>3946 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5553</ID>
<type>AA_AND2</type>
<position>386,386.5</position>
<input>
<ID>IN_0</ID>3948 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3947 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5554</ID>
<type>BA_TRI_STATE</type>
<position>393,386.5</position>
<input>
<ID>ENABLE_0</ID>3947 </input>
<input>
<ID>IN_0</ID>3948 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5555</ID>
<type>AE_DFF_LOW</type>
<position>374,394</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>3948 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5556</ID>
<type>AA_AND2</type>
<position>417.5,386.5</position>
<input>
<ID>IN_0</ID>3950 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3949 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5557</ID>
<type>BA_TRI_STATE</type>
<position>424.5,386.5</position>
<input>
<ID>ENABLE_0</ID>3949 </input>
<input>
<ID>IN_0</ID>3950 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5558</ID>
<type>AE_DFF_LOW</type>
<position>405,394</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>3950 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5559</ID>
<type>AA_AND2</type>
<position>448,386.5</position>
<input>
<ID>IN_0</ID>3952 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3951 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5560</ID>
<type>BA_TRI_STATE</type>
<position>455,386.5</position>
<input>
<ID>ENABLE_0</ID>3951 </input>
<input>
<ID>IN_0</ID>3952 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5561</ID>
<type>AE_DFF_LOW</type>
<position>436,394</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>3952 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5562</ID>
<type>AA_AND2</type>
<position>479.5,386.5</position>
<input>
<ID>IN_0</ID>3954 </input>
<input>
<ID>IN_1</ID>4006 </input>
<output>
<ID>OUT</ID>3953 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5563</ID>
<type>BA_TRI_STATE</type>
<position>486.5,386.5</position>
<input>
<ID>ENABLE_0</ID>3953 </input>
<input>
<ID>IN_0</ID>3954 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5564</ID>
<type>AE_DFF_LOW</type>
<position>467,394</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>3954 </output>
<input>
<ID>clock</ID>4005 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5565</ID>
<type>AA_AND2</type>
<position>263.5,403.5</position>
<input>
<ID>IN_0</ID>3956 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3955 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5566</ID>
<type>BA_TRI_STATE</type>
<position>270.5,403.5</position>
<input>
<ID>ENABLE_0</ID>3955 </input>
<input>
<ID>IN_0</ID>3956 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5567</ID>
<type>AE_DFF_LOW</type>
<position>251.5,411</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>3956 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5568</ID>
<type>AA_AND2</type>
<position>295,403.5</position>
<input>
<ID>IN_0</ID>3958 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3957 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5569</ID>
<type>BA_TRI_STATE</type>
<position>302,403.5</position>
<input>
<ID>ENABLE_0</ID>3957 </input>
<input>
<ID>IN_0</ID>3958 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5570</ID>
<type>AE_DFF_LOW</type>
<position>282.5,411</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>3958 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5571</ID>
<type>AA_AND2</type>
<position>325.5,403.5</position>
<input>
<ID>IN_0</ID>3960 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3959 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5572</ID>
<type>BA_TRI_STATE</type>
<position>332.5,403.5</position>
<input>
<ID>ENABLE_0</ID>3959 </input>
<input>
<ID>IN_0</ID>3960 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5573</ID>
<type>AE_DFF_LOW</type>
<position>313.5,411</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>3960 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5574</ID>
<type>AA_AND2</type>
<position>357,403.5</position>
<input>
<ID>IN_0</ID>3962 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3961 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5575</ID>
<type>BA_TRI_STATE</type>
<position>364,403.5</position>
<input>
<ID>ENABLE_0</ID>3961 </input>
<input>
<ID>IN_0</ID>3962 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5576</ID>
<type>AE_DFF_LOW</type>
<position>344.5,411</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>3962 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5577</ID>
<type>AA_AND2</type>
<position>386.5,403.5</position>
<input>
<ID>IN_0</ID>3964 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3963 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5578</ID>
<type>BA_TRI_STATE</type>
<position>393.5,403.5</position>
<input>
<ID>ENABLE_0</ID>3963 </input>
<input>
<ID>IN_0</ID>3964 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5579</ID>
<type>AE_DFF_LOW</type>
<position>374.5,411</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>3964 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5580</ID>
<type>AA_AND2</type>
<position>418,403.5</position>
<input>
<ID>IN_0</ID>3966 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3965 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5581</ID>
<type>BA_TRI_STATE</type>
<position>425,403.5</position>
<input>
<ID>ENABLE_0</ID>3965 </input>
<input>
<ID>IN_0</ID>3966 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5582</ID>
<type>AE_DFF_LOW</type>
<position>405.5,411</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>3966 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5583</ID>
<type>AA_AND2</type>
<position>448.5,403.5</position>
<input>
<ID>IN_0</ID>3968 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3967 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5584</ID>
<type>BA_TRI_STATE</type>
<position>455.5,403.5</position>
<input>
<ID>ENABLE_0</ID>3967 </input>
<input>
<ID>IN_0</ID>3968 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5585</ID>
<type>AE_DFF_LOW</type>
<position>436.5,411</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>3968 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5586</ID>
<type>AA_AND2</type>
<position>480,403.5</position>
<input>
<ID>IN_0</ID>3970 </input>
<input>
<ID>IN_1</ID>4004 </input>
<output>
<ID>OUT</ID>3969 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5587</ID>
<type>BA_TRI_STATE</type>
<position>487,403.5</position>
<input>
<ID>ENABLE_0</ID>3969 </input>
<input>
<ID>IN_0</ID>3970 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5588</ID>
<type>AE_DFF_LOW</type>
<position>467.5,411</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>3970 </output>
<input>
<ID>clock</ID>4003 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5589</ID>
<type>AA_AND2</type>
<position>264,419.5</position>
<input>
<ID>IN_0</ID>3972 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3971 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5590</ID>
<type>BA_TRI_STATE</type>
<position>271,419.5</position>
<input>
<ID>ENABLE_0</ID>3971 </input>
<input>
<ID>IN_0</ID>3972 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5591</ID>
<type>AE_DFF_LOW</type>
<position>252,427</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>3972 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5592</ID>
<type>AA_AND2</type>
<position>295.5,419.5</position>
<input>
<ID>IN_0</ID>3974 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3973 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5593</ID>
<type>BA_TRI_STATE</type>
<position>302.5,419.5</position>
<input>
<ID>ENABLE_0</ID>3973 </input>
<input>
<ID>IN_0</ID>3974 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5594</ID>
<type>AE_DFF_LOW</type>
<position>283,427</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>3974 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5595</ID>
<type>AA_AND2</type>
<position>326,419.5</position>
<input>
<ID>IN_0</ID>3976 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3975 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5596</ID>
<type>BA_TRI_STATE</type>
<position>333,419.5</position>
<input>
<ID>ENABLE_0</ID>3975 </input>
<input>
<ID>IN_0</ID>3976 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5597</ID>
<type>AE_DFF_LOW</type>
<position>314,427</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>3976 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5598</ID>
<type>AA_AND2</type>
<position>357.5,419.5</position>
<input>
<ID>IN_0</ID>3978 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3977 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5599</ID>
<type>BA_TRI_STATE</type>
<position>364.5,419.5</position>
<input>
<ID>ENABLE_0</ID>3977 </input>
<input>
<ID>IN_0</ID>3978 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5600</ID>
<type>AE_DFF_LOW</type>
<position>345,427</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>3978 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5601</ID>
<type>AA_AND2</type>
<position>387,419.5</position>
<input>
<ID>IN_0</ID>3980 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3979 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5602</ID>
<type>BA_TRI_STATE</type>
<position>394,419.5</position>
<input>
<ID>ENABLE_0</ID>3979 </input>
<input>
<ID>IN_0</ID>3980 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5603</ID>
<type>AE_DFF_LOW</type>
<position>375,427</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>3980 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5604</ID>
<type>AA_AND2</type>
<position>418.5,419.5</position>
<input>
<ID>IN_0</ID>3982 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3981 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5605</ID>
<type>BA_TRI_STATE</type>
<position>425.5,419.5</position>
<input>
<ID>ENABLE_0</ID>3981 </input>
<input>
<ID>IN_0</ID>3982 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5606</ID>
<type>AE_DFF_LOW</type>
<position>406,427</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>3982 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5607</ID>
<type>AA_AND2</type>
<position>449,419.5</position>
<input>
<ID>IN_0</ID>3984 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3983 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5608</ID>
<type>BA_TRI_STATE</type>
<position>456,419.5</position>
<input>
<ID>ENABLE_0</ID>3983 </input>
<input>
<ID>IN_0</ID>3984 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5609</ID>
<type>AE_DFF_LOW</type>
<position>437,427</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>3984 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5610</ID>
<type>AA_AND2</type>
<position>480.5,419.5</position>
<input>
<ID>IN_0</ID>3986 </input>
<input>
<ID>IN_1</ID>3940 </input>
<output>
<ID>OUT</ID>3985 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5611</ID>
<type>BA_TRI_STATE</type>
<position>487.5,419.5</position>
<input>
<ID>ENABLE_0</ID>3985 </input>
<input>
<ID>IN_0</ID>3986 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5612</ID>
<type>AE_DFF_LOW</type>
<position>468,427</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>3986 </output>
<input>
<ID>clock</ID>3939 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5613</ID>
<type>AA_AND2</type>
<position>264.5,435</position>
<input>
<ID>IN_0</ID>3988 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3987 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5614</ID>
<type>BA_TRI_STATE</type>
<position>271.5,435</position>
<input>
<ID>ENABLE_0</ID>3987 </input>
<input>
<ID>IN_0</ID>3988 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5615</ID>
<type>AE_DFF_LOW</type>
<position>252.5,442.5</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>3988 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5616</ID>
<type>AA_AND2</type>
<position>296,435</position>
<input>
<ID>IN_0</ID>3990 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3989 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5617</ID>
<type>BA_TRI_STATE</type>
<position>303,435</position>
<input>
<ID>ENABLE_0</ID>3989 </input>
<input>
<ID>IN_0</ID>3990 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5618</ID>
<type>AE_DFF_LOW</type>
<position>283.5,442.5</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>3990 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5619</ID>
<type>AA_AND2</type>
<position>326.5,435</position>
<input>
<ID>IN_0</ID>3992 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3991 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5620</ID>
<type>BA_TRI_STATE</type>
<position>333.5,435</position>
<input>
<ID>ENABLE_0</ID>3991 </input>
<input>
<ID>IN_0</ID>3992 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5621</ID>
<type>AE_DFF_LOW</type>
<position>314.5,442.5</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>3992 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5622</ID>
<type>AA_AND2</type>
<position>358,435</position>
<input>
<ID>IN_0</ID>3994 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3993 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5623</ID>
<type>BA_TRI_STATE</type>
<position>365,435</position>
<input>
<ID>ENABLE_0</ID>3993 </input>
<input>
<ID>IN_0</ID>3994 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5624</ID>
<type>AE_DFF_LOW</type>
<position>345.5,442.5</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>3994 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5625</ID>
<type>AA_AND2</type>
<position>387.5,435</position>
<input>
<ID>IN_0</ID>3996 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3995 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5626</ID>
<type>BA_TRI_STATE</type>
<position>394.5,435</position>
<input>
<ID>ENABLE_0</ID>3995 </input>
<input>
<ID>IN_0</ID>3996 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5627</ID>
<type>AE_DFF_LOW</type>
<position>375.5,442.5</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>3996 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5628</ID>
<type>AA_AND2</type>
<position>419,435</position>
<input>
<ID>IN_0</ID>3998 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3997 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5629</ID>
<type>BA_TRI_STATE</type>
<position>426,435</position>
<input>
<ID>ENABLE_0</ID>3997 </input>
<input>
<ID>IN_0</ID>3998 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5630</ID>
<type>AE_DFF_LOW</type>
<position>406.5,442.5</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>3998 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5631</ID>
<type>AA_AND2</type>
<position>449.5,435</position>
<input>
<ID>IN_0</ID>4000 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>3999 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5632</ID>
<type>BA_TRI_STATE</type>
<position>456.5,435</position>
<input>
<ID>ENABLE_0</ID>3999 </input>
<input>
<ID>IN_0</ID>4000 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5633</ID>
<type>AE_DFF_LOW</type>
<position>437.5,442.5</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>4000 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5634</ID>
<type>AA_AND2</type>
<position>481,435</position>
<input>
<ID>IN_0</ID>4002 </input>
<input>
<ID>IN_1</ID>3938 </input>
<output>
<ID>OUT</ID>4001 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5635</ID>
<type>BA_TRI_STATE</type>
<position>488,435</position>
<input>
<ID>ENABLE_0</ID>4001 </input>
<input>
<ID>IN_0</ID>4002 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5636</ID>
<type>AE_DFF_LOW</type>
<position>468.5,442.5</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>4002 </output>
<input>
<ID>clock</ID>3937 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5642</ID>
<type>HA_JUNC_2</type>
<position>276,524</position>
<input>
<ID>N_in0</ID>4014 </input>
<input>
<ID>N_in1</ID>9 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5643</ID>
<type>HA_JUNC_2</type>
<position>276,367</position>
<input>
<ID>N_in0</ID>4098 </input>
<input>
<ID>N_in1</ID>4014 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5644</ID>
<type>HA_JUNC_2</type>
<position>339,368</position>
<input>
<ID>N_in0</ID>4103 </input>
<input>
<ID>N_in1</ID>4016 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5645</ID>
<type>HA_JUNC_2</type>
<position>369.5,368.5</position>
<input>
<ID>N_in0</ID>4105 </input>
<input>
<ID>N_in1</ID>4017 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5646</ID>
<type>HA_JUNC_2</type>
<position>400,368.5</position>
<input>
<ID>N_in0</ID>4107 </input>
<input>
<ID>N_in1</ID>4018 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5647</ID>
<type>HA_JUNC_2</type>
<position>431,368.5</position>
<input>
<ID>N_in0</ID>4109 </input>
<input>
<ID>N_in1</ID>4019 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5648</ID>
<type>HA_JUNC_2</type>
<position>462,368</position>
<input>
<ID>N_in0</ID>4111 </input>
<input>
<ID>N_in1</ID>4020 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5649</ID>
<type>HA_JUNC_2</type>
<position>492.5,368.5</position>
<input>
<ID>N_in0</ID>4113 </input>
<input>
<ID>N_in1</ID>4021 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5650</ID>
<type>HA_JUNC_2</type>
<position>492.5,525.5</position>
<input>
<ID>N_in0</ID>4021 </input>
<input>
<ID>N_in1</ID>1 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5651</ID>
<type>HA_JUNC_2</type>
<position>462,525</position>
<input>
<ID>N_in0</ID>4020 </input>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5652</ID>
<type>HA_JUNC_2</type>
<position>431,524</position>
<input>
<ID>N_in0</ID>4019 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5653</ID>
<type>HA_JUNC_2</type>
<position>400,524</position>
<input>
<ID>N_in0</ID>4018 </input>
<input>
<ID>N_in1</ID>5 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5654</ID>
<type>HA_JUNC_2</type>
<position>369.5,524</position>
<input>
<ID>N_in0</ID>4017 </input>
<input>
<ID>N_in1</ID>6 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5655</ID>
<type>HA_JUNC_2</type>
<position>339,524</position>
<input>
<ID>N_in0</ID>4016 </input>
<input>
<ID>N_in1</ID>7 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5656</ID>
<type>HA_JUNC_2</type>
<position>307,524</position>
<input>
<ID>N_in0</ID>4015 </input>
<input>
<ID>N_in1</ID>8 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5657</ID>
<type>BE_DECODER_3x8</type>
<position>197,451.5</position>
<input>
<ID>ENABLE</ID>66 </input>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT_0</ID>4029 </output>
<output>
<ID>OUT_1</ID>4028 </output>
<output>
<ID>OUT_2</ID>4027 </output>
<output>
<ID>OUT_3</ID>4026 </output>
<output>
<ID>OUT_4</ID>4025 </output>
<output>
<ID>OUT_5</ID>4024 </output>
<output>
<ID>OUT_6</ID>4023 </output>
<output>
<ID>OUT_7</ID>4022 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>5658</ID>
<type>BA_TRI_STATE</type>
<position>239,437</position>
<input>
<ID>ENABLE_0</ID>4026 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3938 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5659</ID>
<type>AA_AND2</type>
<position>233,441.5</position>
<input>
<ID>IN_0</ID>4026 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3937 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5660</ID>
<type>BA_TRI_STATE</type>
<position>239,421</position>
<input>
<ID>ENABLE_0</ID>4027 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3940 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5661</ID>
<type>AA_AND2</type>
<position>233,426</position>
<input>
<ID>IN_0</ID>4027 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3939 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5662</ID>
<type>BA_TRI_STATE</type>
<position>239,405</position>
<input>
<ID>ENABLE_0</ID>4028 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>4004 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5663</ID>
<type>AA_AND2</type>
<position>233,410</position>
<input>
<ID>IN_0</ID>4028 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>4003 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5664</ID>
<type>BA_TRI_STATE</type>
<position>239,388</position>
<input>
<ID>ENABLE_0</ID>4029 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>4006 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5665</ID>
<type>AA_AND2</type>
<position>233,393</position>
<input>
<ID>IN_0</ID>4029 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>4005 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5666</ID>
<type>AA_AND2</type>
<position>264,451.5</position>
<input>
<ID>IN_0</ID>4031 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5667</ID>
<type>BA_TRI_STATE</type>
<position>271,451.5</position>
<input>
<ID>ENABLE_0</ID>4030 </input>
<input>
<ID>IN_0</ID>4031 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5668</ID>
<type>AE_DFF_LOW</type>
<position>252,459</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4031 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5669</ID>
<type>BA_TRI_STATE</type>
<position>240,502</position>
<input>
<ID>ENABLE_0</ID>4022 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>4095 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5670</ID>
<type>AA_AND2</type>
<position>233.5,506.5</position>
<input>
<ID>IN_0</ID>4022 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>4096 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5671</ID>
<type>BA_TRI_STATE</type>
<position>240,486</position>
<input>
<ID>ENABLE_0</ID>4023 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3931 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5672</ID>
<type>AA_AND2</type>
<position>295.5,451.5</position>
<input>
<ID>IN_0</ID>4033 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4032 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5673</ID>
<type>AA_AND2</type>
<position>233,491</position>
<input>
<ID>IN_0</ID>4023 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3932 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5674</ID>
<type>BA_TRI_STATE</type>
<position>302.5,451.5</position>
<input>
<ID>ENABLE_0</ID>4032 </input>
<input>
<ID>IN_0</ID>4033 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5675</ID>
<type>BA_TRI_STATE</type>
<position>240,470</position>
<input>
<ID>ENABLE_0</ID>4024 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3933 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5676</ID>
<type>AE_DFF_LOW</type>
<position>283,459</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>4033 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5677</ID>
<type>AA_AND2</type>
<position>233,475</position>
<input>
<ID>IN_0</ID>4024 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3934 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5678</ID>
<type>AA_AND2</type>
<position>326,451.5</position>
<input>
<ID>IN_0</ID>4035 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4034 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5679</ID>
<type>BA_TRI_STATE</type>
<position>240,453</position>
<input>
<ID>ENABLE_0</ID>4025 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3936 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5680</ID>
<type>BA_TRI_STATE</type>
<position>333,451.5</position>
<input>
<ID>ENABLE_0</ID>4034 </input>
<input>
<ID>IN_0</ID>4035 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5681</ID>
<type>AA_AND2</type>
<position>233,458</position>
<input>
<ID>IN_0</ID>4025 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>3935 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5682</ID>
<type>AE_DFF_LOW</type>
<position>314,459</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>4035 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5683</ID>
<type>AA_AND2</type>
<position>357.5,451.5</position>
<input>
<ID>IN_0</ID>4037 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4036 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5684</ID>
<type>BA_TRI_STATE</type>
<position>364.5,451.5</position>
<input>
<ID>ENABLE_0</ID>4036 </input>
<input>
<ID>IN_0</ID>4037 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5685</ID>
<type>AE_DFF_LOW</type>
<position>345,459</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>4037 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5686</ID>
<type>AA_AND2</type>
<position>387,451.5</position>
<input>
<ID>IN_0</ID>4039 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4038 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5687</ID>
<type>BA_TRI_STATE</type>
<position>394,451.5</position>
<input>
<ID>ENABLE_0</ID>4038 </input>
<input>
<ID>IN_0</ID>4039 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5688</ID>
<type>AE_DFF_LOW</type>
<position>375,459</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>4039 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5689</ID>
<type>AA_AND2</type>
<position>418.5,451.5</position>
<input>
<ID>IN_0</ID>4041 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4040 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5690</ID>
<type>BA_TRI_STATE</type>
<position>425.5,451.5</position>
<input>
<ID>ENABLE_0</ID>4040 </input>
<input>
<ID>IN_0</ID>4041 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5691</ID>
<type>AE_DFF_LOW</type>
<position>406,459</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>4041 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5692</ID>
<type>AA_AND2</type>
<position>449,451.5</position>
<input>
<ID>IN_0</ID>4043 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4042 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5693</ID>
<type>BA_TRI_STATE</type>
<position>456,451.5</position>
<input>
<ID>ENABLE_0</ID>4042 </input>
<input>
<ID>IN_0</ID>4043 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5694</ID>
<type>AE_DFF_LOW</type>
<position>437,459</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>4043 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5695</ID>
<type>AA_AND2</type>
<position>480.5,451.5</position>
<input>
<ID>IN_0</ID>4045 </input>
<input>
<ID>IN_1</ID>3936 </input>
<output>
<ID>OUT</ID>4044 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5696</ID>
<type>BA_TRI_STATE</type>
<position>487.5,451.5</position>
<input>
<ID>ENABLE_0</ID>4044 </input>
<input>
<ID>IN_0</ID>4045 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5697</ID>
<type>AE_DFF_LOW</type>
<position>468,459</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>4045 </output>
<input>
<ID>clock</ID>3935 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5698</ID>
<type>AA_AND2</type>
<position>264.5,468.5</position>
<input>
<ID>IN_0</ID>4047 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4046 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5699</ID>
<type>BA_TRI_STATE</type>
<position>271.5,468.5</position>
<input>
<ID>ENABLE_0</ID>4046 </input>
<input>
<ID>IN_0</ID>4047 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5700</ID>
<type>AE_DFF_LOW</type>
<position>252.5,476</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4047 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5701</ID>
<type>AA_AND2</type>
<position>296,468.5</position>
<input>
<ID>IN_0</ID>4049 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4048 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5702</ID>
<type>BA_TRI_STATE</type>
<position>303,468.5</position>
<input>
<ID>ENABLE_0</ID>4048 </input>
<input>
<ID>IN_0</ID>4049 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5703</ID>
<type>AE_DFF_LOW</type>
<position>283.5,476</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>4049 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5704</ID>
<type>AA_AND2</type>
<position>326.5,468.5</position>
<input>
<ID>IN_0</ID>4051 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4050 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5705</ID>
<type>BA_TRI_STATE</type>
<position>333.5,468.5</position>
<input>
<ID>ENABLE_0</ID>4050 </input>
<input>
<ID>IN_0</ID>4051 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5706</ID>
<type>AE_DFF_LOW</type>
<position>314.5,476</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>4051 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5707</ID>
<type>AA_AND2</type>
<position>358,468.5</position>
<input>
<ID>IN_0</ID>4053 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4052 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5708</ID>
<type>BA_TRI_STATE</type>
<position>365,468.5</position>
<input>
<ID>ENABLE_0</ID>4052 </input>
<input>
<ID>IN_0</ID>4053 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5709</ID>
<type>AE_DFF_LOW</type>
<position>345.5,476</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>4053 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5710</ID>
<type>AA_AND2</type>
<position>387.5,468.5</position>
<input>
<ID>IN_0</ID>4055 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4054 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5711</ID>
<type>BA_TRI_STATE</type>
<position>394.5,468.5</position>
<input>
<ID>ENABLE_0</ID>4054 </input>
<input>
<ID>IN_0</ID>4055 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5712</ID>
<type>AE_DFF_LOW</type>
<position>375.5,476</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>4055 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5713</ID>
<type>AA_AND2</type>
<position>419,468.5</position>
<input>
<ID>IN_0</ID>4057 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4056 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5714</ID>
<type>BA_TRI_STATE</type>
<position>426,468.5</position>
<input>
<ID>ENABLE_0</ID>4056 </input>
<input>
<ID>IN_0</ID>4057 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5715</ID>
<type>AE_DFF_LOW</type>
<position>406.5,476</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>4057 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5716</ID>
<type>AA_AND2</type>
<position>449.5,468.5</position>
<input>
<ID>IN_0</ID>4059 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4058 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5717</ID>
<type>BA_TRI_STATE</type>
<position>456.5,468.5</position>
<input>
<ID>ENABLE_0</ID>4058 </input>
<input>
<ID>IN_0</ID>4059 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5718</ID>
<type>AE_DFF_LOW</type>
<position>437.5,476</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>4059 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5719</ID>
<type>AA_AND2</type>
<position>481,468.5</position>
<input>
<ID>IN_0</ID>4061 </input>
<input>
<ID>IN_1</ID>3933 </input>
<output>
<ID>OUT</ID>4060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5720</ID>
<type>BA_TRI_STATE</type>
<position>488,468.5</position>
<input>
<ID>ENABLE_0</ID>4060 </input>
<input>
<ID>IN_0</ID>4061 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5721</ID>
<type>AE_DFF_LOW</type>
<position>468.5,476</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>4061 </output>
<input>
<ID>clock</ID>3934 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5722</ID>
<type>AA_AND2</type>
<position>265,484.5</position>
<input>
<ID>IN_0</ID>4063 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4062 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5723</ID>
<type>BA_TRI_STATE</type>
<position>272,484.5</position>
<input>
<ID>ENABLE_0</ID>4062 </input>
<input>
<ID>IN_0</ID>4063 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5724</ID>
<type>AE_DFF_LOW</type>
<position>253,492</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4063 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5725</ID>
<type>AA_AND2</type>
<position>296.5,484.5</position>
<input>
<ID>IN_0</ID>4065 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5726</ID>
<type>BA_TRI_STATE</type>
<position>303.5,484.5</position>
<input>
<ID>ENABLE_0</ID>4064 </input>
<input>
<ID>IN_0</ID>4065 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5727</ID>
<type>AE_DFF_LOW</type>
<position>284,492</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>4065 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5728</ID>
<type>AA_AND2</type>
<position>327,484.5</position>
<input>
<ID>IN_0</ID>4067 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4066 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5729</ID>
<type>BA_TRI_STATE</type>
<position>334,484.5</position>
<input>
<ID>ENABLE_0</ID>4066 </input>
<input>
<ID>IN_0</ID>4067 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5730</ID>
<type>AE_DFF_LOW</type>
<position>315,492</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>4067 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5731</ID>
<type>AA_AND2</type>
<position>358.5,484.5</position>
<input>
<ID>IN_0</ID>4069 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5732</ID>
<type>BA_TRI_STATE</type>
<position>365.5,484.5</position>
<input>
<ID>ENABLE_0</ID>4068 </input>
<input>
<ID>IN_0</ID>4069 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5733</ID>
<type>AE_DFF_LOW</type>
<position>346,492</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>4069 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5734</ID>
<type>AA_AND2</type>
<position>388,484.5</position>
<input>
<ID>IN_0</ID>4071 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5735</ID>
<type>BA_TRI_STATE</type>
<position>395,484.5</position>
<input>
<ID>ENABLE_0</ID>4070 </input>
<input>
<ID>IN_0</ID>4071 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5736</ID>
<type>AE_DFF_LOW</type>
<position>376,492</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>4071 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5737</ID>
<type>AA_AND2</type>
<position>419.5,484.5</position>
<input>
<ID>IN_0</ID>4073 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4072 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5738</ID>
<type>BA_TRI_STATE</type>
<position>426.5,484.5</position>
<input>
<ID>ENABLE_0</ID>4072 </input>
<input>
<ID>IN_0</ID>4073 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5739</ID>
<type>AE_DFF_LOW</type>
<position>407,492</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>4073 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5740</ID>
<type>AA_AND2</type>
<position>450,484.5</position>
<input>
<ID>IN_0</ID>4075 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5741</ID>
<type>BA_TRI_STATE</type>
<position>457,484.5</position>
<input>
<ID>ENABLE_0</ID>4074 </input>
<input>
<ID>IN_0</ID>4075 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5742</ID>
<type>AE_DFF_LOW</type>
<position>438,492</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>4075 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5743</ID>
<type>AA_AND2</type>
<position>481.5,484.5</position>
<input>
<ID>IN_0</ID>4077 </input>
<input>
<ID>IN_1</ID>3931 </input>
<output>
<ID>OUT</ID>4076 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5744</ID>
<type>BA_TRI_STATE</type>
<position>488.5,484.5</position>
<input>
<ID>ENABLE_0</ID>4076 </input>
<input>
<ID>IN_0</ID>4077 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5745</ID>
<type>AE_DFF_LOW</type>
<position>469,492</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>4077 </output>
<input>
<ID>clock</ID>3932 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5746</ID>
<type>AA_AND2</type>
<position>265.5,500</position>
<input>
<ID>IN_0</ID>4079 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4078 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5747</ID>
<type>BA_TRI_STATE</type>
<position>272.5,500</position>
<input>
<ID>ENABLE_0</ID>4078 </input>
<input>
<ID>IN_0</ID>4079 </input>
<output>
<ID>OUT_0</ID>4014 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5748</ID>
<type>AE_DFF_LOW</type>
<position>253.5,507.5</position>
<input>
<ID>IN_0</ID>4094 </input>
<output>
<ID>OUT_0</ID>4079 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5749</ID>
<type>AA_AND2</type>
<position>297,500</position>
<input>
<ID>IN_0</ID>4081 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5750</ID>
<type>BA_TRI_STATE</type>
<position>304,500</position>
<input>
<ID>ENABLE_0</ID>4080 </input>
<input>
<ID>IN_0</ID>4081 </input>
<output>
<ID>OUT_0</ID>4015 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5751</ID>
<type>AE_DFF_LOW</type>
<position>284.5,507.5</position>
<input>
<ID>IN_0</ID>4007 </input>
<output>
<ID>OUT_0</ID>4081 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5752</ID>
<type>AA_AND2</type>
<position>327.5,500</position>
<input>
<ID>IN_0</ID>4083 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4082 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5753</ID>
<type>BA_TRI_STATE</type>
<position>334.5,500</position>
<input>
<ID>ENABLE_0</ID>4082 </input>
<input>
<ID>IN_0</ID>4083 </input>
<output>
<ID>OUT_0</ID>4016 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5754</ID>
<type>AE_DFF_LOW</type>
<position>315.5,507.5</position>
<input>
<ID>IN_0</ID>4008 </input>
<output>
<ID>OUT_0</ID>4083 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5755</ID>
<type>AA_AND2</type>
<position>359,500</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4084 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5756</ID>
<type>BA_TRI_STATE</type>
<position>366,500</position>
<input>
<ID>ENABLE_0</ID>4084 </input>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>4017 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5757</ID>
<type>AE_DFF_LOW</type>
<position>346.5,507.5</position>
<input>
<ID>IN_0</ID>4009 </input>
<output>
<ID>OUT_0</ID>94 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5758</ID>
<type>AA_AND2</type>
<position>388.5,500</position>
<input>
<ID>IN_0</ID>4087 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4086 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5759</ID>
<type>BA_TRI_STATE</type>
<position>395.5,500</position>
<input>
<ID>ENABLE_0</ID>4086 </input>
<input>
<ID>IN_0</ID>4087 </input>
<output>
<ID>OUT_0</ID>4018 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5760</ID>
<type>AE_DFF_LOW</type>
<position>376.5,507.5</position>
<input>
<ID>IN_0</ID>4010 </input>
<output>
<ID>OUT_0</ID>4087 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5761</ID>
<type>AA_AND2</type>
<position>420,500</position>
<input>
<ID>IN_0</ID>4089 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4088 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5762</ID>
<type>BA_TRI_STATE</type>
<position>427,500</position>
<input>
<ID>ENABLE_0</ID>4088 </input>
<input>
<ID>IN_0</ID>4089 </input>
<output>
<ID>OUT_0</ID>4019 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5763</ID>
<type>AE_DFF_LOW</type>
<position>407.5,507.5</position>
<input>
<ID>IN_0</ID>4011 </input>
<output>
<ID>OUT_0</ID>4089 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5764</ID>
<type>AA_AND2</type>
<position>450.5,500</position>
<input>
<ID>IN_0</ID>4091 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4090 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5765</ID>
<type>BA_TRI_STATE</type>
<position>457.5,500</position>
<input>
<ID>ENABLE_0</ID>4090 </input>
<input>
<ID>IN_0</ID>4091 </input>
<output>
<ID>OUT_0</ID>4020 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5766</ID>
<type>AE_DFF_LOW</type>
<position>438.5,507.5</position>
<input>
<ID>IN_0</ID>4012 </input>
<output>
<ID>OUT_0</ID>4091 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5767</ID>
<type>AA_AND2</type>
<position>482,500</position>
<input>
<ID>IN_0</ID>4093 </input>
<input>
<ID>IN_1</ID>4095 </input>
<output>
<ID>OUT</ID>4092 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5768</ID>
<type>BA_TRI_STATE</type>
<position>489,500</position>
<input>
<ID>ENABLE_0</ID>4092 </input>
<input>
<ID>IN_0</ID>4093 </input>
<output>
<ID>OUT_0</ID>4021 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5769</ID>
<type>AE_DFF_LOW</type>
<position>469.5,507.5</position>
<input>
<ID>IN_0</ID>4013 </input>
<output>
<ID>OUT_0</ID>4093 </output>
<input>
<ID>clock</ID>4096 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5771</ID>
<type>HA_JUNC_2</type>
<position>305.5,367.5</position>
<input>
<ID>N_in0</ID>4101 </input>
<input>
<ID>N_in1</ID>4015 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5773</ID>
<type>HA_JUNC_2</type>
<position>303.5,191.5</position>
<input>
<ID>N_in0</ID>4129 </input>
<input>
<ID>N_in1</ID>3511 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5775</ID>
<type>HA_JUNC_2</type>
<position>309,4</position>
<input>
<ID>N_in0</ID>4133 </input>
<input>
<ID>N_in1</ID>3007 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5777</ID>
<type>HA_JUNC_2</type>
<position>306,-199.5</position>
<input>
<ID>N_in0</ID>4157 </input>
<input>
<ID>N_in1</ID>1663 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5779</ID>
<type>HA_JUNC_2</type>
<position>303.5,-374</position>
<input>
<ID>N_in0</ID>4165 </input>
<input>
<ID>N_in1</ID>2335 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5783</ID>
<type>HA_JUNC_2</type>
<position>306,-554</position>
<input>
<ID>N_in0</ID>4181 </input>
<input>
<ID>N_in1</ID>2503 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>5785</ID>
<type>HA_JUNC_2</type>
<position>301.5,-730</position>
<input>
<ID>N_in0</ID>4206 </input>
<input>
<ID>N_in1</ID>2839 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<wire>
<ID>3086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,12,250.5,151.5</points>
<connection>
<GID>4101</GID>
<name>N_in0</name></connection>
<connection>
<GID>4093</GID>
<name>N_in1</name></connection>
<intersection>31.5 14</intersection>
<intersection>48.5 12</intersection>
<intersection>64.5 10</intersection>
<intersection>80 8</intersection>
<intersection>96.5 6</intersection>
<intersection>113.5 4</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,145,254,145</points>
<connection>
<GID>4308</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,129.5,253.5,129.5</points>
<connection>
<GID>4284</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>250.5,113.5,253,113.5</points>
<connection>
<GID>4260</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>250.5,96.5,252.5,96.5</points>
<connection>
<GID>4228</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>250.5,80,253,80</points>
<connection>
<GID>4175</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>250.5,64.5,252.5,64.5</points>
<connection>
<GID>4151</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>250.5,48.5,252,48.5</points>
<connection>
<GID>4127</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>250.5,31.5,251.5,31.5</points>
<connection>
<GID>4092</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3087</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,134.5,482.5,134.5</points>
<connection>
<GID>4306</GID>
<name>IN_1</name></connection>
<connection>
<GID>4309</GID>
<name>IN_1</name></connection>
<connection>
<GID>4312</GID>
<name>IN_1</name></connection>
<connection>
<GID>4315</GID>
<name>IN_1</name></connection>
<connection>
<GID>4318</GID>
<name>IN_1</name></connection>
<connection>
<GID>4321</GID>
<name>IN_1</name></connection>
<connection>
<GID>4324</GID>
<name>IN_1</name></connection>
<connection>
<GID>4327</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,134.5,246,137.5</points>
<connection>
<GID>4229</GID>
<name>OUT_0</name></connection>
<intersection>134.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,526.5,492.5,534.5</points>
<connection>
<GID>5650</GID>
<name>N_in1</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3088</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,142,470,142</points>
<connection>
<GID>4230</GID>
<name>OUT</name></connection>
<connection>
<GID>4308</GID>
<name>clock</name></connection>
<connection>
<GID>4311</GID>
<name>clock</name></connection>
<connection>
<GID>4314</GID>
<name>clock</name></connection>
<connection>
<GID>4317</GID>
<name>clock</name></connection>
<connection>
<GID>4320</GID>
<name>clock</name></connection>
<connection>
<GID>4323</GID>
<name>clock</name></connection>
<connection>
<GID>4326</GID>
<name>clock</name></connection>
<connection>
<GID>4329</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>274,543,490.5,543</points>
<intersection>274 3</intersection>
<intersection>304 10</intersection>
<intersection>336 9</intersection>
<intersection>365.5 8</intersection>
<intersection>398 7</intersection>
<intersection>429 6</intersection>
<intersection>460 5</intersection>
<intersection>490.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>274,536,274,543</points>
<connection>
<GID>9</GID>
<name>ENABLE_0</name></connection>
<intersection>536 16</intersection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>490.5,537.5,490.5,543</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>460,536.5,460,543</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>429,536.5,429,543</points>
<connection>
<GID>4</GID>
<name>ENABLE_0</name></connection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>398,537,398,543</points>
<connection>
<GID>5</GID>
<name>ENABLE_0</name></connection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>365.5,536,365.5,543</points>
<intersection>536 14</intersection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>336,536.5,336,543</points>
<intersection>536.5 13</intersection>
<intersection>543 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>304,535.5,304,543</points>
<intersection>535.5 12</intersection>
<intersection>543 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>304,535.5,305,535.5</points>
<connection>
<GID>8</GID>
<name>ENABLE_0</name></connection>
<intersection>304 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>336,536.5,337,536.5</points>
<connection>
<GID>7</GID>
<name>ENABLE_0</name></connection>
<intersection>336 9</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>365.5,536,367.5,536</points>
<connection>
<GID>6</GID>
<name>ENABLE_0</name></connection>
<intersection>365.5 8</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>228.5,536,274,536</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>274 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462,526,462,533.5</points>
<connection>
<GID>5651</GID>
<name>N_in1</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431,525,431,533.5</points>
<connection>
<GID>5652</GID>
<name>N_in1</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,525,400,534</points>
<connection>
<GID>5653</GID>
<name>N_in1</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369.5,525,369.5,533</points>
<connection>
<GID>5654</GID>
<name>N_in1</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339,525,339,533.5</points>
<connection>
<GID>5655</GID>
<name>N_in1</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307,525,307,532.5</points>
<connection>
<GID>5656</GID>
<name>N_in1</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,525,276,533</points>
<connection>
<GID>5642</GID>
<name>N_in1</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,540,492.5,548.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462,539,462,549</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431,539,431,549</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,539.5,400,549</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369.5,538.5,369.5,549</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339,539,339,549</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307,538,307,549</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,538.5,276,548.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212.5,-889.5,212.5,523</points>
<intersection>-889.5 1</intersection>
<intersection>-872.5 2</intersection>
<intersection>-856.5 8</intersection>
<intersection>-840.5 6</intersection>
<intersection>-824.5 10</intersection>
<intersection>-807.5 12</intersection>
<intersection>-791.5 14</intersection>
<intersection>-775.5 16</intersection>
<intersection>-715.5 18</intersection>
<intersection>-698.5 20</intersection>
<intersection>-682.5 22</intersection>
<intersection>-666.5 24</intersection>
<intersection>-650.5 26</intersection>
<intersection>-633.5 28</intersection>
<intersection>-617.5 30</intersection>
<intersection>-601.5 32</intersection>
<intersection>-529.5 33</intersection>
<intersection>-512.5 35</intersection>
<intersection>-496.5 37</intersection>
<intersection>-480.5 39</intersection>
<intersection>-464.5 42</intersection>
<intersection>-447.5 44</intersection>
<intersection>-431.5 46</intersection>
<intersection>-415.5 48</intersection>
<intersection>-356.5 49</intersection>
<intersection>-339.5 51</intersection>
<intersection>-323.5 53</intersection>
<intersection>-307.5 55</intersection>
<intersection>-291.5 57</intersection>
<intersection>-274.5 59</intersection>
<intersection>-258.5 61</intersection>
<intersection>-242.5 63</intersection>
<intersection>-180.5 64</intersection>
<intersection>-163.5 66</intersection>
<intersection>-147.5 68</intersection>
<intersection>-131.5 70</intersection>
<intersection>-115.5 72</intersection>
<intersection>-98.5 74</intersection>
<intersection>-82.5 76</intersection>
<intersection>-66.5 78</intersection>
<intersection>23.5 79</intersection>
<intersection>204.5 93</intersection>
<intersection>221.5 95</intersection>
<intersection>237.5 97</intersection>
<intersection>253.5 99</intersection>
<intersection>269.5 101</intersection>
<intersection>286.5 103</intersection>
<intersection>302.5 105</intersection>
<intersection>318.5 107</intersection>
<intersection>388 108</intersection>
<intersection>405 110</intersection>
<intersection>421 112</intersection>
<intersection>437 114</intersection>
<intersection>453 116</intersection>
<intersection>470 118</intersection>
<intersection>486 120</intersection>
<intersection>502 122</intersection>
<intersection>523 123</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-889.5,230.5,-889.5</points>
<connection>
<GID>5424</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212.5,-872.5,230.5,-872.5</points>
<connection>
<GID>5422</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>212.5,-840.5,230.5,-840.5</points>
<connection>
<GID>5418</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>212.5,-856.5,230.5,-856.5</points>
<connection>
<GID>5420</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>212.5,-824.5,231.5,-824.5</points>
<connection>
<GID>5439</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>212.5,-807.5,231.5,-807.5</points>
<connection>
<GID>5435</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>212.5,-791.5,231.5,-791.5</points>
<connection>
<GID>5431</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>212.5,-775.5,231.5,-775.5</points>
<connection>
<GID>5429</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>212.5,-715.5,235.5,-715.5</points>
<connection>
<GID>3984</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>212.5,-698.5,235.5,-698.5</points>
<connection>
<GID>3982</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>212.5,-682.5,235.5,-682.5</points>
<connection>
<GID>3980</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>212.5,-666.5,235.5,-666.5</points>
<connection>
<GID>3978</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>212.5,-650.5,236.5,-650.5</points>
<connection>
<GID>3999</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>212.5,-633.5,236.5,-633.5</points>
<connection>
<GID>3995</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>212.5,-617.5,236.5,-617.5</points>
<connection>
<GID>3991</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>212.5,-601.5,236.5,-601.5</points>
<connection>
<GID>3989</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>212.5,-529.5,239.5,-529.5</points>
<connection>
<GID>3504</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>212.5,-512.5,239.5,-512.5</points>
<connection>
<GID>3502</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>212.5,-496.5,239.5,-496.5</points>
<connection>
<GID>3500</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>212.5,-480.5,239.5,-480.5</points>
<connection>
<GID>3498</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>212.5,-464.5,240.5,-464.5</points>
<connection>
<GID>3519</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>212.5,-447.5,240.5,-447.5</points>
<connection>
<GID>3515</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>212.5,-431.5,240.5,-431.5</points>
<connection>
<GID>3511</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>212.5,-415.5,240.5,-415.5</points>
<connection>
<GID>3509</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>212.5,-356.5,236.5,-356.5</points>
<connection>
<GID>3264</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>212.5,-339.5,236.5,-339.5</points>
<connection>
<GID>3262</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>212.5,-323.5,236.5,-323.5</points>
<connection>
<GID>3260</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>212.5,-307.5,236.5,-307.5</points>
<connection>
<GID>3258</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>212.5,-291.5,237.5,-291.5</points>
<connection>
<GID>3279</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>212.5,-274.5,237.5,-274.5</points>
<connection>
<GID>3275</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>212.5,-258.5,237.5,-258.5</points>
<connection>
<GID>3271</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>212.5,-242.5,237.5,-242.5</points>
<connection>
<GID>3269</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>212.5,-180.5,238.5,-180.5</points>
<connection>
<GID>2304</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>212.5,-163.5,238.5,-163.5</points>
<connection>
<GID>2302</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>212.5,-147.5,238.5,-147.5</points>
<connection>
<GID>2300</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>212.5,-131.5,238.5,-131.5</points>
<connection>
<GID>2298</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>212.5,-115.5,239.5,-115.5</points>
<connection>
<GID>2319</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>212.5,-98.5,239.5,-98.5</points>
<connection>
<GID>2315</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>212.5,-82.5,239.5,-82.5</points>
<connection>
<GID>2311</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>212.5,-66.5,239.5,-66.5</points>
<connection>
<GID>2309</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>212.5,23.5,239.5,23.5</points>
<connection>
<GID>4224</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection>
<intersection>218.5 80</intersection></hsegment>
<vsegment>
<ID>80</ID>
<points>218.5,23.5,218.5,137.5</points>
<intersection>23.5 79</intersection>
<intersection>40.5 81</intersection>
<intersection>56.5 83</intersection>
<intersection>72.5 86</intersection>
<intersection>88.5 85</intersection>
<intersection>105.5 88</intersection>
<intersection>121.5 90</intersection>
<intersection>137.5 92</intersection></vsegment>
<hsegment>
<ID>81</ID>
<points>218.5,40.5,239.5,40.5</points>
<connection>
<GID>4222</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>83</ID>
<points>218.5,56.5,239.5,56.5</points>
<connection>
<GID>4220</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>85</ID>
<points>218.5,88.5,240.5,88.5</points>
<connection>
<GID>4239</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>86</ID>
<points>218.5,72.5,239.5,72.5</points>
<connection>
<GID>4218</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>88</ID>
<points>218.5,105.5,240.5,105.5</points>
<connection>
<GID>4235</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>90</ID>
<points>218.5,121.5,240.5,121.5</points>
<connection>
<GID>4231</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>92</ID>
<points>218.5,137.5,240.5,137.5</points>
<connection>
<GID>4229</GID>
<name>IN_0</name></connection>
<intersection>218.5 80</intersection></hsegment>
<hsegment>
<ID>93</ID>
<points>212.5,204.5,234.5,204.5</points>
<connection>
<GID>4944</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>212.5,221.5,234.5,221.5</points>
<connection>
<GID>4942</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>97</ID>
<points>212.5,237.5,234.5,237.5</points>
<connection>
<GID>4940</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>99</ID>
<points>212.5,253.5,234.5,253.5</points>
<connection>
<GID>4938</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>212.5,269.5,235.5,269.5</points>
<connection>
<GID>4959</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>103</ID>
<points>212.5,286.5,235.5,286.5</points>
<connection>
<GID>4955</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>105</ID>
<points>212.5,302.5,235.5,302.5</points>
<connection>
<GID>4951</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>107</ID>
<points>212.5,318.5,235.5,318.5</points>
<connection>
<GID>4949</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>108</ID>
<points>212.5,388,236,388</points>
<connection>
<GID>5664</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>110</ID>
<points>212.5,405,236,405</points>
<connection>
<GID>5662</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>112</ID>
<points>212.5,421,236,421</points>
<connection>
<GID>5660</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>114</ID>
<points>212.5,437,236,437</points>
<connection>
<GID>5658</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>116</ID>
<points>212.5,453,237,453</points>
<connection>
<GID>5679</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>118</ID>
<points>212.5,470,237,470</points>
<connection>
<GID>5675</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>120</ID>
<points>212.5,486,237,486</points>
<connection>
<GID>5671</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>122</ID>
<points>212.5,502,237,502</points>
<connection>
<GID>5669</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>123</ID>
<points>203,523,212.5,523</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,-935,216,505.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-885.5 7</intersection>
<intersection>-868.5 1</intersection>
<intersection>-852.5 3</intersection>
<intersection>-837 4</intersection>
<intersection>-820.5 5</intersection>
<intersection>-803.5 8</intersection>
<intersection>-787.5 9</intersection>
<intersection>-772 10</intersection>
<intersection>-711.5 11</intersection>
<intersection>-694.5 12</intersection>
<intersection>-678.5 13</intersection>
<intersection>-663 14</intersection>
<intersection>-646.5 15</intersection>
<intersection>-629.5 16</intersection>
<intersection>-613.5 17</intersection>
<intersection>-598 18</intersection>
<intersection>-525.5 19</intersection>
<intersection>-508.5 21</intersection>
<intersection>-460.5 26</intersection>
<intersection>-443.5 29</intersection>
<intersection>-427.5 31</intersection>
<intersection>-412 33</intersection>
<intersection>-352.5 34</intersection>
<intersection>-335.5 35</intersection>
<intersection>-319.5 36</intersection>
<intersection>-304 37</intersection>
<intersection>-287.5 38</intersection>
<intersection>-270.5 39</intersection>
<intersection>-254.5 40</intersection>
<intersection>-239 41</intersection>
<intersection>-176.5 42</intersection>
<intersection>-159.5 43</intersection>
<intersection>-143.5 45</intersection>
<intersection>-128 47</intersection>
<intersection>-111.5 48</intersection>
<intersection>-94.5 49</intersection>
<intersection>-78.5 51</intersection>
<intersection>-63 53</intersection>
<intersection>27.5 54</intersection>
<intersection>208.5 69</intersection>
<intersection>225.5 70</intersection>
<intersection>241.5 71</intersection>
<intersection>257 72</intersection>
<intersection>273.5 73</intersection>
<intersection>290.5 74</intersection>
<intersection>306.5 75</intersection>
<intersection>322 76</intersection>
<intersection>392 77</intersection>
<intersection>409 78</intersection>
<intersection>425 79</intersection>
<intersection>440.5 80</intersection>
<intersection>457 81</intersection>
<intersection>474 82</intersection>
<intersection>490 83</intersection>
<intersection>505.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,-868.5,224.5,-868.5</points>
<connection>
<GID>5423</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,505.5,230.5,505.5</points>
<connection>
<GID>5670</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>216,-852.5,224.5,-852.5</points>
<connection>
<GID>5421</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>216,-837,224.5,-837</points>
<connection>
<GID>5419</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>216,-820.5,224.5,-820.5</points>
<connection>
<GID>5441</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>216,-885.5,224.5,-885.5</points>
<connection>
<GID>5425</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>216,-803.5,224.5,-803.5</points>
<connection>
<GID>5437</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>216,-787.5,224.5,-787.5</points>
<connection>
<GID>5433</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>216,-772,225,-772</points>
<connection>
<GID>5430</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>216,-711.5,229.5,-711.5</points>
<connection>
<GID>3985</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>216,-694.5,229.5,-694.5</points>
<connection>
<GID>3983</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>216,-678.5,229.5,-678.5</points>
<connection>
<GID>3981</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>216,-663,229.5,-663</points>
<connection>
<GID>3979</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>216,-646.5,229.5,-646.5</points>
<connection>
<GID>4001</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>216,-629.5,229.5,-629.5</points>
<connection>
<GID>3997</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>216,-613.5,229.5,-613.5</points>
<connection>
<GID>3993</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>216,-598,230,-598</points>
<connection>
<GID>3990</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>216,-525.5,233.5,-525.5</points>
<connection>
<GID>3505</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>216,-508.5,233.5,-508.5</points>
<connection>
<GID>3503</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection>
<intersection>225 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>225,-508.5,225,-460.5</points>
<intersection>-508.5 21</intersection>
<intersection>-492.5 23</intersection>
<intersection>-477 27</intersection>
<intersection>-460.5 26</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>225,-492.5,233.5,-492.5</points>
<connection>
<GID>3501</GID>
<name>IN_1</name></connection>
<intersection>225 22</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>216,-460.5,233.5,-460.5</points>
<connection>
<GID>3521</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection>
<intersection>225 22</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>225,-477,233.5,-477</points>
<connection>
<GID>3499</GID>
<name>IN_1</name></connection>
<intersection>225 22</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>216,-443.5,233.5,-443.5</points>
<connection>
<GID>3517</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>216,-427.5,233.5,-427.5</points>
<connection>
<GID>3513</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>216,-412,234,-412</points>
<connection>
<GID>3510</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>216,-352.5,230.5,-352.5</points>
<connection>
<GID>3265</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>216,-335.5,230.5,-335.5</points>
<connection>
<GID>3263</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>216,-319.5,230.5,-319.5</points>
<connection>
<GID>3261</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>216,-304,230.5,-304</points>
<connection>
<GID>3259</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>216,-287.5,230.5,-287.5</points>
<connection>
<GID>3281</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>216,-270.5,230.5,-270.5</points>
<connection>
<GID>3277</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>216,-254.5,230.5,-254.5</points>
<connection>
<GID>3273</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>216,-239,231,-239</points>
<connection>
<GID>3270</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>216,-176.5,232.5,-176.5</points>
<connection>
<GID>2305</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>216,-159.5,232.5,-159.5</points>
<connection>
<GID>2303</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>216,-143.5,232.5,-143.5</points>
<connection>
<GID>2301</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>216,-128,232.5,-128</points>
<connection>
<GID>2299</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>216,-111.5,232.5,-111.5</points>
<connection>
<GID>2321</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>216,-94.5,232.5,-94.5</points>
<connection>
<GID>2317</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>216,-78.5,232.5,-78.5</points>
<connection>
<GID>2313</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>216,-63,233,-63</points>
<connection>
<GID>2310</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>216,27.5,233.5,27.5</points>
<connection>
<GID>4225</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection>
<intersection>221.5 55</intersection></hsegment>
<vsegment>
<ID>55</ID>
<points>221.5,27.5,221.5,141</points>
<intersection>27.5 54</intersection>
<intersection>44.5 56</intersection>
<intersection>60.5 58</intersection>
<intersection>76 62</intersection>
<intersection>92.5 61</intersection>
<intersection>109.5 64</intersection>
<intersection>125.5 66</intersection>
<intersection>141 68</intersection></vsegment>
<hsegment>
<ID>56</ID>
<points>221.5,44.5,233.5,44.5</points>
<connection>
<GID>4223</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>221.5,60.5,233.5,60.5</points>
<connection>
<GID>4221</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>221.5,92.5,233.5,92.5</points>
<connection>
<GID>4241</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>221.5,76,233.5,76</points>
<connection>
<GID>4219</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>221.5,109.5,233.5,109.5</points>
<connection>
<GID>4237</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>221.5,125.5,233.5,125.5</points>
<connection>
<GID>4233</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>221.5,141,234,141</points>
<connection>
<GID>4230</GID>
<name>IN_1</name></connection>
<intersection>221.5 55</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>216,208.5,228.5,208.5</points>
<connection>
<GID>4945</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>216,225.5,228.5,225.5</points>
<connection>
<GID>4943</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>216,241.5,228.5,241.5</points>
<connection>
<GID>4941</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>216,257,228.5,257</points>
<connection>
<GID>4939</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>216,273.5,228.5,273.5</points>
<connection>
<GID>4961</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>216,290.5,228.5,290.5</points>
<connection>
<GID>4957</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>75</ID>
<points>216,306.5,228.5,306.5</points>
<connection>
<GID>4953</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>216,322,229,322</points>
<connection>
<GID>4950</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>216,392,230,392</points>
<connection>
<GID>5665</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>216,409,230,409</points>
<connection>
<GID>5663</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>216,425,230,425</points>
<connection>
<GID>5661</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>80</ID>
<points>216,440.5,230,440.5</points>
<connection>
<GID>5659</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>81</ID>
<points>216,457,230,457</points>
<connection>
<GID>5681</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>82</ID>
<points>216,474,230,474</points>
<connection>
<GID>5677</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>83</ID>
<points>216,490,230,490</points>
<connection>
<GID>5673</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-909,241.5,-903</points>
<connection>
<GID>5293</GID>
<name>N_in0</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-909,272.5,-903.5</points>
<connection>
<GID>5294</GID>
<name>N_in0</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,-909,304.5,-903.5</points>
<connection>
<GID>5295</GID>
<name>N_in0</name></connection>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-909,335.5,-902.5</points>
<connection>
<GID>5296</GID>
<name>N_in0</name></connection>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365.5,-909,365.5,-901.5</points>
<connection>
<GID>5297</GID>
<name>N_in0</name></connection>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-909,396.5,-901</points>
<connection>
<GID>5298</GID>
<name>N_in0</name></connection>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-909,427.5,-900</points>
<connection>
<GID>5300</GID>
<name>N_in0</name></connection>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-909,458.5,-902</points>
<connection>
<GID>5299</GID>
<name>N_in0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-911.5,225,-904</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-911.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-911.5,456.5,-911.5</points>
<connection>
<GID>47</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>35</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>37</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>39</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>41</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>43</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>45</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>49</GID>
<name>ENABLE_0</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-917,241.5,-914.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-917,272.5,-914.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,-917.5,304.5,-914.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-917.5,335.5,-914.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365.5,-917.5,365.5,-914.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1577</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268.5,-182,270.5,-182</points>
<connection>
<GID>2170</GID>
<name>OUT</name></connection>
<connection>
<GID>2171</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-918,396.5,-914.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-185.5,272.5,-185</points>
<connection>
<GID>2171</GID>
<name>IN_0</name></connection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,-185.5,272.5,-185.5</points>
<intersection>258.5 2</intersection>
<intersection>272.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258.5,-185.5,258.5,-172.5</points>
<intersection>-185.5 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258.5,-181,262.5,-181</points>
<connection>
<GID>2170</GID>
<name>IN_0</name></connection>
<intersection>258.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256.5,-172.5,258.5,-172.5</points>
<connection>
<GID>2172</GID>
<name>OUT_0</name></connection>
<intersection>258.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-918.5,427.5,-914.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-85,481,-85</points>
<connection>
<GID>2362</GID>
<name>IN_1</name></connection>
<connection>
<GID>2365</GID>
<name>IN_1</name></connection>
<connection>
<GID>2368</GID>
<name>IN_1</name></connection>
<connection>
<GID>2371</GID>
<name>IN_1</name></connection>
<connection>
<GID>2374</GID>
<name>IN_1</name></connection>
<connection>
<GID>2377</GID>
<name>IN_1</name></connection>
<connection>
<GID>2380</GID>
<name>IN_1</name></connection>
<connection>
<GID>2383</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-85,245,-82.5</points>
<connection>
<GID>2311</GID>
<name>OUT_0</name></connection>
<intersection>-85 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-918.5,458.5,-914.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-77.5,468.5,-77.5</points>
<connection>
<GID>2313</GID>
<name>OUT</name></connection>
<connection>
<GID>2364</GID>
<name>clock</name></connection>
<connection>
<GID>2367</GID>
<name>clock</name></connection>
<connection>
<GID>2370</GID>
<name>clock</name></connection>
<connection>
<GID>2373</GID>
<name>clock</name></connection>
<connection>
<GID>2376</GID>
<name>clock</name></connection>
<connection>
<GID>2379</GID>
<name>clock</name></connection>
<connection>
<GID>2382</GID>
<name>clock</name></connection>
<connection>
<GID>2385</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-101,480.5,-101</points>
<connection>
<GID>2338</GID>
<name>IN_1</name></connection>
<connection>
<GID>2341</GID>
<name>IN_1</name></connection>
<connection>
<GID>2344</GID>
<name>IN_1</name></connection>
<connection>
<GID>2347</GID>
<name>IN_1</name></connection>
<connection>
<GID>2350</GID>
<name>IN_1</name></connection>
<connection>
<GID>2353</GID>
<name>IN_1</name></connection>
<connection>
<GID>2356</GID>
<name>IN_1</name></connection>
<connection>
<GID>2359</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-101,245,-98.5</points>
<connection>
<GID>2315</GID>
<name>OUT_0</name></connection>
<intersection>-101 1</intersection></vsegment></shape></wire>
<wire>
<ID>1582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-93.5,468,-93.5</points>
<connection>
<GID>2317</GID>
<name>OUT</name></connection>
<connection>
<GID>2340</GID>
<name>clock</name></connection>
<connection>
<GID>2343</GID>
<name>clock</name></connection>
<connection>
<GID>2346</GID>
<name>clock</name></connection>
<connection>
<GID>2349</GID>
<name>clock</name></connection>
<connection>
<GID>2352</GID>
<name>clock</name></connection>
<connection>
<GID>2355</GID>
<name>clock</name></connection>
<connection>
<GID>2358</GID>
<name>clock</name></connection>
<connection>
<GID>2361</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-110.5,467.5,-110.5</points>
<connection>
<GID>2337</GID>
<name>clock</name></connection>
<connection>
<GID>2334</GID>
<name>clock</name></connection>
<connection>
<GID>2331</GID>
<name>clock</name></connection>
<connection>
<GID>2328</GID>
<name>clock</name></connection>
<connection>
<GID>2325</GID>
<name>clock</name></connection>
<connection>
<GID>2322</GID>
<name>clock</name></connection>
<connection>
<GID>2321</GID>
<name>OUT</name></connection>
<connection>
<GID>2316</GID>
<name>clock</name></connection>
<connection>
<GID>2308</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-827.5,184,452.5</points>
<intersection>-827.5 1</intersection>
<intersection>-653.5 8</intersection>
<intersection>-467.5 7</intersection>
<intersection>-294.5 6</intersection>
<intersection>-118.5 5</intersection>
<intersection>85.5 4</intersection>
<intersection>266.5 3</intersection>
<intersection>450 2</intersection>
<intersection>452.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-827.5,188.5,-827.5</points>
<connection>
<GID>5417</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,450,194,450</points>
<connection>
<GID>5657</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184,266.5,192.5,266.5</points>
<connection>
<GID>4937</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>184,85.5,197.5,85.5</points>
<connection>
<GID>4217</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>184,-118.5,196.5,-118.5</points>
<connection>
<GID>2297</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>184,-294.5,194.5,-294.5</points>
<connection>
<GID>3257</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>184,-467.5,197.5,-467.5</points>
<connection>
<GID>3497</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>184,-653.5,193.5,-653.5</points>
<connection>
<GID>3977</GID>
<name>IN_2</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>138.5,452.5,184,452.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>1584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-118,480,-118</points>
<connection>
<GID>2306</GID>
<name>IN_1</name></connection>
<connection>
<GID>2312</GID>
<name>IN_1</name></connection>
<connection>
<GID>2318</GID>
<name>IN_1</name></connection>
<connection>
<GID>2323</GID>
<name>IN_1</name></connection>
<connection>
<GID>2326</GID>
<name>IN_1</name></connection>
<connection>
<GID>2329</GID>
<name>IN_1</name></connection>
<connection>
<GID>2332</GID>
<name>IN_1</name></connection>
<connection>
<GID>2335</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-118,245,-115.5</points>
<connection>
<GID>2319</GID>
<name>OUT_0</name></connection>
<intersection>-118 1</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-828.5,182,449</points>
<intersection>-828.5 1</intersection>
<intersection>-654.5 3</intersection>
<intersection>-468.5 4</intersection>
<intersection>-295.5 5</intersection>
<intersection>-119.5 6</intersection>
<intersection>84.5 7</intersection>
<intersection>265.5 8</intersection>
<intersection>449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>182,-828.5,188.5,-828.5</points>
<connection>
<GID>5417</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,449,194,449</points>
<connection>
<GID>5657</GID>
<name>IN_1</name></connection>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>182,-654.5,193.5,-654.5</points>
<connection>
<GID>3977</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>182,-468.5,197.5,-468.5</points>
<connection>
<GID>3497</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182,-295.5,194.5,-295.5</points>
<connection>
<GID>3257</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>182,-119.5,196.5,-119.5</points>
<connection>
<GID>2297</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>182,84.5,197.5,84.5</points>
<connection>
<GID>4217</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>182,265.5,192.5,265.5</points>
<connection>
<GID>4937</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>1585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-127,468,-127</points>
<connection>
<GID>2299</GID>
<name>OUT</name></connection>
<connection>
<GID>2276</GID>
<name>clock</name></connection>
<connection>
<GID>2273</GID>
<name>clock</name></connection>
<connection>
<GID>2270</GID>
<name>clock</name></connection>
<connection>
<GID>2267</GID>
<name>clock</name></connection>
<connection>
<GID>2264</GID>
<name>clock</name></connection>
<connection>
<GID>2261</GID>
<name>clock</name></connection>
<connection>
<GID>2258</GID>
<name>clock</name></connection>
<connection>
<GID>2255</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-829.5,179,445.5</points>
<intersection>-829.5 1</intersection>
<intersection>-655.5 3</intersection>
<intersection>-469.5 4</intersection>
<intersection>-296.5 5</intersection>
<intersection>-120.5 6</intersection>
<intersection>83.5 7</intersection>
<intersection>264.5 8</intersection>
<intersection>445.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179,-829.5,188.5,-829.5</points>
<connection>
<GID>5417</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,445.5,186,445.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>179 0</intersection>
<intersection>186 13</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>179,-655.5,193.5,-655.5</points>
<connection>
<GID>3977</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>179,-469.5,197.5,-469.5</points>
<connection>
<GID>3497</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>179,-296.5,194.5,-296.5</points>
<connection>
<GID>3257</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>179,-120.5,196.5,-120.5</points>
<connection>
<GID>2297</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>179,83.5,197.5,83.5</points>
<connection>
<GID>4217</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>179,264.5,192.5,264.5</points>
<connection>
<GID>4937</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>186,445.5,186,448</points>
<intersection>445.5 2</intersection>
<intersection>448 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>186,448,194,448</points>
<connection>
<GID>5657</GID>
<name>IN_0</name></connection>
<intersection>186 13</intersection></hsegment></shape></wire>
<wire>
<ID>1586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-134.5,480.5,-134.5</points>
<connection>
<GID>2253</GID>
<name>IN_1</name></connection>
<connection>
<GID>2256</GID>
<name>IN_1</name></connection>
<connection>
<GID>2259</GID>
<name>IN_1</name></connection>
<connection>
<GID>2262</GID>
<name>IN_1</name></connection>
<connection>
<GID>2265</GID>
<name>IN_1</name></connection>
<connection>
<GID>2268</GID>
<name>IN_1</name></connection>
<connection>
<GID>2271</GID>
<name>IN_1</name></connection>
<connection>
<GID>2274</GID>
<name>IN_1</name></connection>
<intersection>244 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>244,-134.5,244,-131.5</points>
<connection>
<GID>2298</GID>
<name>OUT_0</name></connection>
<intersection>-134.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-142.5,467.5,-142.5</points>
<connection>
<GID>2301</GID>
<name>OUT</name></connection>
<connection>
<GID>2252</GID>
<name>clock</name></connection>
<connection>
<GID>2249</GID>
<name>clock</name></connection>
<connection>
<GID>2246</GID>
<name>clock</name></connection>
<connection>
<GID>2243</GID>
<name>clock</name></connection>
<connection>
<GID>2240</GID>
<name>clock</name></connection>
<connection>
<GID>2237</GID>
<name>clock</name></connection>
<connection>
<GID>2234</GID>
<name>clock</name></connection>
<connection>
<GID>2231</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1588</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-150,480,-150</points>
<connection>
<GID>2229</GID>
<name>IN_1</name></connection>
<connection>
<GID>2232</GID>
<name>IN_1</name></connection>
<connection>
<GID>2235</GID>
<name>IN_1</name></connection>
<connection>
<GID>2238</GID>
<name>IN_1</name></connection>
<connection>
<GID>2241</GID>
<name>IN_1</name></connection>
<connection>
<GID>2244</GID>
<name>IN_1</name></connection>
<connection>
<GID>2247</GID>
<name>IN_1</name></connection>
<connection>
<GID>2250</GID>
<name>IN_1</name></connection>
<intersection>244 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>244,-150,244,-147.5</points>
<connection>
<GID>2300</GID>
<name>OUT_0</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>1589</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>300,-182,302,-182</points>
<connection>
<GID>2184</GID>
<name>OUT</name></connection>
<connection>
<GID>2185</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1590</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-185,304,-185</points>
<connection>
<GID>2185</GID>
<name>IN_0</name></connection>
<intersection>290 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>290,-185,290,-172.5</points>
<intersection>-185 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>290,-181,294,-181</points>
<connection>
<GID>2184</GID>
<name>IN_0</name></connection>
<intersection>290 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287.5,-172.5,290,-172.5</points>
<connection>
<GID>2186</GID>
<name>OUT_0</name></connection>
<intersection>290 2</intersection></hsegment></shape></wire>
<wire>
<ID>1591</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330.5,-182,332.5,-182</points>
<connection>
<GID>2187</GID>
<name>OUT</name></connection>
<connection>
<GID>2188</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,-185.5,334.5,-185</points>
<connection>
<GID>2188</GID>
<name>IN_0</name></connection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-185.5,334.5,-185.5</points>
<intersection>320.5 2</intersection>
<intersection>334.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320.5,-185.5,320.5,-172.5</points>
<intersection>-185.5 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320.5,-181,324.5,-181</points>
<connection>
<GID>2187</GID>
<name>IN_0</name></connection>
<intersection>320.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318.5,-172.5,320.5,-172.5</points>
<connection>
<GID>2189</GID>
<name>OUT_0</name></connection>
<intersection>320.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1593</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>362,-182,364,-182</points>
<connection>
<GID>2190</GID>
<name>OUT</name></connection>
<connection>
<GID>2191</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>352,-185,366,-185</points>
<connection>
<GID>2191</GID>
<name>IN_0</name></connection>
<intersection>352 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>352,-185,352,-172.5</points>
<intersection>-185 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>352,-181,356,-181</points>
<connection>
<GID>2190</GID>
<name>IN_0</name></connection>
<intersection>352 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>349.5,-172.5,352,-172.5</points>
<connection>
<GID>2192</GID>
<name>OUT_0</name></connection>
<intersection>352 2</intersection></hsegment></shape></wire>
<wire>
<ID>1595</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391.5,-182,393.5,-182</points>
<connection>
<GID>2193</GID>
<name>OUT</name></connection>
<connection>
<GID>2194</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395.5,-185.5,395.5,-185</points>
<connection>
<GID>2194</GID>
<name>IN_0</name></connection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381.5,-185.5,395.5,-185.5</points>
<intersection>381.5 2</intersection>
<intersection>395.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381.5,-185.5,381.5,-172.5</points>
<intersection>-185.5 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381.5,-181,385.5,-181</points>
<connection>
<GID>2193</GID>
<name>IN_0</name></connection>
<intersection>381.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379.5,-172.5,381.5,-172.5</points>
<connection>
<GID>2195</GID>
<name>OUT_0</name></connection>
<intersection>381.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1597</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>423,-182,425,-182</points>
<connection>
<GID>2196</GID>
<name>OUT</name></connection>
<connection>
<GID>2197</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1598</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413,-185,427,-185</points>
<connection>
<GID>2197</GID>
<name>IN_0</name></connection>
<intersection>413 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>413,-185,413,-172.5</points>
<intersection>-185 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>413,-181,417,-181</points>
<connection>
<GID>2196</GID>
<name>IN_0</name></connection>
<intersection>413 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410.5,-172.5,413,-172.5</points>
<connection>
<GID>2198</GID>
<name>OUT_0</name></connection>
<intersection>413 2</intersection></hsegment></shape></wire>
<wire>
<ID>1599</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453.5,-182,455.5,-182</points>
<connection>
<GID>2199</GID>
<name>OUT</name></connection>
<connection>
<GID>2200</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,-185.5,457.5,-185</points>
<connection>
<GID>2200</GID>
<name>IN_0</name></connection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443.5,-185.5,457.5,-185.5</points>
<intersection>443.5 2</intersection>
<intersection>457.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443.5,-185.5,443.5,-172.5</points>
<intersection>-185.5 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443.5,-181,447.5,-181</points>
<connection>
<GID>2199</GID>
<name>IN_0</name></connection>
<intersection>443.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441.5,-172.5,443.5,-172.5</points>
<connection>
<GID>2201</GID>
<name>OUT_0</name></connection>
<intersection>443.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1601</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>485,-182,487,-182</points>
<connection>
<GID>2202</GID>
<name>OUT</name></connection>
<connection>
<GID>2203</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1602</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475,-185,489,-185</points>
<connection>
<GID>2203</GID>
<name>IN_0</name></connection>
<intersection>475 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>475,-185,475,-172.5</points>
<intersection>-185 1</intersection>
<intersection>-181 4</intersection>
<intersection>-172.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>475,-181,479,-181</points>
<connection>
<GID>2202</GID>
<name>IN_0</name></connection>
<intersection>475 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472.5,-172.5,475,-172.5</points>
<connection>
<GID>2204</GID>
<name>OUT_0</name></connection>
<intersection>475 2</intersection></hsegment></shape></wire>
<wire>
<ID>1603</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>269,-165,271,-165</points>
<connection>
<GID>2205</GID>
<name>OUT</name></connection>
<connection>
<GID>2206</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-168.5,273,-168</points>
<connection>
<GID>2206</GID>
<name>IN_0</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259,-168.5,273,-168.5</points>
<intersection>259 2</intersection>
<intersection>273 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>259,-168.5,259,-155.5</points>
<intersection>-168.5 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259,-164,263,-164</points>
<connection>
<GID>2205</GID>
<name>IN_0</name></connection>
<intersection>259 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>257,-155.5,259,-155.5</points>
<connection>
<GID>2207</GID>
<name>OUT_0</name></connection>
<intersection>259 2</intersection></hsegment></shape></wire>
<wire>
<ID>1605</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>300.5,-165,302.5,-165</points>
<connection>
<GID>2208</GID>
<name>OUT</name></connection>
<connection>
<GID>2209</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,442.5,161.5,442.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>161.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>161.5,442.5,161.5,442.5</points>
<connection>
<GID>122</GID>
<name>ENABLE</name></connection>
<intersection>442.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1606</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-168,304.5,-168</points>
<connection>
<GID>2209</GID>
<name>IN_0</name></connection>
<intersection>290.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>290.5,-168,290.5,-155.5</points>
<intersection>-168 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>290.5,-164,294.5,-164</points>
<connection>
<GID>2208</GID>
<name>IN_0</name></connection>
<intersection>290.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>288,-155.5,290.5,-155.5</points>
<connection>
<GID>2210</GID>
<name>OUT_0</name></connection>
<intersection>290.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138.5,440,161.5,440</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>161.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>161.5,437.5,161.5,440</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>440 1</intersection></vsegment></shape></wire>
<wire>
<ID>1607</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>331,-165,333,-165</points>
<connection>
<GID>2211</GID>
<name>OUT</name></connection>
<connection>
<GID>2212</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138.5,436,161.5,436</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>161.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>161.5,436,161.5,436.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>436 1</intersection></vsegment></shape></wire>
<wire>
<ID>1608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-168.5,335,-168</points>
<connection>
<GID>2212</GID>
<name>IN_0</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,-168.5,335,-168.5</points>
<intersection>321 2</intersection>
<intersection>335 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321,-168.5,321,-155.5</points>
<intersection>-168.5 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321,-164,325,-164</points>
<connection>
<GID>2211</GID>
<name>IN_0</name></connection>
<intersection>321 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>319,-155.5,321,-155.5</points>
<connection>
<GID>2213</GID>
<name>OUT_0</name></connection>
<intersection>321 2</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,432,161.5,435.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>432 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,432,161.5,432</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1609</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>362.5,-165,364.5,-165</points>
<connection>
<GID>2214</GID>
<name>OUT</name></connection>
<connection>
<GID>2215</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,455,194,455</points>
<connection>
<GID>5657</GID>
<name>ENABLE</name></connection>
<intersection>192 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>192,442.5,192,455</points>
<intersection>442.5 4</intersection>
<intersection>455 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>167.5,442.5,192,442.5</points>
<connection>
<GID>122</GID>
<name>OUT_7</name></connection>
<intersection>192 3</intersection></hsegment></shape></wire>
<wire>
<ID>1610</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>352.5,-168,366.5,-168</points>
<connection>
<GID>2215</GID>
<name>IN_0</name></connection>
<intersection>352.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>352.5,-168,352.5,-155.5</points>
<intersection>-168 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>352.5,-164,356.5,-164</points>
<connection>
<GID>2214</GID>
<name>IN_0</name></connection>
<intersection>352.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>350,-155.5,352.5,-155.5</points>
<connection>
<GID>2216</GID>
<name>OUT_0</name></connection>
<intersection>352.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,271.5,192,441.5</points>
<intersection>271.5 1</intersection>
<intersection>441.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,271.5,192.5,271.5</points>
<connection>
<GID>4937</GID>
<name>ENABLE</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167.5,441.5,192,441.5</points>
<connection>
<GID>122</GID>
<name>OUT_6</name></connection>
<intersection>192 0</intersection></hsegment></shape></wire>
<wire>
<ID>1611</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>392,-165,394,-165</points>
<connection>
<GID>2217</GID>
<name>OUT</name></connection>
<connection>
<GID>2218</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,90.5,191,440.5</points>
<intersection>90.5 1</intersection>
<intersection>440.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,90.5,197.5,90.5</points>
<connection>
<GID>4217</GID>
<name>ENABLE</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167.5,440.5,191,440.5</points>
<connection>
<GID>122</GID>
<name>OUT_5</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>1612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396,-168.5,396,-168</points>
<connection>
<GID>2218</GID>
<name>IN_0</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382,-168.5,396,-168.5</points>
<intersection>382 2</intersection>
<intersection>396 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>382,-168.5,382,-155.5</points>
<intersection>-168.5 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>382,-164,386,-164</points>
<connection>
<GID>2217</GID>
<name>IN_0</name></connection>
<intersection>382 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380,-155.5,382,-155.5</points>
<connection>
<GID>2219</GID>
<name>OUT_0</name></connection>
<intersection>382 2</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-113.5,187.5,439.5</points>
<intersection>-113.5 1</intersection>
<intersection>439.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,-113.5,196.5,-113.5</points>
<connection>
<GID>2297</GID>
<name>ENABLE</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167.5,439.5,187.5,439.5</points>
<connection>
<GID>122</GID>
<name>OUT_4</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1613</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>423.5,-165,425.5,-165</points>
<connection>
<GID>2220</GID>
<name>OUT</name></connection>
<connection>
<GID>2221</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-289.5,176.5,438.5</points>
<intersection>-289.5 2</intersection>
<intersection>438.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,438.5,176.5,438.5</points>
<connection>
<GID>122</GID>
<name>OUT_3</name></connection>
<intersection>176.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176.5,-289.5,194.5,-289.5</points>
<connection>
<GID>3257</GID>
<name>ENABLE</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1614</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413.5,-168,427.5,-168</points>
<connection>
<GID>2221</GID>
<name>IN_0</name></connection>
<intersection>413.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>413.5,-168,413.5,-155.5</points>
<intersection>-168 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>413.5,-164,417.5,-164</points>
<connection>
<GID>2220</GID>
<name>IN_0</name></connection>
<intersection>413.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411,-155.5,413.5,-155.5</points>
<connection>
<GID>2222</GID>
<name>OUT_0</name></connection>
<intersection>413.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1615</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>454,-165,456,-165</points>
<connection>
<GID>2223</GID>
<name>OUT</name></connection>
<connection>
<GID>2224</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-462.5,176,437.5</points>
<intersection>-462.5 2</intersection>
<intersection>437.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,437.5,176,437.5</points>
<connection>
<GID>122</GID>
<name>OUT_2</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176,-462.5,197.5,-462.5</points>
<connection>
<GID>3497</GID>
<name>ENABLE</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>1616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,-168.5,458,-168</points>
<connection>
<GID>2224</GID>
<name>IN_0</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444,-168.5,458,-168.5</points>
<intersection>444 2</intersection>
<intersection>458 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>444,-168.5,444,-155.5</points>
<intersection>-168.5 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>444,-164,448,-164</points>
<connection>
<GID>2223</GID>
<name>IN_0</name></connection>
<intersection>444 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>442,-155.5,444,-155.5</points>
<connection>
<GID>2225</GID>
<name>OUT_0</name></connection>
<intersection>444 2</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,-648.5,177.5,436.5</points>
<intersection>-648.5 1</intersection>
<intersection>436.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177.5,-648.5,193.5,-648.5</points>
<connection>
<GID>3977</GID>
<name>ENABLE</name></connection>
<intersection>177.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167.5,436.5,177.5,436.5</points>
<connection>
<GID>122</GID>
<name>OUT_1</name></connection>
<intersection>177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1617</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>485.5,-165,487.5,-165</points>
<connection>
<GID>2226</GID>
<name>OUT</name></connection>
<connection>
<GID>2227</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-822.5,174,435.5</points>
<intersection>-822.5 2</intersection>
<intersection>435.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,435.5,174,435.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-822.5,188.5,-822.5</points>
<connection>
<GID>5417</GID>
<name>ENABLE</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>1618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475.5,-168,489.5,-168</points>
<connection>
<GID>2227</GID>
<name>IN_0</name></connection>
<intersection>475.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>475.5,-168,475.5,-155.5</points>
<intersection>-168 1</intersection>
<intersection>-164 4</intersection>
<intersection>-155.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>475.5,-164,479.5,-164</points>
<connection>
<GID>2226</GID>
<name>IN_0</name></connection>
<intersection>475.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>473,-155.5,475.5,-155.5</points>
<connection>
<GID>2228</GID>
<name>OUT_0</name></connection>
<intersection>475.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,449.5,119.5,449.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1619</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>269.5,-149,271.5,-149</points>
<connection>
<GID>2229</GID>
<name>OUT</name></connection>
<connection>
<GID>2230</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115.5,441,119,441</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,-152.5,273.5,-152</points>
<connection>
<GID>2230</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-152.5,273.5,-152.5</points>
<intersection>259.5 2</intersection>
<intersection>273.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>259.5,-152.5,259.5,-139.5</points>
<intersection>-152.5 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,-148,263.5,-148</points>
<connection>
<GID>2229</GID>
<name>IN_0</name></connection>
<intersection>259.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>257.5,-139.5,259.5,-139.5</points>
<connection>
<GID>2231</GID>
<name>OUT_0</name></connection>
<intersection>259.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,433.5,118.5,433.5</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>118.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>118.5,433.5,118.5,433.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>433.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1621</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301,-149,303,-149</points>
<connection>
<GID>2232</GID>
<name>OUT</name></connection>
<connection>
<GID>2233</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,462,124,466</points>
<connection>
<GID>147</GID>
<name>N_in3</name></connection>
<connection>
<GID>156</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291,-152,305,-152</points>
<connection>
<GID>2233</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291,-152,291,-139.5</points>
<intersection>-152 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291,-148,295,-148</points>
<connection>
<GID>2232</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>288.5,-139.5,291,-139.5</points>
<connection>
<GID>2234</GID>
<name>OUT_0</name></connection>
<intersection>291 2</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,462,134.5,466</points>
<connection>
<GID>148</GID>
<name>N_in3</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1623</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>331.5,-149,333.5,-149</points>
<connection>
<GID>2235</GID>
<name>OUT</name></connection>
<connection>
<GID>2236</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,462,144.5,466</points>
<connection>
<GID>149</GID>
<name>N_in3</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-152.5,335.5,-152</points>
<connection>
<GID>2236</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-152.5,335.5,-152.5</points>
<intersection>321.5 2</intersection>
<intersection>335.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321.5,-152.5,321.5,-139.5</points>
<intersection>-152.5 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321.5,-148,325.5,-148</points>
<connection>
<GID>2235</GID>
<name>IN_0</name></connection>
<intersection>321.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>319.5,-139.5,321.5,-139.5</points>
<connection>
<GID>2237</GID>
<name>OUT_0</name></connection>
<intersection>321.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,462,152,466</points>
<connection>
<GID>150</GID>
<name>N_in3</name></connection>
<connection>
<GID>159</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1625</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363,-149,365,-149</points>
<connection>
<GID>2238</GID>
<name>OUT</name></connection>
<connection>
<GID>2239</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,462,163.5,466</points>
<connection>
<GID>151</GID>
<name>N_in3</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353,-152,367,-152</points>
<connection>
<GID>2239</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353,-152,353,-139.5</points>
<intersection>-152 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353,-148,357,-148</points>
<connection>
<GID>2238</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>350.5,-139.5,353,-139.5</points>
<connection>
<GID>2240</GID>
<name>OUT_0</name></connection>
<intersection>353 2</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,462,172.5,466</points>
<connection>
<GID>153</GID>
<name>N_in3</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1627</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>392.5,-149,394.5,-149</points>
<connection>
<GID>2241</GID>
<name>OUT</name></connection>
<connection>
<GID>2242</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,462,182.5,466</points>
<connection>
<GID>152</GID>
<name>N_in3</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-152.5,396.5,-152</points>
<connection>
<GID>2242</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382.5,-152.5,396.5,-152.5</points>
<intersection>382.5 2</intersection>
<intersection>396.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>382.5,-152.5,382.5,-139.5</points>
<intersection>-152.5 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>382.5,-148,386.5,-148</points>
<connection>
<GID>2241</GID>
<name>IN_0</name></connection>
<intersection>382.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380.5,-139.5,382.5,-139.5</points>
<connection>
<GID>2243</GID>
<name>OUT_0</name></connection>
<intersection>382.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,462,190.5,466</points>
<connection>
<GID>154</GID>
<name>N_in3</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1629</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424,-149,426,-149</points>
<connection>
<GID>2244</GID>
<name>OUT</name></connection>
<connection>
<GID>2245</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,478,124,481</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<connection>
<GID>173</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1630</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414,-152,428,-152</points>
<connection>
<GID>2245</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414,-152,414,-139.5</points>
<intersection>-152 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414,-148,418,-148</points>
<connection>
<GID>2244</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411.5,-139.5,414,-139.5</points>
<connection>
<GID>2246</GID>
<name>OUT_0</name></connection>
<intersection>414 2</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,478,144,481</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1631</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>454.5,-149,456.5,-149</points>
<connection>
<GID>2247</GID>
<name>OUT</name></connection>
<connection>
<GID>2248</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-152.5,458.5,-152</points>
<connection>
<GID>2248</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,-152.5,458.5,-152.5</points>
<intersection>444.5 2</intersection>
<intersection>458.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>444.5,-152.5,444.5,-139.5</points>
<intersection>-152.5 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>444.5,-148,448.5,-148</points>
<connection>
<GID>2247</GID>
<name>IN_0</name></connection>
<intersection>444.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>442.5,-139.5,444.5,-139.5</points>
<connection>
<GID>2249</GID>
<name>OUT_0</name></connection>
<intersection>444.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,478,163,481</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1633</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486,-149,488,-149</points>
<connection>
<GID>2250</GID>
<name>OUT</name></connection>
<connection>
<GID>2251</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,478,172.5,481</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1634</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476,-152,490,-152</points>
<connection>
<GID>2251</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476,-152,476,-139.5</points>
<intersection>-152 1</intersection>
<intersection>-148 4</intersection>
<intersection>-139.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476,-148,480,-148</points>
<connection>
<GID>2250</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>473.5,-139.5,476,-139.5</points>
<connection>
<GID>2252</GID>
<name>OUT_0</name></connection>
<intersection>476 2</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,478,182,481</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>481 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>182,481,182.5,481</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>1635</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270,-133.5,272,-133.5</points>
<connection>
<GID>2253</GID>
<name>OUT</name></connection>
<connection>
<GID>2254</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,478,190.5,481</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-137,274,-136.5</points>
<connection>
<GID>2254</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-137,274,-137</points>
<intersection>260 2</intersection>
<intersection>274 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260,-137,260,-124</points>
<intersection>-137 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260,-132.5,264,-132.5</points>
<connection>
<GID>2253</GID>
<name>IN_0</name></connection>
<intersection>260 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258,-124,260,-124</points>
<connection>
<GID>2255</GID>
<name>OUT_0</name></connection>
<intersection>260 2</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,478,133.5,481</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>481 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,481,134,481</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>355,496.5,355,509.5</points>
<intersection>496.5 1</intersection>
<intersection>509.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,496.5,366,496.5</points>
<intersection>355 0</intersection>
<intersection>356 4</intersection>
<intersection>366 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,509.5,355,509.5</points>
<connection>
<GID>5757</GID>
<name>OUT_0</name></connection>
<intersection>355 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>366,496.5,366,497</points>
<connection>
<GID>5756</GID>
<name>IN_0</name></connection>
<intersection>496.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>356,496.5,356,501</points>
<connection>
<GID>5755</GID>
<name>IN_0</name></connection>
<intersection>496.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1637</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,-133.5,303.5,-133.5</points>
<connection>
<GID>2256</GID>
<name>OUT</name></connection>
<connection>
<GID>2257</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,-136.5,305.5,-136.5</points>
<connection>
<GID>2257</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291.5,-136.5,291.5,-124</points>
<intersection>-136.5 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291.5,-132.5,295.5,-132.5</points>
<connection>
<GID>2256</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289,-124,291.5,-124</points>
<connection>
<GID>2258</GID>
<name>OUT_0</name></connection>
<intersection>291.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1639</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332,-133.5,334,-133.5</points>
<connection>
<GID>2259</GID>
<name>OUT</name></connection>
<connection>
<GID>2260</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,-137,336,-136.5</points>
<connection>
<GID>2260</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-137,336,-137</points>
<intersection>322 2</intersection>
<intersection>336 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322,-137,322,-124</points>
<intersection>-137 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322,-132.5,326,-132.5</points>
<connection>
<GID>2259</GID>
<name>IN_0</name></connection>
<intersection>322 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320,-124,322,-124</points>
<connection>
<GID>2261</GID>
<name>OUT_0</name></connection>
<intersection>322 2</intersection></hsegment></shape></wire>
<wire>
<ID>1641</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363.5,-133.5,365.5,-133.5</points>
<connection>
<GID>2262</GID>
<name>OUT</name></connection>
<connection>
<GID>2263</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1642</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353.5,-136.5,367.5,-136.5</points>
<connection>
<GID>2263</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353.5,-136.5,353.5,-124</points>
<intersection>-136.5 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353.5,-132.5,357.5,-132.5</points>
<connection>
<GID>2262</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351,-124,353.5,-124</points>
<connection>
<GID>2264</GID>
<name>OUT_0</name></connection>
<intersection>353.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1643</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393,-133.5,395,-133.5</points>
<connection>
<GID>2265</GID>
<name>OUT</name></connection>
<connection>
<GID>2266</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,-137,397,-136.5</points>
<connection>
<GID>2266</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383,-137,397,-137</points>
<intersection>383 2</intersection>
<intersection>397 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,-137,383,-124</points>
<intersection>-137 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383,-132.5,387,-132.5</points>
<connection>
<GID>2265</GID>
<name>IN_0</name></connection>
<intersection>383 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381,-124,383,-124</points>
<connection>
<GID>2267</GID>
<name>OUT_0</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>1645</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424.5,-133.5,426.5,-133.5</points>
<connection>
<GID>2268</GID>
<name>OUT</name></connection>
<connection>
<GID>2269</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414.5,-136.5,428.5,-136.5</points>
<connection>
<GID>2269</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414.5,-136.5,414.5,-124</points>
<intersection>-136.5 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414.5,-132.5,418.5,-132.5</points>
<connection>
<GID>2268</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412,-124,414.5,-124</points>
<connection>
<GID>2270</GID>
<name>OUT_0</name></connection>
<intersection>414.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1647</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455,-133.5,457,-133.5</points>
<connection>
<GID>2271</GID>
<name>OUT</name></connection>
<connection>
<GID>2272</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-137,459,-136.5</points>
<connection>
<GID>2272</GID>
<name>IN_0</name></connection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,-137,459,-137</points>
<intersection>445 2</intersection>
<intersection>459 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445,-137,445,-124</points>
<intersection>-137 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445,-132.5,449,-132.5</points>
<connection>
<GID>2271</GID>
<name>IN_0</name></connection>
<intersection>445 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443,-124,445,-124</points>
<connection>
<GID>2273</GID>
<name>OUT_0</name></connection>
<intersection>445 2</intersection></hsegment></shape></wire>
<wire>
<ID>1649</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486.5,-133.5,488.5,-133.5</points>
<connection>
<GID>2274</GID>
<name>OUT</name></connection>
<connection>
<GID>2275</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476.5,-136.5,490.5,-136.5</points>
<connection>
<GID>2275</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476.5,-136.5,476.5,-124</points>
<intersection>-136.5 1</intersection>
<intersection>-132.5 4</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476.5,-132.5,480.5,-132.5</points>
<connection>
<GID>2274</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474,-124,476.5,-124</points>
<connection>
<GID>2276</GID>
<name>OUT_0</name></connection>
<intersection>476.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-158.5,467,-158.5</points>
<connection>
<GID>2303</GID>
<name>OUT</name></connection>
<connection>
<GID>2228</GID>
<name>clock</name></connection>
<connection>
<GID>2225</GID>
<name>clock</name></connection>
<connection>
<GID>2222</GID>
<name>clock</name></connection>
<connection>
<GID>2219</GID>
<name>clock</name></connection>
<connection>
<GID>2216</GID>
<name>clock</name></connection>
<connection>
<GID>2213</GID>
<name>clock</name></connection>
<connection>
<GID>2210</GID>
<name>clock</name></connection>
<connection>
<GID>2207</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1652</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-166,479.5,-166</points>
<connection>
<GID>2205</GID>
<name>IN_1</name></connection>
<connection>
<GID>2208</GID>
<name>IN_1</name></connection>
<connection>
<GID>2211</GID>
<name>IN_1</name></connection>
<connection>
<GID>2214</GID>
<name>IN_1</name></connection>
<connection>
<GID>2217</GID>
<name>IN_1</name></connection>
<connection>
<GID>2220</GID>
<name>IN_1</name></connection>
<connection>
<GID>2223</GID>
<name>IN_1</name></connection>
<connection>
<GID>2226</GID>
<name>IN_1</name></connection>
<intersection>244 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>244,-166,244,-163.5</points>
<connection>
<GID>2302</GID>
<name>OUT_0</name></connection>
<intersection>-166 1</intersection></vsegment></shape></wire>
<wire>
<ID>1653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-175.5,466.5,-175.5</points>
<connection>
<GID>2305</GID>
<name>OUT</name></connection>
<connection>
<GID>2204</GID>
<name>clock</name></connection>
<connection>
<GID>2201</GID>
<name>clock</name></connection>
<connection>
<GID>2198</GID>
<name>clock</name></connection>
<connection>
<GID>2195</GID>
<name>clock</name></connection>
<connection>
<GID>2192</GID>
<name>clock</name></connection>
<connection>
<GID>2189</GID>
<name>clock</name></connection>
<connection>
<GID>2186</GID>
<name>clock</name></connection>
<connection>
<GID>2172</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-183,245,-180.5</points>
<intersection>-183 2</intersection>
<intersection>-180.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>245,-183,479,-183</points>
<connection>
<GID>2170</GID>
<name>IN_1</name></connection>
<connection>
<GID>2184</GID>
<name>IN_1</name></connection>
<connection>
<GID>2187</GID>
<name>IN_1</name></connection>
<connection>
<GID>2190</GID>
<name>IN_1</name></connection>
<connection>
<GID>2193</GID>
<name>IN_1</name></connection>
<connection>
<GID>2196</GID>
<name>IN_1</name></connection>
<connection>
<GID>2199</GID>
<name>IN_1</name></connection>
<connection>
<GID>2202</GID>
<name>IN_1</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>244,-180.5,245,-180.5</points>
<connection>
<GID>2304</GID>
<name>OUT_0</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>1655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-192.5,280.5,-52.5</points>
<connection>
<GID>2174</GID>
<name>N_in1</name></connection>
<connection>
<GID>2182</GID>
<name>N_in0</name></connection>
<intersection>-172.5 1</intersection>
<intersection>-155.5 3</intersection>
<intersection>-139.5 4</intersection>
<intersection>-124 5</intersection>
<intersection>-107.5 6</intersection>
<intersection>-90.5 7</intersection>
<intersection>-74.5 8</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280.5,-172.5,281.5,-172.5</points>
<connection>
<GID>2186</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-59,284,-59</points>
<connection>
<GID>2391</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280.5,-155.5,282,-155.5</points>
<connection>
<GID>2210</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>280.5,-139.5,282.5,-139.5</points>
<connection>
<GID>2234</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>280.5,-124,283,-124</points>
<connection>
<GID>2258</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>280.5,-107.5,282.5,-107.5</points>
<connection>
<GID>2316</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>280.5,-90.5,283,-90.5</points>
<connection>
<GID>2343</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>280.5,-74.5,283.5,-74.5</points>
<connection>
<GID>2367</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-192.5,312.5,-52.5</points>
<connection>
<GID>2189</GID>
<name>IN_0</name></connection>
<connection>
<GID>2175</GID>
<name>N_in1</name></connection>
<connection>
<GID>2183</GID>
<name>N_in0</name></connection>
<intersection>-155.5 9</intersection>
<intersection>-139.5 10</intersection>
<intersection>-124 7</intersection>
<intersection>-107.5 11</intersection>
<intersection>-90.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-59,315,-59</points>
<connection>
<GID>2394</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>312.5,-74.5,314.5,-74.5</points>
<connection>
<GID>2370</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>312.5,-90.5,314,-90.5</points>
<connection>
<GID>2346</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>312.5,-124,314,-124</points>
<connection>
<GID>2261</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>312.5,-155.5,313,-155.5</points>
<connection>
<GID>2213</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>312.5,-139.5,313.5,-139.5</points>
<connection>
<GID>2237</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>312.5,-107.5,313.5,-107.5</points>
<connection>
<GID>2322</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343.5,-191.5,343.5,-52.5</points>
<connection>
<GID>2192</GID>
<name>IN_0</name></connection>
<connection>
<GID>2176</GID>
<name>N_in1</name></connection>
<connection>
<GID>2277</GID>
<name>N_in0</name></connection>
<intersection>-155.5 38</intersection>
<intersection>-139.5 21</intersection>
<intersection>-124 7</intersection>
<intersection>-107.5 20</intersection>
<intersection>-90.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>343.5,-59,346,-59</points>
<connection>
<GID>2397</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343.5,-74.5,345.5,-74.5</points>
<connection>
<GID>2373</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>343.5,-90.5,345,-90.5</points>
<connection>
<GID>2349</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>343.5,-124,345,-124</points>
<connection>
<GID>2264</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>343.5,-107.5,344.5,-107.5</points>
<connection>
<GID>2325</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>343.5,-139.5,344.5,-139.5</points>
<connection>
<GID>2240</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>343.5,-155.5,344,-155.5</points>
<connection>
<GID>2216</GID>
<name>IN_0</name></connection>
<intersection>343.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374.5,-155.5,374.5,-53</points>
<connection>
<GID>2328</GID>
<name>IN_0</name></connection>
<connection>
<GID>2243</GID>
<name>IN_0</name></connection>
<connection>
<GID>2278</GID>
<name>N_in0</name></connection>
<intersection>-155.5 9</intersection>
<intersection>-124 7</intersection>
<intersection>-90.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-59,376,-59</points>
<connection>
<GID>2400</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>374.5,-74.5,375.5,-74.5</points>
<connection>
<GID>2376</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>374.5,-90.5,375,-90.5</points>
<connection>
<GID>2352</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>374.5,-124,375,-124</points>
<connection>
<GID>2267</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>373.5,-155.5,374.5,-155.5</points>
<connection>
<GID>2219</GID>
<name>IN_0</name></connection>
<intersection>373.5 10</intersection>
<intersection>374.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>373.5,-190.5,373.5,-155.5</points>
<connection>
<GID>2195</GID>
<name>IN_0</name></connection>
<connection>
<GID>2177</GID>
<name>N_in1</name></connection>
<intersection>-155.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>1659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404.5,-190,404.5,-52.5</points>
<connection>
<GID>2198</GID>
<name>IN_0</name></connection>
<connection>
<GID>2178</GID>
<name>N_in1</name></connection>
<connection>
<GID>2279</GID>
<name>N_in0</name></connection>
<intersection>-155.5 13</intersection>
<intersection>-139.5 11</intersection>
<intersection>-124 9</intersection>
<intersection>-107.5 7</intersection>
<intersection>-90.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>404.5,-59,407,-59</points>
<connection>
<GID>2403</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>404.5,-74.5,406.5,-74.5</points>
<connection>
<GID>2379</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>404.5,-90.5,406,-90.5</points>
<connection>
<GID>2355</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>404.5,-107.5,405.5,-107.5</points>
<connection>
<GID>2331</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>404.5,-124,406,-124</points>
<connection>
<GID>2270</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>404.5,-139.5,405.5,-139.5</points>
<connection>
<GID>2246</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>404.5,-155.5,405,-155.5</points>
<connection>
<GID>2222</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,-189,435.5,-52.5</points>
<connection>
<GID>2201</GID>
<name>IN_0</name></connection>
<connection>
<GID>2180</GID>
<name>N_in1</name></connection>
<connection>
<GID>2280</GID>
<name>N_in0</name></connection>
<intersection>-155.5 13</intersection>
<intersection>-139.5 11</intersection>
<intersection>-124 9</intersection>
<intersection>-107.5 7</intersection>
<intersection>-90.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435.5,-59,438,-59</points>
<connection>
<GID>2406</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>435.5,-74.5,437.5,-74.5</points>
<connection>
<GID>2382</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>435.5,-90.5,437,-90.5</points>
<connection>
<GID>2358</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>435.5,-107.5,436.5,-107.5</points>
<connection>
<GID>2334</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>435.5,-124,437,-124</points>
<connection>
<GID>2273</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>435.5,-139.5,436.5,-139.5</points>
<connection>
<GID>2249</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>435.5,-155.5,436,-155.5</points>
<connection>
<GID>2225</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466.5,-191,466.5,-53</points>
<connection>
<GID>2204</GID>
<name>IN_0</name></connection>
<connection>
<GID>2179</GID>
<name>N_in1</name></connection>
<connection>
<GID>2281</GID>
<name>N_in0</name></connection>
<intersection>-155.5 13</intersection>
<intersection>-139.5 10</intersection>
<intersection>-124 8</intersection>
<intersection>-107.5 6</intersection>
<intersection>-90.5 4</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>466.5,-59,469,-59</points>
<connection>
<GID>2409</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>466.5,-74.5,468.5,-74.5</points>
<connection>
<GID>2385</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>466.5,-90.5,468,-90.5</points>
<connection>
<GID>2361</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>466.5,-107.5,467.5,-107.5</points>
<connection>
<GID>2337</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>466.5,-124,468,-124</points>
<connection>
<GID>2276</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>466.5,-139.5,467.5,-139.5</points>
<connection>
<GID>2252</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>466.5,-155.5,467,-155.5</points>
<connection>
<GID>2228</GID>
<name>IN_0</name></connection>
<intersection>466.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-200.5,278.5,-45.5</points>
<connection>
<GID>2283</GID>
<name>N_in1</name></connection>
<connection>
<GID>2282</GID>
<name>N_in0</name></connection>
<intersection>-178.5 13</intersection>
<intersection>-161.5 12</intersection>
<intersection>-145.5 11</intersection>
<intersection>-130 10</intersection>
<intersection>-113.5 9</intersection>
<intersection>-96.5 8</intersection>
<intersection>-80.5 7</intersection>
<intersection>-65 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>275,-65,278.5,-65</points>
<intersection>275 23</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>274.5,-80.5,278.5,-80.5</points>
<intersection>274.5 22</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>274,-96.5,278.5,-96.5</points>
<intersection>274 21</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>273.5,-113.5,278.5,-113.5</points>
<intersection>273.5 20</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>274,-130,278.5,-130</points>
<intersection>274 17</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>273.5,-145.5,278.5,-145.5</points>
<intersection>273.5 16</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>273,-161.5,278.5,-161.5</points>
<intersection>273 15</intersection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>272.5,-178.5,278.5,-178.5</points>
<intersection>272.5 14</intersection>
<intersection>278.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>272.5,-179.5,272.5,-178.5</points>
<connection>
<GID>2171</GID>
<name>OUT_0</name></connection>
<intersection>-178.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>273,-162.5,273,-161.5</points>
<connection>
<GID>2206</GID>
<name>OUT_0</name></connection>
<intersection>-161.5 12</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>273.5,-146.5,273.5,-145.5</points>
<connection>
<GID>2230</GID>
<name>OUT_0</name></connection>
<intersection>-145.5 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>274,-131,274,-130</points>
<connection>
<GID>2254</GID>
<name>OUT_0</name></connection>
<intersection>-130 10</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>273.5,-114.5,273.5,-113.5</points>
<connection>
<GID>2307</GID>
<name>OUT_0</name></connection>
<intersection>-113.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>274,-97.5,274,-96.5</points>
<connection>
<GID>2339</GID>
<name>OUT_0</name></connection>
<intersection>-96.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>274.5,-81.5,274.5,-80.5</points>
<connection>
<GID>2363</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 7</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>275,-66,275,-65</points>
<connection>
<GID>2387</GID>
<name>OUT_0</name></connection>
<intersection>-65 6</intersection></vsegment></shape></wire>
<wire>
<ID>1663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-179.5,309.5,-45.5</points>
<connection>
<GID>2296</GID>
<name>N_in0</name></connection>
<intersection>-179.5 13</intersection>
<intersection>-162.5 12</intersection>
<intersection>-146.5 11</intersection>
<intersection>-131 10</intersection>
<intersection>-114.5 9</intersection>
<intersection>-97.5 8</intersection>
<intersection>-81.5 7</intersection>
<intersection>-66 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>306.5,-66,309.5,-66</points>
<connection>
<GID>2390</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>306,-81.5,309.5,-81.5</points>
<connection>
<GID>2366</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>305.5,-97.5,309.5,-97.5</points>
<connection>
<GID>2342</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>305,-114.5,309.5,-114.5</points>
<connection>
<GID>2314</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>305.5,-131,309.5,-131</points>
<connection>
<GID>2257</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>305,-146.5,309.5,-146.5</points>
<connection>
<GID>2233</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>304.5,-162.5,309.5,-162.5</points>
<connection>
<GID>2209</GID>
<name>OUT_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>304,-179.5,309.5,-179.5</points>
<connection>
<GID>2185</GID>
<name>OUT_0</name></connection>
<intersection>306 22</intersection>
<intersection>309.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>306,-198.5,306,-179.5</points>
<connection>
<GID>5777</GID>
<name>N_in1</name></connection>
<intersection>-179.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-199.5,341.5,-45.5</points>
<connection>
<GID>2284</GID>
<name>N_in1</name></connection>
<connection>
<GID>2295</GID>
<name>N_in0</name></connection>
<intersection>-179.5 13</intersection>
<intersection>-162.5 12</intersection>
<intersection>-146.5 11</intersection>
<intersection>-131 10</intersection>
<intersection>-114.5 9</intersection>
<intersection>-97.5 8</intersection>
<intersection>-81.5 7</intersection>
<intersection>-66 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>337,-66,341.5,-66</points>
<connection>
<GID>2393</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>336.5,-81.5,341.5,-81.5</points>
<connection>
<GID>2369</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>336,-97.5,341.5,-97.5</points>
<connection>
<GID>2345</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>335.5,-114.5,341.5,-114.5</points>
<connection>
<GID>2320</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>336,-131,341.5,-131</points>
<connection>
<GID>2260</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>335.5,-146.5,341.5,-146.5</points>
<connection>
<GID>2236</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>335,-162.5,341.5,-162.5</points>
<connection>
<GID>2212</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>334.5,-179.5,341.5,-179.5</points>
<connection>
<GID>2188</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-199,372,-45.5</points>
<connection>
<GID>2285</GID>
<name>N_in1</name></connection>
<connection>
<GID>2294</GID>
<name>N_in0</name></connection>
<intersection>-179.5 18</intersection>
<intersection>-162.5 17</intersection>
<intersection>-146.5 16</intersection>
<intersection>-131 15</intersection>
<intersection>-114.5 14</intersection>
<intersection>-97.5 13</intersection>
<intersection>-81.5 12</intersection>
<intersection>-66 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>368.5,-66,372,-66</points>
<connection>
<GID>2396</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>368,-81.5,372,-81.5</points>
<connection>
<GID>2372</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>367.5,-97.5,372,-97.5</points>
<connection>
<GID>2348</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>367,-114.5,372,-114.5</points>
<connection>
<GID>2324</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>367.5,-131,372,-131</points>
<connection>
<GID>2263</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>367,-146.5,372,-146.5</points>
<connection>
<GID>2239</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>366.5,-162.5,372,-162.5</points>
<connection>
<GID>2215</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>366,-179.5,372,-179.5</points>
<connection>
<GID>2191</GID>
<name>OUT_0</name></connection>
<intersection>372 0</intersection></hsegment></shape></wire>
<wire>
<ID>1666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-199,402.5,-45.5</points>
<connection>
<GID>2286</GID>
<name>N_in1</name></connection>
<connection>
<GID>2293</GID>
<name>N_in0</name></connection>
<intersection>-179.5 9</intersection>
<intersection>-162.5 10</intersection>
<intersection>-146.5 11</intersection>
<intersection>-131 12</intersection>
<intersection>-114.5 13</intersection>
<intersection>-97.5 14</intersection>
<intersection>-81.5 15</intersection>
<intersection>-66 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>395.5,-179.5,402.5,-179.5</points>
<connection>
<GID>2194</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>396,-162.5,402.5,-162.5</points>
<connection>
<GID>2218</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>396.5,-146.5,402.5,-146.5</points>
<connection>
<GID>2242</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>397,-131,402.5,-131</points>
<connection>
<GID>2266</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>396.5,-114.5,402.5,-114.5</points>
<connection>
<GID>2327</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>397,-97.5,402.5,-97.5</points>
<connection>
<GID>2351</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>397.5,-81.5,402.5,-81.5</points>
<connection>
<GID>2375</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>398,-66,402.5,-66</points>
<connection>
<GID>2399</GID>
<name>OUT_0</name></connection>
<intersection>402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,-199,433.5,-45.5</points>
<connection>
<GID>2287</GID>
<name>N_in1</name></connection>
<connection>
<GID>2292</GID>
<name>N_in0</name></connection>
<intersection>-179.5 6</intersection>
<intersection>-162.5 7</intersection>
<intersection>-146.5 8</intersection>
<intersection>-131 9</intersection>
<intersection>-114.5 10</intersection>
<intersection>-97.5 11</intersection>
<intersection>-81.5 12</intersection>
<intersection>-66 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>427,-179.5,433.5,-179.5</points>
<connection>
<GID>2197</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>427.5,-162.5,433.5,-162.5</points>
<connection>
<GID>2221</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>428,-146.5,433.5,-146.5</points>
<connection>
<GID>2245</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>428.5,-131,433.5,-131</points>
<connection>
<GID>2269</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>428,-114.5,433.5,-114.5</points>
<connection>
<GID>2330</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>428.5,-97.5,433.5,-97.5</points>
<connection>
<GID>2354</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>429,-81.5,433.5,-81.5</points>
<connection>
<GID>2378</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>429.5,-66,433.5,-66</points>
<connection>
<GID>2402</GID>
<name>OUT_0</name></connection>
<intersection>433.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,-199.5,464.5,-44.5</points>
<connection>
<GID>2288</GID>
<name>N_in1</name></connection>
<connection>
<GID>2291</GID>
<name>N_in0</name></connection>
<intersection>-179.5 6</intersection>
<intersection>-162.5 7</intersection>
<intersection>-146.5 8</intersection>
<intersection>-131 9</intersection>
<intersection>-114.5 10</intersection>
<intersection>-97.5 11</intersection>
<intersection>-81.5 12</intersection>
<intersection>-66 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>457.5,-179.5,464.5,-179.5</points>
<connection>
<GID>2200</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>458,-162.5,464.5,-162.5</points>
<connection>
<GID>2224</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>458.5,-146.5,464.5,-146.5</points>
<connection>
<GID>2248</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>459,-131,464.5,-131</points>
<connection>
<GID>2272</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>458.5,-114.5,464.5,-114.5</points>
<connection>
<GID>2333</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>459,-97.5,464.5,-97.5</points>
<connection>
<GID>2357</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>459.5,-81.5,464.5,-81.5</points>
<connection>
<GID>2381</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>460,-66,464.5,-66</points>
<connection>
<GID>2405</GID>
<name>OUT_0</name></connection>
<intersection>464.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495,-199,495,-44</points>
<connection>
<GID>2289</GID>
<name>N_in1</name></connection>
<connection>
<GID>2290</GID>
<name>N_in0</name></connection>
<intersection>-179.5 3</intersection>
<intersection>-162.5 4</intersection>
<intersection>-146.5 5</intersection>
<intersection>-131 6</intersection>
<intersection>-114.5 7</intersection>
<intersection>-97.5 8</intersection>
<intersection>-81.5 9</intersection>
<intersection>-66 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>489,-179.5,495,-179.5</points>
<connection>
<GID>2203</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>489.5,-162.5,495,-162.5</points>
<connection>
<GID>2227</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>490,-146.5,495,-146.5</points>
<connection>
<GID>2251</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>490.5,-131,495,-131</points>
<connection>
<GID>2275</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>490,-114.5,495,-114.5</points>
<connection>
<GID>2336</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>490.5,-97.5,495,-97.5</points>
<connection>
<GID>2360</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>491,-81.5,495,-81.5</points>
<connection>
<GID>2384</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>491.5,-66,495,-66</points>
<connection>
<GID>2408</GID>
<name>OUT_0</name></connection>
<intersection>495 0</intersection></hsegment></shape></wire>
<wire>
<ID>1670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-113.5,203.5,-64.5</points>
<intersection>-113.5 2</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-64.5,242.5,-64.5</points>
<connection>
<GID>2309</GID>
<name>ENABLE_0</name></connection>
<intersection>203.5 0</intersection>
<intersection>228.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-113.5,203.5,-113.5</points>
<connection>
<GID>2297</GID>
<name>OUT_7</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228.5,-64.5,228.5,-61</points>
<intersection>-64.5 1</intersection>
<intersection>-61 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-61,233,-61</points>
<connection>
<GID>2310</GID>
<name>IN_0</name></connection>
<intersection>228.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-114.5,205.5,-80</points>
<intersection>-114.5 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-80,242.5,-80</points>
<intersection>205.5 0</intersection>
<intersection>228.5 4</intersection>
<intersection>242.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-114.5,205.5,-114.5</points>
<connection>
<GID>2297</GID>
<name>OUT_6</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,-80.5,242.5,-80</points>
<connection>
<GID>2311</GID>
<name>ENABLE_0</name></connection>
<intersection>-80 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>228.5,-80,228.5,-76.5</points>
<intersection>-80 1</intersection>
<intersection>-76.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-76.5,232.5,-76.5</points>
<connection>
<GID>2313</GID>
<name>IN_0</name></connection>
<intersection>228.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-115.5,207.5,-92.5</points>
<intersection>-115.5 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-92.5,232.5,-92.5</points>
<connection>
<GID>2317</GID>
<name>IN_0</name></connection>
<intersection>207.5 0</intersection>
<intersection>228.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-115.5,207.5,-115.5</points>
<connection>
<GID>2297</GID>
<name>OUT_5</name></connection>
<intersection>207.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>228.5,-96.5,228.5,-92.5</points>
<intersection>-96.5 4</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>228.5,-96.5,242.5,-96.5</points>
<connection>
<GID>2315</GID>
<name>ENABLE_0</name></connection>
<intersection>228.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209.5,-116.5,209.5,-109.5</points>
<intersection>-116.5 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-109.5,232.5,-109.5</points>
<connection>
<GID>2321</GID>
<name>IN_0</name></connection>
<intersection>209.5 0</intersection>
<intersection>228.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-116.5,209.5,-116.5</points>
<connection>
<GID>2297</GID>
<name>OUT_4</name></connection>
<intersection>209.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>228.5,-113.5,228.5,-109.5</points>
<intersection>-113.5 4</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>228.5,-113.5,242.5,-113.5</points>
<connection>
<GID>2319</GID>
<name>ENABLE_0</name></connection>
<intersection>228.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209.5,-129.5,209.5,-117.5</points>
<intersection>-129.5 1</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-129.5,241.5,-129.5</points>
<connection>
<GID>2298</GID>
<name>ENABLE_0</name></connection>
<intersection>209.5 0</intersection>
<intersection>228.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-117.5,209.5,-117.5</points>
<connection>
<GID>2297</GID>
<name>OUT_3</name></connection>
<intersection>209.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228.5,-129.5,228.5,-126</points>
<intersection>-129.5 1</intersection>
<intersection>-126 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-126,232.5,-126</points>
<connection>
<GID>2299</GID>
<name>IN_0</name></connection>
<intersection>228.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-145.5,207.5,-118.5</points>
<intersection>-145.5 1</intersection>
<intersection>-118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-145.5,241.5,-145.5</points>
<connection>
<GID>2300</GID>
<name>ENABLE_0</name></connection>
<intersection>207.5 0</intersection>
<intersection>228.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-118.5,207.5,-118.5</points>
<connection>
<GID>2297</GID>
<name>OUT_2</name></connection>
<intersection>207.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228.5,-145.5,228.5,-141.5</points>
<intersection>-145.5 1</intersection>
<intersection>-141.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-141.5,232.5,-141.5</points>
<connection>
<GID>2301</GID>
<name>IN_0</name></connection>
<intersection>228.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-161,205.5,-119.5</points>
<intersection>-161 1</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-161,241.5,-161</points>
<intersection>205.5 0</intersection>
<intersection>228.5 4</intersection>
<intersection>241.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-119.5,205.5,-119.5</points>
<connection>
<GID>2297</GID>
<name>OUT_1</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241.5,-161.5,241.5,-161</points>
<connection>
<GID>2302</GID>
<name>ENABLE_0</name></connection>
<intersection>-161 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>228.5,-161,228.5,-157.5</points>
<intersection>-161 1</intersection>
<intersection>-157.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-157.5,232.5,-157.5</points>
<connection>
<GID>2303</GID>
<name>IN_0</name></connection>
<intersection>228.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-178.5,203.5,-120.5</points>
<intersection>-178.5 1</intersection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-178.5,241.5,-178.5</points>
<connection>
<GID>2304</GID>
<name>ENABLE_0</name></connection>
<intersection>203.5 0</intersection>
<intersection>228.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-120.5,203.5,-120.5</points>
<connection>
<GID>2297</GID>
<name>OUT_0</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228.5,-178.5,228.5,-174.5</points>
<intersection>-178.5 1</intersection>
<intersection>-174.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-174.5,232.5,-174.5</points>
<connection>
<GID>2305</GID>
<name>IN_0</name></connection>
<intersection>228.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1678</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>269.5,-117,271.5,-117</points>
<connection>
<GID>2306</GID>
<name>OUT</name></connection>
<connection>
<GID>2307</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,-120.5,273.5,-120</points>
<connection>
<GID>2307</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-120.5,273.5,-120.5</points>
<intersection>259.5 2</intersection>
<intersection>273.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>259.5,-120.5,259.5,-107.5</points>
<intersection>-120.5 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,-116,263.5,-116</points>
<connection>
<GID>2306</GID>
<name>IN_0</name></connection>
<intersection>259.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>257.5,-107.5,259.5,-107.5</points>
<connection>
<GID>2308</GID>
<name>OUT_0</name></connection>
<intersection>259.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1680</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301,-117,303,-117</points>
<connection>
<GID>2312</GID>
<name>OUT</name></connection>
<connection>
<GID>2314</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1681</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291,-120,305,-120</points>
<connection>
<GID>2314</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291,-120,291,-107.5</points>
<intersection>-120 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291,-116,295,-116</points>
<connection>
<GID>2312</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>288.5,-107.5,291,-107.5</points>
<connection>
<GID>2316</GID>
<name>OUT_0</name></connection>
<intersection>291 2</intersection></hsegment></shape></wire>
<wire>
<ID>1682</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>331.5,-117,333.5,-117</points>
<connection>
<GID>2318</GID>
<name>OUT</name></connection>
<connection>
<GID>2320</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-120.5,335.5,-120</points>
<connection>
<GID>2320</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-120.5,335.5,-120.5</points>
<intersection>321.5 2</intersection>
<intersection>335.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321.5,-120.5,321.5,-107.5</points>
<intersection>-120.5 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321.5,-116,325.5,-116</points>
<connection>
<GID>2318</GID>
<name>IN_0</name></connection>
<intersection>321.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>319.5,-107.5,321.5,-107.5</points>
<connection>
<GID>2322</GID>
<name>OUT_0</name></connection>
<intersection>321.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1684</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363,-117,365,-117</points>
<connection>
<GID>2323</GID>
<name>OUT</name></connection>
<connection>
<GID>2324</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1685</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353,-120,367,-120</points>
<connection>
<GID>2324</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353,-120,353,-107.5</points>
<intersection>-120 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353,-116,357,-116</points>
<connection>
<GID>2323</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>350.5,-107.5,353,-107.5</points>
<connection>
<GID>2325</GID>
<name>OUT_0</name></connection>
<intersection>353 2</intersection></hsegment></shape></wire>
<wire>
<ID>1686</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>392.5,-117,394.5,-117</points>
<connection>
<GID>2326</GID>
<name>OUT</name></connection>
<connection>
<GID>2327</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-120.5,396.5,-120</points>
<connection>
<GID>2327</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382.5,-120.5,396.5,-120.5</points>
<intersection>382.5 2</intersection>
<intersection>396.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>382.5,-120.5,382.5,-107.5</points>
<intersection>-120.5 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>382.5,-116,386.5,-116</points>
<connection>
<GID>2326</GID>
<name>IN_0</name></connection>
<intersection>382.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380.5,-107.5,382.5,-107.5</points>
<connection>
<GID>2328</GID>
<name>OUT_0</name></connection>
<intersection>382.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1688</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424,-117,426,-117</points>
<connection>
<GID>2329</GID>
<name>OUT</name></connection>
<connection>
<GID>2330</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1689</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414,-120,428,-120</points>
<connection>
<GID>2330</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414,-120,414,-107.5</points>
<intersection>-120 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414,-116,418,-116</points>
<connection>
<GID>2329</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411.5,-107.5,414,-107.5</points>
<connection>
<GID>2331</GID>
<name>OUT_0</name></connection>
<intersection>414 2</intersection></hsegment></shape></wire>
<wire>
<ID>1690</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>454.5,-117,456.5,-117</points>
<connection>
<GID>2332</GID>
<name>OUT</name></connection>
<connection>
<GID>2333</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-120.5,458.5,-120</points>
<connection>
<GID>2333</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,-120.5,458.5,-120.5</points>
<intersection>444.5 2</intersection>
<intersection>458.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>444.5,-120.5,444.5,-107.5</points>
<intersection>-120.5 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>444.5,-116,448.5,-116</points>
<connection>
<GID>2332</GID>
<name>IN_0</name></connection>
<intersection>444.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>442.5,-107.5,444.5,-107.5</points>
<connection>
<GID>2334</GID>
<name>OUT_0</name></connection>
<intersection>444.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1692</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486,-117,488,-117</points>
<connection>
<GID>2335</GID>
<name>OUT</name></connection>
<connection>
<GID>2336</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1693</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476,-120,490,-120</points>
<connection>
<GID>2336</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476,-120,476,-107.5</points>
<intersection>-120 1</intersection>
<intersection>-116 4</intersection>
<intersection>-107.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476,-116,480,-116</points>
<connection>
<GID>2335</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>473.5,-107.5,476,-107.5</points>
<connection>
<GID>2337</GID>
<name>OUT_0</name></connection>
<intersection>476 2</intersection></hsegment></shape></wire>
<wire>
<ID>1694</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270,-100,272,-100</points>
<connection>
<GID>2338</GID>
<name>OUT</name></connection>
<connection>
<GID>2339</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-103.5,274,-103</points>
<connection>
<GID>2339</GID>
<name>IN_0</name></connection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-103.5,274,-103.5</points>
<intersection>260 2</intersection>
<intersection>274 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260,-103.5,260,-90.5</points>
<intersection>-103.5 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260,-99,264,-99</points>
<connection>
<GID>2338</GID>
<name>IN_0</name></connection>
<intersection>260 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258,-90.5,260,-90.5</points>
<connection>
<GID>2340</GID>
<name>OUT_0</name></connection>
<intersection>260 2</intersection></hsegment></shape></wire>
<wire>
<ID>1696</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,-100,303.5,-100</points>
<connection>
<GID>2341</GID>
<name>OUT</name></connection>
<connection>
<GID>2342</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,-103,305.5,-103</points>
<connection>
<GID>2342</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291.5,-103,291.5,-90.5</points>
<intersection>-103 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291.5,-99,295.5,-99</points>
<connection>
<GID>2341</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289,-90.5,291.5,-90.5</points>
<connection>
<GID>2343</GID>
<name>OUT_0</name></connection>
<intersection>291.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1698</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332,-100,334,-100</points>
<connection>
<GID>2344</GID>
<name>OUT</name></connection>
<connection>
<GID>2345</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,-103.5,336,-103</points>
<connection>
<GID>2345</GID>
<name>IN_0</name></connection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-103.5,336,-103.5</points>
<intersection>322 2</intersection>
<intersection>336 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322,-103.5,322,-90.5</points>
<intersection>-103.5 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322,-99,326,-99</points>
<connection>
<GID>2344</GID>
<name>IN_0</name></connection>
<intersection>322 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320,-90.5,322,-90.5</points>
<connection>
<GID>2346</GID>
<name>OUT_0</name></connection>
<intersection>322 2</intersection></hsegment></shape></wire>
<wire>
<ID>1700</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363.5,-100,365.5,-100</points>
<connection>
<GID>2347</GID>
<name>OUT</name></connection>
<connection>
<GID>2348</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1701</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353.5,-103,367.5,-103</points>
<connection>
<GID>2348</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353.5,-103,353.5,-90.5</points>
<intersection>-103 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353.5,-99,357.5,-99</points>
<connection>
<GID>2347</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351,-90.5,353.5,-90.5</points>
<connection>
<GID>2349</GID>
<name>OUT_0</name></connection>
<intersection>353.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1702</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393,-100,395,-100</points>
<connection>
<GID>2350</GID>
<name>OUT</name></connection>
<connection>
<GID>2351</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,-103.5,397,-103</points>
<connection>
<GID>2351</GID>
<name>IN_0</name></connection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383,-103.5,397,-103.5</points>
<intersection>383 2</intersection>
<intersection>397 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,-103.5,383,-90.5</points>
<intersection>-103.5 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383,-99,387,-99</points>
<connection>
<GID>2350</GID>
<name>IN_0</name></connection>
<intersection>383 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381,-90.5,383,-90.5</points>
<connection>
<GID>2352</GID>
<name>OUT_0</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>1704</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424.5,-100,426.5,-100</points>
<connection>
<GID>2353</GID>
<name>OUT</name></connection>
<connection>
<GID>2354</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414.5,-103,428.5,-103</points>
<connection>
<GID>2354</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414.5,-103,414.5,-90.5</points>
<intersection>-103 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414.5,-99,418.5,-99</points>
<connection>
<GID>2353</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412,-90.5,414.5,-90.5</points>
<connection>
<GID>2355</GID>
<name>OUT_0</name></connection>
<intersection>414.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1706</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455,-100,457,-100</points>
<connection>
<GID>2356</GID>
<name>OUT</name></connection>
<connection>
<GID>2357</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-103.5,459,-103</points>
<connection>
<GID>2357</GID>
<name>IN_0</name></connection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,-103.5,459,-103.5</points>
<intersection>445 2</intersection>
<intersection>459 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445,-103.5,445,-90.5</points>
<intersection>-103.5 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445,-99,449,-99</points>
<connection>
<GID>2356</GID>
<name>IN_0</name></connection>
<intersection>445 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443,-90.5,445,-90.5</points>
<connection>
<GID>2358</GID>
<name>OUT_0</name></connection>
<intersection>445 2</intersection></hsegment></shape></wire>
<wire>
<ID>1708</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486.5,-100,488.5,-100</points>
<connection>
<GID>2359</GID>
<name>OUT</name></connection>
<connection>
<GID>2360</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1709</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476.5,-103,490.5,-103</points>
<connection>
<GID>2360</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476.5,-103,476.5,-90.5</points>
<intersection>-103 1</intersection>
<intersection>-99 4</intersection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476.5,-99,480.5,-99</points>
<connection>
<GID>2359</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474,-90.5,476.5,-90.5</points>
<connection>
<GID>2361</GID>
<name>OUT_0</name></connection>
<intersection>476.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1710</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270.5,-84,272.5,-84</points>
<connection>
<GID>2362</GID>
<name>OUT</name></connection>
<connection>
<GID>2363</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-87.5,274.5,-87</points>
<connection>
<GID>2363</GID>
<name>IN_0</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-87.5,274.5,-87.5</points>
<intersection>260.5 2</intersection>
<intersection>274.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260.5,-87.5,260.5,-74.5</points>
<intersection>-87.5 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,-83,264.5,-83</points>
<connection>
<GID>2362</GID>
<name>IN_0</name></connection>
<intersection>260.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258.5,-74.5,260.5,-74.5</points>
<connection>
<GID>2364</GID>
<name>OUT_0</name></connection>
<intersection>260.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1712</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302,-84,304,-84</points>
<connection>
<GID>2365</GID>
<name>OUT</name></connection>
<connection>
<GID>2366</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-87,306,-87</points>
<connection>
<GID>2366</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292,-87,292,-74.5</points>
<intersection>-87 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292,-83,296,-83</points>
<connection>
<GID>2365</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289.5,-74.5,292,-74.5</points>
<connection>
<GID>2367</GID>
<name>OUT_0</name></connection>
<intersection>292 2</intersection></hsegment></shape></wire>
<wire>
<ID>1714</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332.5,-84,334.5,-84</points>
<connection>
<GID>2368</GID>
<name>OUT</name></connection>
<connection>
<GID>2369</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,-87.5,336.5,-87</points>
<connection>
<GID>2369</GID>
<name>IN_0</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,-87.5,336.5,-87.5</points>
<intersection>322.5 2</intersection>
<intersection>336.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322.5,-87.5,322.5,-74.5</points>
<intersection>-87.5 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322.5,-83,326.5,-83</points>
<connection>
<GID>2368</GID>
<name>IN_0</name></connection>
<intersection>322.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320.5,-74.5,322.5,-74.5</points>
<connection>
<GID>2370</GID>
<name>OUT_0</name></connection>
<intersection>322.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1716</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364,-84,366,-84</points>
<connection>
<GID>2371</GID>
<name>OUT</name></connection>
<connection>
<GID>2372</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1717</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354,-87,368,-87</points>
<connection>
<GID>2372</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354,-87,354,-74.5</points>
<intersection>-87 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354,-83,358,-83</points>
<connection>
<GID>2371</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351.5,-74.5,354,-74.5</points>
<connection>
<GID>2373</GID>
<name>OUT_0</name></connection>
<intersection>354 2</intersection></hsegment></shape></wire>
<wire>
<ID>1718</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393.5,-84,395.5,-84</points>
<connection>
<GID>2374</GID>
<name>OUT</name></connection>
<connection>
<GID>2375</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,-87.5,397.5,-87</points>
<connection>
<GID>2375</GID>
<name>IN_0</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,-87.5,397.5,-87.5</points>
<intersection>383.5 2</intersection>
<intersection>397.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,-87.5,383.5,-74.5</points>
<intersection>-87.5 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383.5,-83,387.5,-83</points>
<connection>
<GID>2374</GID>
<name>IN_0</name></connection>
<intersection>383.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381.5,-74.5,383.5,-74.5</points>
<connection>
<GID>2376</GID>
<name>OUT_0</name></connection>
<intersection>383.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1720</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425,-84,427,-84</points>
<connection>
<GID>2377</GID>
<name>OUT</name></connection>
<connection>
<GID>2378</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415,-87,429,-87</points>
<connection>
<GID>2378</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415,-87,415,-74.5</points>
<intersection>-87 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415,-83,419,-83</points>
<connection>
<GID>2377</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412.5,-74.5,415,-74.5</points>
<connection>
<GID>2379</GID>
<name>OUT_0</name></connection>
<intersection>415 2</intersection></hsegment></shape></wire>
<wire>
<ID>1722</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455.5,-84,457.5,-84</points>
<connection>
<GID>2380</GID>
<name>OUT</name></connection>
<connection>
<GID>2381</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-87.5,459.5,-87</points>
<connection>
<GID>2381</GID>
<name>IN_0</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,-87.5,459.5,-87.5</points>
<intersection>445.5 2</intersection>
<intersection>459.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445.5,-87.5,445.5,-74.5</points>
<intersection>-87.5 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445.5,-83,449.5,-83</points>
<connection>
<GID>2380</GID>
<name>IN_0</name></connection>
<intersection>445.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443.5,-74.5,445.5,-74.5</points>
<connection>
<GID>2382</GID>
<name>OUT_0</name></connection>
<intersection>445.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1724</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487,-84,489,-84</points>
<connection>
<GID>2383</GID>
<name>OUT</name></connection>
<connection>
<GID>2384</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,-87,491,-87</points>
<connection>
<GID>2384</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477,-87,477,-74.5</points>
<intersection>-87 1</intersection>
<intersection>-83 4</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477,-83,481,-83</points>
<connection>
<GID>2383</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474.5,-74.5,477,-74.5</points>
<connection>
<GID>2385</GID>
<name>OUT_0</name></connection>
<intersection>477 2</intersection></hsegment></shape></wire>
<wire>
<ID>1726</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271,-68.5,273,-68.5</points>
<connection>
<GID>2386</GID>
<name>OUT</name></connection>
<connection>
<GID>2387</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-72,275,-71.5</points>
<connection>
<GID>2387</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-72,275,-72</points>
<intersection>261 2</intersection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261,-72,261,-59</points>
<intersection>-72 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,-67.5,265,-67.5</points>
<connection>
<GID>2386</GID>
<name>IN_0</name></connection>
<intersection>261 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259,-59,261,-59</points>
<connection>
<GID>2388</GID>
<name>OUT_0</name></connection>
<intersection>261 2</intersection></hsegment></shape></wire>
<wire>
<ID>1728</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302.5,-68.5,304.5,-68.5</points>
<connection>
<GID>2389</GID>
<name>OUT</name></connection>
<connection>
<GID>2390</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1729</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-71.5,306.5,-71.5</points>
<connection>
<GID>2390</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292.5,-71.5,292.5,-59</points>
<intersection>-71.5 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-67.5,296.5,-67.5</points>
<connection>
<GID>2389</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290,-59,292.5,-59</points>
<connection>
<GID>2391</GID>
<name>OUT_0</name></connection>
<intersection>292.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1730</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333,-68.5,335,-68.5</points>
<connection>
<GID>2392</GID>
<name>OUT</name></connection>
<connection>
<GID>2393</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-72,337,-71.5</points>
<connection>
<GID>2393</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,-72,337,-72</points>
<intersection>323 2</intersection>
<intersection>337 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323,-72,323,-59</points>
<intersection>-72 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323,-67.5,327,-67.5</points>
<connection>
<GID>2392</GID>
<name>IN_0</name></connection>
<intersection>323 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321,-59,323,-59</points>
<connection>
<GID>2394</GID>
<name>OUT_0</name></connection>
<intersection>323 2</intersection></hsegment></shape></wire>
<wire>
<ID>1732</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364.5,-68.5,366.5,-68.5</points>
<connection>
<GID>2395</GID>
<name>OUT</name></connection>
<connection>
<GID>2396</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1733</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-71.5,368.5,-71.5</points>
<connection>
<GID>2396</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354.5,-71.5,354.5,-59</points>
<intersection>-71.5 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354.5,-67.5,358.5,-67.5</points>
<connection>
<GID>2395</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352,-59,354.5,-59</points>
<connection>
<GID>2397</GID>
<name>OUT_0</name></connection>
<intersection>354.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1734</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394,-68.5,396,-68.5</points>
<connection>
<GID>2398</GID>
<name>OUT</name></connection>
<connection>
<GID>2399</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,-72,398,-71.5</points>
<connection>
<GID>2399</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-72,398,-72</points>
<intersection>384 2</intersection>
<intersection>398 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384,-72,384,-59</points>
<intersection>-72 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384,-67.5,388,-67.5</points>
<connection>
<GID>2398</GID>
<name>IN_0</name></connection>
<intersection>384 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382,-59,384,-59</points>
<connection>
<GID>2400</GID>
<name>OUT_0</name></connection>
<intersection>384 2</intersection></hsegment></shape></wire>
<wire>
<ID>1736</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425.5,-68.5,427.5,-68.5</points>
<connection>
<GID>2401</GID>
<name>OUT</name></connection>
<connection>
<GID>2402</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1737</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415.5,-71.5,429.5,-71.5</points>
<connection>
<GID>2402</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415.5,-71.5,415.5,-59</points>
<intersection>-71.5 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415.5,-67.5,419.5,-67.5</points>
<connection>
<GID>2401</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413,-59,415.5,-59</points>
<connection>
<GID>2403</GID>
<name>OUT_0</name></connection>
<intersection>415.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1738</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456,-68.5,458,-68.5</points>
<connection>
<GID>2404</GID>
<name>OUT</name></connection>
<connection>
<GID>2405</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460,-72,460,-71.5</points>
<connection>
<GID>2405</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446,-72,460,-72</points>
<intersection>446 2</intersection>
<intersection>460 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446,-72,446,-59</points>
<intersection>-72 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446,-67.5,450,-67.5</points>
<connection>
<GID>2404</GID>
<name>IN_0</name></connection>
<intersection>446 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444,-59,446,-59</points>
<connection>
<GID>2406</GID>
<name>OUT_0</name></connection>
<intersection>446 2</intersection></hsegment></shape></wire>
<wire>
<ID>1740</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487.5,-68.5,489.5,-68.5</points>
<connection>
<GID>2407</GID>
<name>OUT</name></connection>
<connection>
<GID>2408</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-71.5,491.5,-71.5</points>
<connection>
<GID>2408</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477.5,-71.5,477.5,-59</points>
<intersection>-71.5 1</intersection>
<intersection>-67.5 4</intersection>
<intersection>-59 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477.5,-67.5,481.5,-67.5</points>
<connection>
<GID>2407</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475,-59,477.5,-59</points>
<connection>
<GID>2409</GID>
<name>OUT_0</name></connection>
<intersection>477.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-192,249.5,-52.5</points>
<connection>
<GID>2173</GID>
<name>N_in1</name></connection>
<connection>
<GID>2181</GID>
<name>N_in0</name></connection>
<intersection>-172.5 14</intersection>
<intersection>-155.5 12</intersection>
<intersection>-139.5 10</intersection>
<intersection>-124 8</intersection>
<intersection>-107.5 6</intersection>
<intersection>-90.5 4</intersection>
<intersection>-74.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,-59,253,-59</points>
<connection>
<GID>2388</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-74.5,252.5,-74.5</points>
<connection>
<GID>2364</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>249.5,-90.5,252,-90.5</points>
<connection>
<GID>2340</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>249.5,-107.5,251.5,-107.5</points>
<connection>
<GID>2308</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>249.5,-124,252,-124</points>
<connection>
<GID>2255</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>249.5,-139.5,251.5,-139.5</points>
<connection>
<GID>2231</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>249.5,-155.5,251,-155.5</points>
<connection>
<GID>2207</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>249.5,-172.5,250.5,-172.5</points>
<connection>
<GID>2172</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1743</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-69.5,481.5,-69.5</points>
<connection>
<GID>2386</GID>
<name>IN_1</name></connection>
<connection>
<GID>2389</GID>
<name>IN_1</name></connection>
<connection>
<GID>2392</GID>
<name>IN_1</name></connection>
<connection>
<GID>2395</GID>
<name>IN_1</name></connection>
<connection>
<GID>2398</GID>
<name>IN_1</name></connection>
<connection>
<GID>2401</GID>
<name>IN_1</name></connection>
<connection>
<GID>2404</GID>
<name>IN_1</name></connection>
<connection>
<GID>2407</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-69.5,245,-66.5</points>
<connection>
<GID>2309</GID>
<name>OUT_0</name></connection>
<intersection>-69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239,-62,469,-62</points>
<connection>
<GID>2310</GID>
<name>OUT</name></connection>
<connection>
<GID>2388</GID>
<name>clock</name></connection>
<connection>
<GID>2391</GID>
<name>clock</name></connection>
<connection>
<GID>2394</GID>
<name>clock</name></connection>
<connection>
<GID>2397</GID>
<name>clock</name></connection>
<connection>
<GID>2400</GID>
<name>clock</name></connection>
<connection>
<GID>2403</GID>
<name>clock</name></connection>
<connection>
<GID>2406</GID>
<name>clock</name></connection>
<connection>
<GID>2409</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3425</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>264.5,203,266.5,203</points>
<connection>
<GID>4810</GID>
<name>OUT</name></connection>
<connection>
<GID>4811</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,199.5,268.5,200</points>
<connection>
<GID>4811</GID>
<name>IN_0</name></connection>
<intersection>199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>254.5,199.5,268.5,199.5</points>
<intersection>254.5 2</intersection>
<intersection>268.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>254.5,199.5,254.5,212.5</points>
<intersection>199.5 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>254.5,204,258.5,204</points>
<connection>
<GID>4810</GID>
<name>IN_0</name></connection>
<intersection>254.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>252.5,212.5,254.5,212.5</points>
<connection>
<GID>4812</GID>
<name>OUT_0</name></connection>
<intersection>254.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,300,477,300</points>
<connection>
<GID>5002</GID>
<name>IN_1</name></connection>
<connection>
<GID>5005</GID>
<name>IN_1</name></connection>
<connection>
<GID>5008</GID>
<name>IN_1</name></connection>
<connection>
<GID>5011</GID>
<name>IN_1</name></connection>
<connection>
<GID>5014</GID>
<name>IN_1</name></connection>
<connection>
<GID>5017</GID>
<name>IN_1</name></connection>
<connection>
<GID>5020</GID>
<name>IN_1</name></connection>
<connection>
<GID>5023</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,300,241,302.5</points>
<connection>
<GID>4951</GID>
<name>OUT_0</name></connection>
<intersection>300 1</intersection></vsegment></shape></wire>
<wire>
<ID>3428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,307.5,464.5,307.5</points>
<connection>
<GID>4953</GID>
<name>OUT</name></connection>
<connection>
<GID>5004</GID>
<name>clock</name></connection>
<connection>
<GID>5007</GID>
<name>clock</name></connection>
<connection>
<GID>5010</GID>
<name>clock</name></connection>
<connection>
<GID>5013</GID>
<name>clock</name></connection>
<connection>
<GID>5016</GID>
<name>clock</name></connection>
<connection>
<GID>5019</GID>
<name>clock</name></connection>
<connection>
<GID>5022</GID>
<name>clock</name></connection>
<connection>
<GID>5025</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3429</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,284,476.5,284</points>
<connection>
<GID>4978</GID>
<name>IN_1</name></connection>
<connection>
<GID>4981</GID>
<name>IN_1</name></connection>
<connection>
<GID>4984</GID>
<name>IN_1</name></connection>
<connection>
<GID>4987</GID>
<name>IN_1</name></connection>
<connection>
<GID>4990</GID>
<name>IN_1</name></connection>
<connection>
<GID>4993</GID>
<name>IN_1</name></connection>
<connection>
<GID>4996</GID>
<name>IN_1</name></connection>
<connection>
<GID>4999</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,284,241,286.5</points>
<connection>
<GID>4955</GID>
<name>OUT_0</name></connection>
<intersection>284 1</intersection></vsegment></shape></wire>
<wire>
<ID>3430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,291.5,464,291.5</points>
<connection>
<GID>4957</GID>
<name>OUT</name></connection>
<connection>
<GID>4980</GID>
<name>clock</name></connection>
<connection>
<GID>4983</GID>
<name>clock</name></connection>
<connection>
<GID>4986</GID>
<name>clock</name></connection>
<connection>
<GID>4989</GID>
<name>clock</name></connection>
<connection>
<GID>4992</GID>
<name>clock</name></connection>
<connection>
<GID>4995</GID>
<name>clock</name></connection>
<connection>
<GID>4998</GID>
<name>clock</name></connection>
<connection>
<GID>5001</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3431</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,274.5,463.5,274.5</points>
<connection>
<GID>4977</GID>
<name>clock</name></connection>
<connection>
<GID>4974</GID>
<name>clock</name></connection>
<connection>
<GID>4971</GID>
<name>clock</name></connection>
<connection>
<GID>4968</GID>
<name>clock</name></connection>
<connection>
<GID>4965</GID>
<name>clock</name></connection>
<connection>
<GID>4962</GID>
<name>clock</name></connection>
<connection>
<GID>4961</GID>
<name>OUT</name></connection>
<connection>
<GID>4956</GID>
<name>clock</name></connection>
<connection>
<GID>4948</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3432</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,267,476,267</points>
<connection>
<GID>4946</GID>
<name>IN_1</name></connection>
<connection>
<GID>4952</GID>
<name>IN_1</name></connection>
<connection>
<GID>4958</GID>
<name>IN_1</name></connection>
<connection>
<GID>4963</GID>
<name>IN_1</name></connection>
<connection>
<GID>4966</GID>
<name>IN_1</name></connection>
<connection>
<GID>4969</GID>
<name>IN_1</name></connection>
<connection>
<GID>4972</GID>
<name>IN_1</name></connection>
<connection>
<GID>4975</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,267,241,269.5</points>
<connection>
<GID>4959</GID>
<name>OUT_0</name></connection>
<intersection>267 1</intersection></vsegment></shape></wire>
<wire>
<ID>3433</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,258,464,258</points>
<connection>
<GID>4939</GID>
<name>OUT</name></connection>
<connection>
<GID>4916</GID>
<name>clock</name></connection>
<connection>
<GID>4913</GID>
<name>clock</name></connection>
<connection>
<GID>4910</GID>
<name>clock</name></connection>
<connection>
<GID>4907</GID>
<name>clock</name></connection>
<connection>
<GID>4904</GID>
<name>clock</name></connection>
<connection>
<GID>4901</GID>
<name>clock</name></connection>
<connection>
<GID>4898</GID>
<name>clock</name></connection>
<connection>
<GID>4895</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,250.5,476.5,250.5</points>
<connection>
<GID>4893</GID>
<name>IN_1</name></connection>
<connection>
<GID>4896</GID>
<name>IN_1</name></connection>
<connection>
<GID>4899</GID>
<name>IN_1</name></connection>
<connection>
<GID>4902</GID>
<name>IN_1</name></connection>
<connection>
<GID>4905</GID>
<name>IN_1</name></connection>
<connection>
<GID>4908</GID>
<name>IN_1</name></connection>
<connection>
<GID>4911</GID>
<name>IN_1</name></connection>
<connection>
<GID>4914</GID>
<name>IN_1</name></connection>
<intersection>240 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240,250.5,240,253.5</points>
<connection>
<GID>4938</GID>
<name>OUT_0</name></connection>
<intersection>250.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,242.5,463.5,242.5</points>
<connection>
<GID>4941</GID>
<name>OUT</name></connection>
<connection>
<GID>4892</GID>
<name>clock</name></connection>
<connection>
<GID>4889</GID>
<name>clock</name></connection>
<connection>
<GID>4886</GID>
<name>clock</name></connection>
<connection>
<GID>4883</GID>
<name>clock</name></connection>
<connection>
<GID>4880</GID>
<name>clock</name></connection>
<connection>
<GID>4877</GID>
<name>clock</name></connection>
<connection>
<GID>4874</GID>
<name>clock</name></connection>
<connection>
<GID>4871</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,235,476,235</points>
<connection>
<GID>4869</GID>
<name>IN_1</name></connection>
<connection>
<GID>4872</GID>
<name>IN_1</name></connection>
<connection>
<GID>4875</GID>
<name>IN_1</name></connection>
<connection>
<GID>4878</GID>
<name>IN_1</name></connection>
<connection>
<GID>4881</GID>
<name>IN_1</name></connection>
<connection>
<GID>4884</GID>
<name>IN_1</name></connection>
<connection>
<GID>4887</GID>
<name>IN_1</name></connection>
<connection>
<GID>4890</GID>
<name>IN_1</name></connection>
<intersection>240 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240,235,240,237.5</points>
<connection>
<GID>4940</GID>
<name>OUT_0</name></connection>
<intersection>235 1</intersection></vsegment></shape></wire>
<wire>
<ID>3437</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>296,203,298,203</points>
<connection>
<GID>4824</GID>
<name>OUT</name></connection>
<connection>
<GID>4825</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286,200,300,200</points>
<connection>
<GID>4825</GID>
<name>IN_0</name></connection>
<intersection>286 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>286,200,286,212.5</points>
<intersection>200 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>286,204,290,204</points>
<connection>
<GID>4824</GID>
<name>IN_0</name></connection>
<intersection>286 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>283.5,212.5,286,212.5</points>
<connection>
<GID>4826</GID>
<name>OUT_0</name></connection>
<intersection>286 2</intersection></hsegment></shape></wire>
<wire>
<ID>3439</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>326.5,203,328.5,203</points>
<connection>
<GID>4827</GID>
<name>OUT</name></connection>
<connection>
<GID>4828</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,199.5,330.5,200</points>
<connection>
<GID>4828</GID>
<name>IN_0</name></connection>
<intersection>199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316.5,199.5,330.5,199.5</points>
<intersection>316.5 2</intersection>
<intersection>330.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>316.5,199.5,316.5,212.5</points>
<intersection>199.5 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>316.5,204,320.5,204</points>
<connection>
<GID>4827</GID>
<name>IN_0</name></connection>
<intersection>316.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>314.5,212.5,316.5,212.5</points>
<connection>
<GID>4829</GID>
<name>OUT_0</name></connection>
<intersection>316.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3441</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>358,203,360,203</points>
<connection>
<GID>4830</GID>
<name>OUT</name></connection>
<connection>
<GID>4831</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3442</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>348,200,362,200</points>
<connection>
<GID>4831</GID>
<name>IN_0</name></connection>
<intersection>348 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>348,200,348,212.5</points>
<intersection>200 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>348,204,352,204</points>
<connection>
<GID>4830</GID>
<name>IN_0</name></connection>
<intersection>348 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>345.5,212.5,348,212.5</points>
<connection>
<GID>4832</GID>
<name>OUT_0</name></connection>
<intersection>348 2</intersection></hsegment></shape></wire>
<wire>
<ID>3443</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>387.5,203,389.5,203</points>
<connection>
<GID>4833</GID>
<name>OUT</name></connection>
<connection>
<GID>4834</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>391.5,199.5,391.5,200</points>
<connection>
<GID>4834</GID>
<name>IN_0</name></connection>
<intersection>199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377.5,199.5,391.5,199.5</points>
<intersection>377.5 2</intersection>
<intersection>391.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>377.5,199.5,377.5,212.5</points>
<intersection>199.5 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>377.5,204,381.5,204</points>
<connection>
<GID>4833</GID>
<name>IN_0</name></connection>
<intersection>377.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>375.5,212.5,377.5,212.5</points>
<connection>
<GID>4835</GID>
<name>OUT_0</name></connection>
<intersection>377.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3445</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>419,203,421,203</points>
<connection>
<GID>4836</GID>
<name>OUT</name></connection>
<connection>
<GID>4837</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>409,200,423,200</points>
<connection>
<GID>4837</GID>
<name>IN_0</name></connection>
<intersection>409 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>409,200,409,212.5</points>
<intersection>200 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>409,204,413,204</points>
<connection>
<GID>4836</GID>
<name>IN_0</name></connection>
<intersection>409 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>406.5,212.5,409,212.5</points>
<connection>
<GID>4838</GID>
<name>OUT_0</name></connection>
<intersection>409 2</intersection></hsegment></shape></wire>
<wire>
<ID>3447</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>449.5,203,451.5,203</points>
<connection>
<GID>4839</GID>
<name>OUT</name></connection>
<connection>
<GID>4840</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453.5,199.5,453.5,200</points>
<connection>
<GID>4840</GID>
<name>IN_0</name></connection>
<intersection>199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>439.5,199.5,453.5,199.5</points>
<intersection>439.5 2</intersection>
<intersection>453.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>439.5,199.5,439.5,212.5</points>
<intersection>199.5 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>439.5,204,443.5,204</points>
<connection>
<GID>4839</GID>
<name>IN_0</name></connection>
<intersection>439.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>437.5,212.5,439.5,212.5</points>
<connection>
<GID>4841</GID>
<name>OUT_0</name></connection>
<intersection>439.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3449</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>481,203,483,203</points>
<connection>
<GID>4842</GID>
<name>OUT</name></connection>
<connection>
<GID>4843</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>471,200,485,200</points>
<connection>
<GID>4843</GID>
<name>IN_0</name></connection>
<intersection>471 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>471,200,471,212.5</points>
<intersection>200 1</intersection>
<intersection>204 4</intersection>
<intersection>212.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>471,204,475,204</points>
<connection>
<GID>4842</GID>
<name>IN_0</name></connection>
<intersection>471 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>468.5,212.5,471,212.5</points>
<connection>
<GID>4844</GID>
<name>OUT_0</name></connection>
<intersection>471 2</intersection></hsegment></shape></wire>
<wire>
<ID>3451</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>265,220,267,220</points>
<connection>
<GID>4845</GID>
<name>OUT</name></connection>
<connection>
<GID>4846</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,216.5,269,217</points>
<connection>
<GID>4846</GID>
<name>IN_0</name></connection>
<intersection>216.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,216.5,269,216.5</points>
<intersection>255 2</intersection>
<intersection>269 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>255,216.5,255,229.5</points>
<intersection>216.5 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>255,221,259,221</points>
<connection>
<GID>4845</GID>
<name>IN_0</name></connection>
<intersection>255 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>253,229.5,255,229.5</points>
<connection>
<GID>4847</GID>
<name>OUT_0</name></connection>
<intersection>255 2</intersection></hsegment></shape></wire>
<wire>
<ID>3453</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>296.5,220,298.5,220</points>
<connection>
<GID>4848</GID>
<name>OUT</name></connection>
<connection>
<GID>4849</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286.5,217,300.5,217</points>
<connection>
<GID>4849</GID>
<name>IN_0</name></connection>
<intersection>286.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>286.5,217,286.5,229.5</points>
<intersection>217 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>286.5,221,290.5,221</points>
<connection>
<GID>4848</GID>
<name>IN_0</name></connection>
<intersection>286.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>284,229.5,286.5,229.5</points>
<connection>
<GID>4850</GID>
<name>OUT_0</name></connection>
<intersection>286.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3455</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>327,220,329,220</points>
<connection>
<GID>4851</GID>
<name>OUT</name></connection>
<connection>
<GID>4852</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331,216.5,331,217</points>
<connection>
<GID>4852</GID>
<name>IN_0</name></connection>
<intersection>216.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,216.5,331,216.5</points>
<intersection>317 2</intersection>
<intersection>331 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>317,216.5,317,229.5</points>
<intersection>216.5 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>317,221,321,221</points>
<connection>
<GID>4851</GID>
<name>IN_0</name></connection>
<intersection>317 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>315,229.5,317,229.5</points>
<connection>
<GID>4853</GID>
<name>OUT_0</name></connection>
<intersection>317 2</intersection></hsegment></shape></wire>
<wire>
<ID>3457</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>358.5,220,360.5,220</points>
<connection>
<GID>4854</GID>
<name>OUT</name></connection>
<connection>
<GID>4855</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>348.5,217,362.5,217</points>
<connection>
<GID>4855</GID>
<name>IN_0</name></connection>
<intersection>348.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>348.5,217,348.5,229.5</points>
<intersection>217 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>348.5,221,352.5,221</points>
<connection>
<GID>4854</GID>
<name>IN_0</name></connection>
<intersection>348.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>346,229.5,348.5,229.5</points>
<connection>
<GID>4856</GID>
<name>OUT_0</name></connection>
<intersection>348.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3459</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>388,220,390,220</points>
<connection>
<GID>4857</GID>
<name>OUT</name></connection>
<connection>
<GID>4858</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392,216.5,392,217</points>
<connection>
<GID>4858</GID>
<name>IN_0</name></connection>
<intersection>216.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378,216.5,392,216.5</points>
<intersection>378 2</intersection>
<intersection>392 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>378,216.5,378,229.5</points>
<intersection>216.5 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>378,221,382,221</points>
<connection>
<GID>4857</GID>
<name>IN_0</name></connection>
<intersection>378 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>376,229.5,378,229.5</points>
<connection>
<GID>4859</GID>
<name>OUT_0</name></connection>
<intersection>378 2</intersection></hsegment></shape></wire>
<wire>
<ID>3461</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>419.5,220,421.5,220</points>
<connection>
<GID>4860</GID>
<name>OUT</name></connection>
<connection>
<GID>4861</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>409.5,217,423.5,217</points>
<connection>
<GID>4861</GID>
<name>IN_0</name></connection>
<intersection>409.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>409.5,217,409.5,229.5</points>
<intersection>217 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>409.5,221,413.5,221</points>
<connection>
<GID>4860</GID>
<name>IN_0</name></connection>
<intersection>409.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>407,229.5,409.5,229.5</points>
<connection>
<GID>4862</GID>
<name>OUT_0</name></connection>
<intersection>409.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3463</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>450,220,452,220</points>
<connection>
<GID>4863</GID>
<name>OUT</name></connection>
<connection>
<GID>4864</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,216.5,454,217</points>
<connection>
<GID>4864</GID>
<name>IN_0</name></connection>
<intersection>216.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>440,216.5,454,216.5</points>
<intersection>440 2</intersection>
<intersection>454 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>440,216.5,440,229.5</points>
<intersection>216.5 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>440,221,444,221</points>
<connection>
<GID>4863</GID>
<name>IN_0</name></connection>
<intersection>440 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>438,229.5,440,229.5</points>
<connection>
<GID>4865</GID>
<name>OUT_0</name></connection>
<intersection>440 2</intersection></hsegment></shape></wire>
<wire>
<ID>3465</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>481.5,220,483.5,220</points>
<connection>
<GID>4866</GID>
<name>OUT</name></connection>
<connection>
<GID>4867</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>471.5,217,485.5,217</points>
<connection>
<GID>4867</GID>
<name>IN_0</name></connection>
<intersection>471.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>471.5,217,471.5,229.5</points>
<intersection>217 1</intersection>
<intersection>221 4</intersection>
<intersection>229.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>471.5,221,475.5,221</points>
<connection>
<GID>4866</GID>
<name>IN_0</name></connection>
<intersection>471.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>469,229.5,471.5,229.5</points>
<connection>
<GID>4868</GID>
<name>OUT_0</name></connection>
<intersection>471.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3467</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>265.5,236,267.5,236</points>
<connection>
<GID>4869</GID>
<name>OUT</name></connection>
<connection>
<GID>4870</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,232.5,269.5,233</points>
<connection>
<GID>4870</GID>
<name>IN_0</name></connection>
<intersection>232.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,232.5,269.5,232.5</points>
<intersection>255.5 2</intersection>
<intersection>269.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>255.5,232.5,255.5,245.5</points>
<intersection>232.5 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>255.5,237,259.5,237</points>
<connection>
<GID>4869</GID>
<name>IN_0</name></connection>
<intersection>255.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>253.5,245.5,255.5,245.5</points>
<connection>
<GID>4871</GID>
<name>OUT_0</name></connection>
<intersection>255.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3469</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297,236,299,236</points>
<connection>
<GID>4872</GID>
<name>OUT</name></connection>
<connection>
<GID>4873</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,233,301,233</points>
<connection>
<GID>4873</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287,233,287,245.5</points>
<intersection>233 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287,237,291,237</points>
<connection>
<GID>4872</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>284.5,245.5,287,245.5</points>
<connection>
<GID>4874</GID>
<name>OUT_0</name></connection>
<intersection>287 2</intersection></hsegment></shape></wire>
<wire>
<ID>3471</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>327.5,236,329.5,236</points>
<connection>
<GID>4875</GID>
<name>OUT</name></connection>
<connection>
<GID>4876</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,232.5,331.5,233</points>
<connection>
<GID>4876</GID>
<name>IN_0</name></connection>
<intersection>232.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,232.5,331.5,232.5</points>
<intersection>317.5 2</intersection>
<intersection>331.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>317.5,232.5,317.5,245.5</points>
<intersection>232.5 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>317.5,237,321.5,237</points>
<connection>
<GID>4875</GID>
<name>IN_0</name></connection>
<intersection>317.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>315.5,245.5,317.5,245.5</points>
<connection>
<GID>4877</GID>
<name>OUT_0</name></connection>
<intersection>317.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3473</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359,236,361,236</points>
<connection>
<GID>4878</GID>
<name>OUT</name></connection>
<connection>
<GID>4879</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,233,363,233</points>
<connection>
<GID>4879</GID>
<name>IN_0</name></connection>
<intersection>349 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349,233,349,245.5</points>
<intersection>233 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349,237,353,237</points>
<connection>
<GID>4878</GID>
<name>IN_0</name></connection>
<intersection>349 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>346.5,245.5,349,245.5</points>
<connection>
<GID>4880</GID>
<name>OUT_0</name></connection>
<intersection>349 2</intersection></hsegment></shape></wire>
<wire>
<ID>3475</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>388.5,236,390.5,236</points>
<connection>
<GID>4881</GID>
<name>OUT</name></connection>
<connection>
<GID>4882</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392.5,232.5,392.5,233</points>
<connection>
<GID>4882</GID>
<name>IN_0</name></connection>
<intersection>232.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378.5,232.5,392.5,232.5</points>
<intersection>378.5 2</intersection>
<intersection>392.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>378.5,232.5,378.5,245.5</points>
<intersection>232.5 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>378.5,237,382.5,237</points>
<connection>
<GID>4881</GID>
<name>IN_0</name></connection>
<intersection>378.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>376.5,245.5,378.5,245.5</points>
<connection>
<GID>4883</GID>
<name>OUT_0</name></connection>
<intersection>378.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3477</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420,236,422,236</points>
<connection>
<GID>4884</GID>
<name>OUT</name></connection>
<connection>
<GID>4885</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410,233,424,233</points>
<connection>
<GID>4885</GID>
<name>IN_0</name></connection>
<intersection>410 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410,233,410,245.5</points>
<intersection>233 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410,237,414,237</points>
<connection>
<GID>4884</GID>
<name>IN_0</name></connection>
<intersection>410 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>407.5,245.5,410,245.5</points>
<connection>
<GID>4886</GID>
<name>OUT_0</name></connection>
<intersection>410 2</intersection></hsegment></shape></wire>
<wire>
<ID>3479</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>450.5,236,452.5,236</points>
<connection>
<GID>4887</GID>
<name>OUT</name></connection>
<connection>
<GID>4888</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,232.5,454.5,233</points>
<connection>
<GID>4888</GID>
<name>IN_0</name></connection>
<intersection>232.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>440.5,232.5,454.5,232.5</points>
<intersection>440.5 2</intersection>
<intersection>454.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>440.5,232.5,440.5,245.5</points>
<intersection>232.5 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>440.5,237,444.5,237</points>
<connection>
<GID>4887</GID>
<name>IN_0</name></connection>
<intersection>440.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>438.5,245.5,440.5,245.5</points>
<connection>
<GID>4889</GID>
<name>OUT_0</name></connection>
<intersection>440.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3481</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482,236,484,236</points>
<connection>
<GID>4890</GID>
<name>OUT</name></connection>
<connection>
<GID>4891</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3482</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472,233,486,233</points>
<connection>
<GID>4891</GID>
<name>IN_0</name></connection>
<intersection>472 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472,233,472,245.5</points>
<intersection>233 1</intersection>
<intersection>237 4</intersection>
<intersection>245.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472,237,476,237</points>
<connection>
<GID>4890</GID>
<name>IN_0</name></connection>
<intersection>472 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>469.5,245.5,472,245.5</points>
<connection>
<GID>4892</GID>
<name>OUT_0</name></connection>
<intersection>472 2</intersection></hsegment></shape></wire>
<wire>
<ID>3483</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266,251.5,268,251.5</points>
<connection>
<GID>4893</GID>
<name>OUT</name></connection>
<connection>
<GID>4894</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,248,270,248.5</points>
<connection>
<GID>4894</GID>
<name>IN_0</name></connection>
<intersection>248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,248,270,248</points>
<intersection>256 2</intersection>
<intersection>270 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256,248,256,261</points>
<intersection>248 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256,252.5,260,252.5</points>
<connection>
<GID>4893</GID>
<name>IN_0</name></connection>
<intersection>256 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254,261,256,261</points>
<connection>
<GID>4895</GID>
<name>OUT_0</name></connection>
<intersection>256 2</intersection></hsegment></shape></wire>
<wire>
<ID>3485</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297.5,251.5,299.5,251.5</points>
<connection>
<GID>4896</GID>
<name>OUT</name></connection>
<connection>
<GID>4897</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287.5,248.5,301.5,248.5</points>
<connection>
<GID>4897</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287.5,248.5,287.5,261</points>
<intersection>248.5 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,252.5,291.5,252.5</points>
<connection>
<GID>4896</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285,261,287.5,261</points>
<connection>
<GID>4898</GID>
<name>OUT_0</name></connection>
<intersection>287.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3487</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328,251.5,330,251.5</points>
<connection>
<GID>4899</GID>
<name>OUT</name></connection>
<connection>
<GID>4900</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,248,332,248.5</points>
<connection>
<GID>4900</GID>
<name>IN_0</name></connection>
<intersection>248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,248,332,248</points>
<intersection>318 2</intersection>
<intersection>332 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318,248,318,261</points>
<intersection>248 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318,252.5,322,252.5</points>
<connection>
<GID>4899</GID>
<name>IN_0</name></connection>
<intersection>318 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316,261,318,261</points>
<connection>
<GID>4901</GID>
<name>OUT_0</name></connection>
<intersection>318 2</intersection></hsegment></shape></wire>
<wire>
<ID>3489</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359.5,251.5,361.5,251.5</points>
<connection>
<GID>4902</GID>
<name>OUT</name></connection>
<connection>
<GID>4903</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3490</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349.5,248.5,363.5,248.5</points>
<connection>
<GID>4903</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349.5,248.5,349.5,261</points>
<intersection>248.5 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349.5,252.5,353.5,252.5</points>
<connection>
<GID>4902</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347,261,349.5,261</points>
<connection>
<GID>4904</GID>
<name>OUT_0</name></connection>
<intersection>349.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3491</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389,251.5,391,251.5</points>
<connection>
<GID>4905</GID>
<name>OUT</name></connection>
<connection>
<GID>4906</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,248,393,248.5</points>
<connection>
<GID>4906</GID>
<name>IN_0</name></connection>
<intersection>248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,248,393,248</points>
<intersection>379 2</intersection>
<intersection>393 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379,248,379,261</points>
<intersection>248 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379,252.5,383,252.5</points>
<connection>
<GID>4905</GID>
<name>IN_0</name></connection>
<intersection>379 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377,261,379,261</points>
<connection>
<GID>4907</GID>
<name>OUT_0</name></connection>
<intersection>379 2</intersection></hsegment></shape></wire>
<wire>
<ID>3493</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420.5,251.5,422.5,251.5</points>
<connection>
<GID>4908</GID>
<name>OUT</name></connection>
<connection>
<GID>4909</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410.5,248.5,424.5,248.5</points>
<connection>
<GID>4909</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410.5,248.5,410.5,261</points>
<intersection>248.5 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410.5,252.5,414.5,252.5</points>
<connection>
<GID>4908</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408,261,410.5,261</points>
<connection>
<GID>4910</GID>
<name>OUT_0</name></connection>
<intersection>410.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3495</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451,251.5,453,251.5</points>
<connection>
<GID>4911</GID>
<name>OUT</name></connection>
<connection>
<GID>4912</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,248,455,248.5</points>
<connection>
<GID>4912</GID>
<name>IN_0</name></connection>
<intersection>248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,248,455,248</points>
<intersection>441 2</intersection>
<intersection>455 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441,248,441,261</points>
<intersection>248 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441,252.5,445,252.5</points>
<connection>
<GID>4911</GID>
<name>IN_0</name></connection>
<intersection>441 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439,261,441,261</points>
<connection>
<GID>4913</GID>
<name>OUT_0</name></connection>
<intersection>441 2</intersection></hsegment></shape></wire>
<wire>
<ID>3497</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482.5,251.5,484.5,251.5</points>
<connection>
<GID>4914</GID>
<name>OUT</name></connection>
<connection>
<GID>4915</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472.5,248.5,486.5,248.5</points>
<connection>
<GID>4915</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472.5,248.5,472.5,261</points>
<intersection>248.5 1</intersection>
<intersection>252.5 4</intersection>
<intersection>261 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472.5,252.5,476.5,252.5</points>
<connection>
<GID>4914</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470,261,472.5,261</points>
<connection>
<GID>4916</GID>
<name>OUT_0</name></connection>
<intersection>472.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,226.5,463,226.5</points>
<connection>
<GID>4943</GID>
<name>OUT</name></connection>
<connection>
<GID>4868</GID>
<name>clock</name></connection>
<connection>
<GID>4865</GID>
<name>clock</name></connection>
<connection>
<GID>4862</GID>
<name>clock</name></connection>
<connection>
<GID>4859</GID>
<name>clock</name></connection>
<connection>
<GID>4856</GID>
<name>clock</name></connection>
<connection>
<GID>4853</GID>
<name>clock</name></connection>
<connection>
<GID>4850</GID>
<name>clock</name></connection>
<connection>
<GID>4847</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,219,475.5,219</points>
<connection>
<GID>4845</GID>
<name>IN_1</name></connection>
<connection>
<GID>4848</GID>
<name>IN_1</name></connection>
<connection>
<GID>4851</GID>
<name>IN_1</name></connection>
<connection>
<GID>4854</GID>
<name>IN_1</name></connection>
<connection>
<GID>4857</GID>
<name>IN_1</name></connection>
<connection>
<GID>4860</GID>
<name>IN_1</name></connection>
<connection>
<GID>4863</GID>
<name>IN_1</name></connection>
<connection>
<GID>4866</GID>
<name>IN_1</name></connection>
<intersection>240 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240,219,240,221.5</points>
<connection>
<GID>4942</GID>
<name>OUT_0</name></connection>
<intersection>219 1</intersection></vsegment></shape></wire>
<wire>
<ID>3501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,209.5,462.5,209.5</points>
<connection>
<GID>4945</GID>
<name>OUT</name></connection>
<connection>
<GID>4844</GID>
<name>clock</name></connection>
<connection>
<GID>4841</GID>
<name>clock</name></connection>
<connection>
<GID>4838</GID>
<name>clock</name></connection>
<connection>
<GID>4835</GID>
<name>clock</name></connection>
<connection>
<GID>4832</GID>
<name>clock</name></connection>
<connection>
<GID>4829</GID>
<name>clock</name></connection>
<connection>
<GID>4826</GID>
<name>clock</name></connection>
<connection>
<GID>4812</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,202,241,204.5</points>
<intersection>202 2</intersection>
<intersection>204.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>241,202,475,202</points>
<connection>
<GID>4810</GID>
<name>IN_1</name></connection>
<connection>
<GID>4824</GID>
<name>IN_1</name></connection>
<connection>
<GID>4827</GID>
<name>IN_1</name></connection>
<connection>
<GID>4830</GID>
<name>IN_1</name></connection>
<connection>
<GID>4833</GID>
<name>IN_1</name></connection>
<connection>
<GID>4836</GID>
<name>IN_1</name></connection>
<connection>
<GID>4839</GID>
<name>IN_1</name></connection>
<connection>
<GID>4842</GID>
<name>IN_1</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>240,204.5,241,204.5</points>
<connection>
<GID>4944</GID>
<name>OUT_0</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>3503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,192.5,276.5,332.5</points>
<connection>
<GID>4822</GID>
<name>N_in0</name></connection>
<connection>
<GID>4814</GID>
<name>N_in1</name></connection>
<intersection>212.5 1</intersection>
<intersection>229.5 3</intersection>
<intersection>245.5 4</intersection>
<intersection>261 5</intersection>
<intersection>277.5 6</intersection>
<intersection>294.5 7</intersection>
<intersection>310.5 8</intersection>
<intersection>326 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276.5,212.5,277.5,212.5</points>
<connection>
<GID>4826</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276.5,326,280,326</points>
<connection>
<GID>5031</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>276.5,229.5,278,229.5</points>
<connection>
<GID>4850</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>276.5,245.5,278.5,245.5</points>
<connection>
<GID>4874</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>276.5,261,279,261</points>
<connection>
<GID>4898</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>276.5,277.5,278.5,277.5</points>
<connection>
<GID>4956</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>276.5,294.5,279,294.5</points>
<connection>
<GID>4983</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>276.5,310.5,279.5,310.5</points>
<connection>
<GID>5007</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,192.5,308.5,332.5</points>
<connection>
<GID>4823</GID>
<name>N_in0</name></connection>
<connection>
<GID>4829</GID>
<name>IN_0</name></connection>
<connection>
<GID>4815</GID>
<name>N_in1</name></connection>
<intersection>229.5 9</intersection>
<intersection>245.5 10</intersection>
<intersection>261 7</intersection>
<intersection>277.5 11</intersection>
<intersection>294.5 5</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308.5,326,311,326</points>
<connection>
<GID>5034</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,310.5,310.5,310.5</points>
<connection>
<GID>5010</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>308.5,294.5,310,294.5</points>
<connection>
<GID>4986</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>308.5,261,310,261</points>
<connection>
<GID>4901</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>308.5,229.5,309,229.5</points>
<connection>
<GID>4853</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>308.5,245.5,309.5,245.5</points>
<connection>
<GID>4877</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>308.5,277.5,309.5,277.5</points>
<connection>
<GID>4962</GID>
<name>IN_0</name></connection>
<intersection>308.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,193.5,339.5,332.5</points>
<connection>
<GID>4917</GID>
<name>N_in0</name></connection>
<connection>
<GID>4832</GID>
<name>IN_0</name></connection>
<connection>
<GID>4816</GID>
<name>N_in1</name></connection>
<intersection>229.5 38</intersection>
<intersection>245.5 21</intersection>
<intersection>261 7</intersection>
<intersection>277.5 20</intersection>
<intersection>294.5 5</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>339.5,326,342,326</points>
<connection>
<GID>5037</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,310.5,341.5,310.5</points>
<connection>
<GID>5013</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>339.5,294.5,341,294.5</points>
<connection>
<GID>4989</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>339.5,261,341,261</points>
<connection>
<GID>4904</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>339.5,277.5,340.5,277.5</points>
<connection>
<GID>4965</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>339.5,245.5,340.5,245.5</points>
<connection>
<GID>4880</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>339.5,229.5,340,229.5</points>
<connection>
<GID>4856</GID>
<name>IN_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370.5,229.5,370.5,332</points>
<connection>
<GID>4968</GID>
<name>IN_0</name></connection>
<connection>
<GID>4883</GID>
<name>IN_0</name></connection>
<connection>
<GID>4918</GID>
<name>N_in0</name></connection>
<intersection>229.5 9</intersection>
<intersection>261 7</intersection>
<intersection>294.5 5</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>370.5,326,372,326</points>
<connection>
<GID>5040</GID>
<name>IN_0</name></connection>
<intersection>370.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>370.5,310.5,371.5,310.5</points>
<connection>
<GID>5016</GID>
<name>IN_0</name></connection>
<intersection>370.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>370.5,294.5,371,294.5</points>
<connection>
<GID>4992</GID>
<name>IN_0</name></connection>
<intersection>370.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>370.5,261,371,261</points>
<connection>
<GID>4907</GID>
<name>IN_0</name></connection>
<intersection>370.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>369.5,229.5,370.5,229.5</points>
<connection>
<GID>4859</GID>
<name>IN_0</name></connection>
<intersection>369.5 10</intersection>
<intersection>370.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>369.5,194.5,369.5,229.5</points>
<connection>
<GID>4835</GID>
<name>IN_0</name></connection>
<connection>
<GID>4817</GID>
<name>N_in1</name></connection>
<intersection>229.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>3507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,195,400.5,332.5</points>
<connection>
<GID>4919</GID>
<name>N_in0</name></connection>
<connection>
<GID>4838</GID>
<name>IN_0</name></connection>
<connection>
<GID>4818</GID>
<name>N_in1</name></connection>
<intersection>229.5 13</intersection>
<intersection>245.5 11</intersection>
<intersection>261 9</intersection>
<intersection>277.5 7</intersection>
<intersection>294.5 5</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>400.5,326,403,326</points>
<connection>
<GID>5043</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>400.5,310.5,402.5,310.5</points>
<connection>
<GID>5019</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>400.5,294.5,402,294.5</points>
<connection>
<GID>4995</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>400.5,277.5,401.5,277.5</points>
<connection>
<GID>4971</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>400.5,261,402,261</points>
<connection>
<GID>4910</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>400.5,245.5,401.5,245.5</points>
<connection>
<GID>4886</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>400.5,229.5,401,229.5</points>
<connection>
<GID>4862</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,196,431.5,332.5</points>
<connection>
<GID>4920</GID>
<name>N_in0</name></connection>
<connection>
<GID>4841</GID>
<name>IN_0</name></connection>
<connection>
<GID>4820</GID>
<name>N_in1</name></connection>
<intersection>229.5 13</intersection>
<intersection>245.5 11</intersection>
<intersection>261 9</intersection>
<intersection>277.5 7</intersection>
<intersection>294.5 5</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,326,434,326</points>
<connection>
<GID>5046</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,310.5,433.5,310.5</points>
<connection>
<GID>5022</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>431.5,294.5,433,294.5</points>
<connection>
<GID>4998</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>431.5,277.5,432.5,277.5</points>
<connection>
<GID>4974</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>431.5,261,433,261</points>
<connection>
<GID>4913</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>431.5,245.5,432.5,245.5</points>
<connection>
<GID>4889</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>431.5,229.5,432,229.5</points>
<connection>
<GID>4865</GID>
<name>IN_0</name></connection>
<intersection>431.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,194,462.5,332</points>
<connection>
<GID>4921</GID>
<name>N_in0</name></connection>
<connection>
<GID>4844</GID>
<name>IN_0</name></connection>
<connection>
<GID>4819</GID>
<name>N_in1</name></connection>
<intersection>229.5 13</intersection>
<intersection>245.5 10</intersection>
<intersection>261 8</intersection>
<intersection>277.5 6</intersection>
<intersection>294.5 4</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>462.5,326,465,326</points>
<connection>
<GID>5049</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>462.5,310.5,464.5,310.5</points>
<connection>
<GID>5025</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>462.5,294.5,464,294.5</points>
<connection>
<GID>5001</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>462.5,277.5,463.5,277.5</points>
<connection>
<GID>4977</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>462.5,261,464,261</points>
<connection>
<GID>4916</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>462.5,245.5,463.5,245.5</points>
<connection>
<GID>4892</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>462.5,229.5,463,229.5</points>
<connection>
<GID>4868</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,184.5,274.5,339.5</points>
<connection>
<GID>4923</GID>
<name>N_in1</name></connection>
<connection>
<GID>4922</GID>
<name>N_in0</name></connection>
<intersection>205.5 13</intersection>
<intersection>222.5 12</intersection>
<intersection>238.5 11</intersection>
<intersection>254 10</intersection>
<intersection>270.5 9</intersection>
<intersection>287.5 8</intersection>
<intersection>303.5 7</intersection>
<intersection>319 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>271,319,274.5,319</points>
<connection>
<GID>5027</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>270.5,303.5,274.5,303.5</points>
<connection>
<GID>5003</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>270,287.5,274.5,287.5</points>
<connection>
<GID>4979</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>269.5,270.5,274.5,270.5</points>
<connection>
<GID>4947</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>270,254,274.5,254</points>
<connection>
<GID>4894</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>269.5,238.5,274.5,238.5</points>
<connection>
<GID>4870</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>269,222.5,274.5,222.5</points>
<connection>
<GID>4846</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>268.5,205.5,274.5,205.5</points>
<connection>
<GID>4811</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,205.5,305.5,339.5</points>
<connection>
<GID>4936</GID>
<name>N_in0</name></connection>
<intersection>205.5 13</intersection>
<intersection>222.5 12</intersection>
<intersection>238.5 11</intersection>
<intersection>254 10</intersection>
<intersection>270.5 9</intersection>
<intersection>287.5 8</intersection>
<intersection>303.5 7</intersection>
<intersection>319 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>302.5,319,305.5,319</points>
<connection>
<GID>5030</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>302,303.5,305.5,303.5</points>
<connection>
<GID>5006</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>301.5,287.5,305.5,287.5</points>
<connection>
<GID>4982</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>301,270.5,305.5,270.5</points>
<connection>
<GID>4954</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>301.5,254,305.5,254</points>
<connection>
<GID>4897</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>301,238.5,305.5,238.5</points>
<connection>
<GID>4873</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>300.5,222.5,305.5,222.5</points>
<connection>
<GID>4849</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>300,205.5,305.5,205.5</points>
<connection>
<GID>4825</GID>
<name>OUT_0</name></connection>
<intersection>303.5 22</intersection>
<intersection>305.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>303.5,192.5,303.5,205.5</points>
<connection>
<GID>5773</GID>
<name>N_in1</name></connection>
<intersection>205.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,185.5,337.5,339.5</points>
<connection>
<GID>4935</GID>
<name>N_in0</name></connection>
<connection>
<GID>4924</GID>
<name>N_in1</name></connection>
<intersection>205.5 13</intersection>
<intersection>222.5 12</intersection>
<intersection>238.5 11</intersection>
<intersection>254 10</intersection>
<intersection>270.5 9</intersection>
<intersection>287.5 8</intersection>
<intersection>303.5 7</intersection>
<intersection>319 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>333,319,337.5,319</points>
<connection>
<GID>5033</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>332.5,303.5,337.5,303.5</points>
<connection>
<GID>5009</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>332,287.5,337.5,287.5</points>
<connection>
<GID>4985</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>331.5,270.5,337.5,270.5</points>
<connection>
<GID>4960</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>332,254,337.5,254</points>
<connection>
<GID>4900</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>331.5,238.5,337.5,238.5</points>
<connection>
<GID>4876</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>331,222.5,337.5,222.5</points>
<connection>
<GID>4852</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>330.5,205.5,337.5,205.5</points>
<connection>
<GID>4828</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,186,368,339.5</points>
<connection>
<GID>4934</GID>
<name>N_in0</name></connection>
<connection>
<GID>4925</GID>
<name>N_in1</name></connection>
<intersection>205.5 18</intersection>
<intersection>222.5 17</intersection>
<intersection>238.5 16</intersection>
<intersection>254 15</intersection>
<intersection>270.5 14</intersection>
<intersection>287.5 13</intersection>
<intersection>303.5 12</intersection>
<intersection>319 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>364.5,319,368,319</points>
<connection>
<GID>5036</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>364,303.5,368,303.5</points>
<connection>
<GID>5012</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>363.5,287.5,368,287.5</points>
<connection>
<GID>4988</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>363,270.5,368,270.5</points>
<connection>
<GID>4964</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>363.5,254,368,254</points>
<connection>
<GID>4903</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>363,238.5,368,238.5</points>
<connection>
<GID>4879</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>362.5,222.5,368,222.5</points>
<connection>
<GID>4855</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>362,205.5,368,205.5</points>
<connection>
<GID>4831</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment></shape></wire>
<wire>
<ID>3514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398.5,186,398.5,339.5</points>
<connection>
<GID>4933</GID>
<name>N_in0</name></connection>
<connection>
<GID>4926</GID>
<name>N_in1</name></connection>
<intersection>205.5 9</intersection>
<intersection>222.5 10</intersection>
<intersection>238.5 11</intersection>
<intersection>254 12</intersection>
<intersection>270.5 13</intersection>
<intersection>287.5 14</intersection>
<intersection>303.5 15</intersection>
<intersection>319 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>391.5,205.5,398.5,205.5</points>
<connection>
<GID>4834</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>392,222.5,398.5,222.5</points>
<connection>
<GID>4858</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>392.5,238.5,398.5,238.5</points>
<connection>
<GID>4882</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>393,254,398.5,254</points>
<connection>
<GID>4906</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>392.5,270.5,398.5,270.5</points>
<connection>
<GID>4967</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>393,287.5,398.5,287.5</points>
<connection>
<GID>4991</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>393.5,303.5,398.5,303.5</points>
<connection>
<GID>5015</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>394,319,398.5,319</points>
<connection>
<GID>5039</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,186,429.5,339.5</points>
<connection>
<GID>4932</GID>
<name>N_in0</name></connection>
<connection>
<GID>4927</GID>
<name>N_in1</name></connection>
<intersection>205.5 6</intersection>
<intersection>222.5 7</intersection>
<intersection>238.5 8</intersection>
<intersection>254 9</intersection>
<intersection>270.5 10</intersection>
<intersection>287.5 11</intersection>
<intersection>303.5 12</intersection>
<intersection>319 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>423,205.5,429.5,205.5</points>
<connection>
<GID>4837</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>423.5,222.5,429.5,222.5</points>
<connection>
<GID>4861</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>424,238.5,429.5,238.5</points>
<connection>
<GID>4885</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>424.5,254,429.5,254</points>
<connection>
<GID>4909</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>424,270.5,429.5,270.5</points>
<connection>
<GID>4970</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>424.5,287.5,429.5,287.5</points>
<connection>
<GID>4994</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>425,303.5,429.5,303.5</points>
<connection>
<GID>5018</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>425.5,319,429.5,319</points>
<connection>
<GID>5042</GID>
<name>OUT_0</name></connection>
<intersection>429.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460.5,185.5,460.5,340.5</points>
<connection>
<GID>4931</GID>
<name>N_in0</name></connection>
<connection>
<GID>4928</GID>
<name>N_in1</name></connection>
<intersection>205.5 6</intersection>
<intersection>222.5 7</intersection>
<intersection>238.5 8</intersection>
<intersection>254 9</intersection>
<intersection>270.5 10</intersection>
<intersection>287.5 11</intersection>
<intersection>303.5 12</intersection>
<intersection>319 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>453.5,205.5,460.5,205.5</points>
<connection>
<GID>4840</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>454,222.5,460.5,222.5</points>
<connection>
<GID>4864</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>454.5,238.5,460.5,238.5</points>
<connection>
<GID>4888</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>455,254,460.5,254</points>
<connection>
<GID>4912</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>454.5,270.5,460.5,270.5</points>
<connection>
<GID>4973</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>455,287.5,460.5,287.5</points>
<connection>
<GID>4997</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>455.5,303.5,460.5,303.5</points>
<connection>
<GID>5021</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>456,319,460.5,319</points>
<connection>
<GID>5045</GID>
<name>OUT_0</name></connection>
<intersection>460.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,186,491,341</points>
<connection>
<GID>4930</GID>
<name>N_in0</name></connection>
<connection>
<GID>4929</GID>
<name>N_in1</name></connection>
<intersection>205.5 3</intersection>
<intersection>222.5 4</intersection>
<intersection>238.5 5</intersection>
<intersection>254 6</intersection>
<intersection>270.5 7</intersection>
<intersection>287.5 8</intersection>
<intersection>303.5 9</intersection>
<intersection>319 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>485,205.5,491,205.5</points>
<connection>
<GID>4843</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>485.5,222.5,491,222.5</points>
<connection>
<GID>4867</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>486,238.5,491,238.5</points>
<connection>
<GID>4891</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>486.5,254,491,254</points>
<connection>
<GID>4915</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>486,270.5,491,270.5</points>
<connection>
<GID>4976</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>486.5,287.5,491,287.5</points>
<connection>
<GID>5000</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>487,303.5,491,303.5</points>
<connection>
<GID>5024</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>487.5,319,491,319</points>
<connection>
<GID>5048</GID>
<name>OUT_0</name></connection>
<intersection>491 0</intersection></hsegment></shape></wire>
<wire>
<ID>3518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,271.5,199.5,320.5</points>
<intersection>271.5 2</intersection>
<intersection>320.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,320.5,238.5,320.5</points>
<connection>
<GID>4949</GID>
<name>ENABLE_0</name></connection>
<intersection>199.5 0</intersection>
<intersection>224.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,271.5,199.5,271.5</points>
<connection>
<GID>4937</GID>
<name>OUT_7</name></connection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>224.5,320.5,224.5,324</points>
<intersection>320.5 1</intersection>
<intersection>324 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,324,229,324</points>
<connection>
<GID>4950</GID>
<name>IN_0</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,270.5,201.5,305</points>
<intersection>270.5 2</intersection>
<intersection>305 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,305,238.5,305</points>
<intersection>201.5 0</intersection>
<intersection>224.5 4</intersection>
<intersection>238.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,270.5,201.5,270.5</points>
<connection>
<GID>4937</GID>
<name>OUT_6</name></connection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>238.5,304.5,238.5,305</points>
<connection>
<GID>4951</GID>
<name>ENABLE_0</name></connection>
<intersection>305 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>224.5,305,224.5,308.5</points>
<intersection>305 1</intersection>
<intersection>308.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,308.5,228.5,308.5</points>
<connection>
<GID>4953</GID>
<name>IN_0</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,269.5,203.5,292.5</points>
<intersection>269.5 2</intersection>
<intersection>292.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,292.5,228.5,292.5</points>
<connection>
<GID>4957</GID>
<name>IN_0</name></connection>
<intersection>203.5 0</intersection>
<intersection>224.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,269.5,203.5,269.5</points>
<connection>
<GID>4937</GID>
<name>OUT_5</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>224.5,288.5,224.5,292.5</points>
<intersection>288.5 4</intersection>
<intersection>292.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>224.5,288.5,238.5,288.5</points>
<connection>
<GID>4955</GID>
<name>ENABLE_0</name></connection>
<intersection>224.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,268.5,205.5,275.5</points>
<intersection>268.5 2</intersection>
<intersection>275.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,275.5,228.5,275.5</points>
<connection>
<GID>4961</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection>
<intersection>224.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,268.5,205.5,268.5</points>
<connection>
<GID>4937</GID>
<name>OUT_4</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>224.5,271.5,224.5,275.5</points>
<intersection>271.5 4</intersection>
<intersection>275.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>224.5,271.5,238.5,271.5</points>
<connection>
<GID>4959</GID>
<name>ENABLE_0</name></connection>
<intersection>224.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,255.5,205.5,267.5</points>
<intersection>255.5 1</intersection>
<intersection>267.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,255.5,237.5,255.5</points>
<connection>
<GID>4938</GID>
<name>ENABLE_0</name></connection>
<intersection>205.5 0</intersection>
<intersection>224.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,267.5,205.5,267.5</points>
<connection>
<GID>4937</GID>
<name>OUT_3</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>224.5,255.5,224.5,259</points>
<intersection>255.5 1</intersection>
<intersection>259 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,259,228.5,259</points>
<connection>
<GID>4939</GID>
<name>IN_0</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,239.5,203.5,266.5</points>
<intersection>239.5 1</intersection>
<intersection>266.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,239.5,237.5,239.5</points>
<connection>
<GID>4940</GID>
<name>ENABLE_0</name></connection>
<intersection>203.5 0</intersection>
<intersection>224.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,266.5,203.5,266.5</points>
<connection>
<GID>4937</GID>
<name>OUT_2</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>224.5,239.5,224.5,243.5</points>
<intersection>239.5 1</intersection>
<intersection>243.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,243.5,228.5,243.5</points>
<connection>
<GID>4941</GID>
<name>IN_0</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,224,201.5,265.5</points>
<intersection>224 1</intersection>
<intersection>265.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,224,237.5,224</points>
<intersection>201.5 0</intersection>
<intersection>224.5 4</intersection>
<intersection>237.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,265.5,201.5,265.5</points>
<connection>
<GID>4937</GID>
<name>OUT_1</name></connection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>237.5,223.5,237.5,224</points>
<connection>
<GID>4942</GID>
<name>ENABLE_0</name></connection>
<intersection>224 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>224.5,224,224.5,227.5</points>
<intersection>224 1</intersection>
<intersection>227.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,227.5,228.5,227.5</points>
<connection>
<GID>4943</GID>
<name>IN_0</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,206.5,199.5,264.5</points>
<intersection>206.5 1</intersection>
<intersection>264.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,206.5,237.5,206.5</points>
<connection>
<GID>4944</GID>
<name>ENABLE_0</name></connection>
<intersection>199.5 0</intersection>
<intersection>224.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198.5,264.5,199.5,264.5</points>
<connection>
<GID>4937</GID>
<name>OUT_0</name></connection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>224.5,206.5,224.5,210.5</points>
<intersection>206.5 1</intersection>
<intersection>210.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,210.5,228.5,210.5</points>
<connection>
<GID>4945</GID>
<name>IN_0</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3526</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>265.5,268,267.5,268</points>
<connection>
<GID>4946</GID>
<name>OUT</name></connection>
<connection>
<GID>4947</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,264.5,269.5,265</points>
<connection>
<GID>4947</GID>
<name>IN_0</name></connection>
<intersection>264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,264.5,269.5,264.5</points>
<intersection>255.5 2</intersection>
<intersection>269.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>255.5,264.5,255.5,277.5</points>
<intersection>264.5 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>255.5,269,259.5,269</points>
<connection>
<GID>4946</GID>
<name>IN_0</name></connection>
<intersection>255.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>253.5,277.5,255.5,277.5</points>
<connection>
<GID>4948</GID>
<name>OUT_0</name></connection>
<intersection>255.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3528</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297,268,299,268</points>
<connection>
<GID>4952</GID>
<name>OUT</name></connection>
<connection>
<GID>4954</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,265,301,265</points>
<connection>
<GID>4954</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287,265,287,277.5</points>
<intersection>265 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287,269,291,269</points>
<connection>
<GID>4952</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>284.5,277.5,287,277.5</points>
<connection>
<GID>4956</GID>
<name>OUT_0</name></connection>
<intersection>287 2</intersection></hsegment></shape></wire>
<wire>
<ID>3530</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>327.5,268,329.5,268</points>
<connection>
<GID>4958</GID>
<name>OUT</name></connection>
<connection>
<GID>4960</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,264.5,331.5,265</points>
<connection>
<GID>4960</GID>
<name>IN_0</name></connection>
<intersection>264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,264.5,331.5,264.5</points>
<intersection>317.5 2</intersection>
<intersection>331.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>317.5,264.5,317.5,277.5</points>
<intersection>264.5 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>317.5,269,321.5,269</points>
<connection>
<GID>4958</GID>
<name>IN_0</name></connection>
<intersection>317.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>315.5,277.5,317.5,277.5</points>
<connection>
<GID>4962</GID>
<name>OUT_0</name></connection>
<intersection>317.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3532</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359,268,361,268</points>
<connection>
<GID>4963</GID>
<name>OUT</name></connection>
<connection>
<GID>4964</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,265,363,265</points>
<connection>
<GID>4964</GID>
<name>IN_0</name></connection>
<intersection>349 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349,265,349,277.5</points>
<intersection>265 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349,269,353,269</points>
<connection>
<GID>4963</GID>
<name>IN_0</name></connection>
<intersection>349 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>346.5,277.5,349,277.5</points>
<connection>
<GID>4965</GID>
<name>OUT_0</name></connection>
<intersection>349 2</intersection></hsegment></shape></wire>
<wire>
<ID>3534</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>388.5,268,390.5,268</points>
<connection>
<GID>4966</GID>
<name>OUT</name></connection>
<connection>
<GID>4967</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392.5,264.5,392.5,265</points>
<connection>
<GID>4967</GID>
<name>IN_0</name></connection>
<intersection>264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378.5,264.5,392.5,264.5</points>
<intersection>378.5 2</intersection>
<intersection>392.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>378.5,264.5,378.5,277.5</points>
<intersection>264.5 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>378.5,269,382.5,269</points>
<connection>
<GID>4966</GID>
<name>IN_0</name></connection>
<intersection>378.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>376.5,277.5,378.5,277.5</points>
<connection>
<GID>4968</GID>
<name>OUT_0</name></connection>
<intersection>378.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3536</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420,268,422,268</points>
<connection>
<GID>4969</GID>
<name>OUT</name></connection>
<connection>
<GID>4970</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410,265,424,265</points>
<connection>
<GID>4970</GID>
<name>IN_0</name></connection>
<intersection>410 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410,265,410,277.5</points>
<intersection>265 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410,269,414,269</points>
<connection>
<GID>4969</GID>
<name>IN_0</name></connection>
<intersection>410 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>407.5,277.5,410,277.5</points>
<connection>
<GID>4971</GID>
<name>OUT_0</name></connection>
<intersection>410 2</intersection></hsegment></shape></wire>
<wire>
<ID>3538</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>450.5,268,452.5,268</points>
<connection>
<GID>4972</GID>
<name>OUT</name></connection>
<connection>
<GID>4973</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,264.5,454.5,265</points>
<connection>
<GID>4973</GID>
<name>IN_0</name></connection>
<intersection>264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>440.5,264.5,454.5,264.5</points>
<intersection>440.5 2</intersection>
<intersection>454.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>440.5,264.5,440.5,277.5</points>
<intersection>264.5 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>440.5,269,444.5,269</points>
<connection>
<GID>4972</GID>
<name>IN_0</name></connection>
<intersection>440.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>438.5,277.5,440.5,277.5</points>
<connection>
<GID>4974</GID>
<name>OUT_0</name></connection>
<intersection>440.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3540</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482,268,484,268</points>
<connection>
<GID>4975</GID>
<name>OUT</name></connection>
<connection>
<GID>4976</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3541</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472,265,486,265</points>
<connection>
<GID>4976</GID>
<name>IN_0</name></connection>
<intersection>472 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472,265,472,277.5</points>
<intersection>265 1</intersection>
<intersection>269 4</intersection>
<intersection>277.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472,269,476,269</points>
<connection>
<GID>4975</GID>
<name>IN_0</name></connection>
<intersection>472 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>469.5,277.5,472,277.5</points>
<connection>
<GID>4977</GID>
<name>OUT_0</name></connection>
<intersection>472 2</intersection></hsegment></shape></wire>
<wire>
<ID>3542</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266,285,268,285</points>
<connection>
<GID>4978</GID>
<name>OUT</name></connection>
<connection>
<GID>4979</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,281.5,270,282</points>
<connection>
<GID>4979</GID>
<name>IN_0</name></connection>
<intersection>281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,281.5,270,281.5</points>
<intersection>256 2</intersection>
<intersection>270 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256,281.5,256,294.5</points>
<intersection>281.5 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256,286,260,286</points>
<connection>
<GID>4978</GID>
<name>IN_0</name></connection>
<intersection>256 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254,294.5,256,294.5</points>
<connection>
<GID>4980</GID>
<name>OUT_0</name></connection>
<intersection>256 2</intersection></hsegment></shape></wire>
<wire>
<ID>3544</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297.5,285,299.5,285</points>
<connection>
<GID>4981</GID>
<name>OUT</name></connection>
<connection>
<GID>4982</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3545</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287.5,282,301.5,282</points>
<connection>
<GID>4982</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287.5,282,287.5,294.5</points>
<intersection>282 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,286,291.5,286</points>
<connection>
<GID>4981</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285,294.5,287.5,294.5</points>
<connection>
<GID>4983</GID>
<name>OUT_0</name></connection>
<intersection>287.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3546</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328,285,330,285</points>
<connection>
<GID>4984</GID>
<name>OUT</name></connection>
<connection>
<GID>4985</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,281.5,332,282</points>
<connection>
<GID>4985</GID>
<name>IN_0</name></connection>
<intersection>281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,281.5,332,281.5</points>
<intersection>318 2</intersection>
<intersection>332 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318,281.5,318,294.5</points>
<intersection>281.5 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318,286,322,286</points>
<connection>
<GID>4984</GID>
<name>IN_0</name></connection>
<intersection>318 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316,294.5,318,294.5</points>
<connection>
<GID>4986</GID>
<name>OUT_0</name></connection>
<intersection>318 2</intersection></hsegment></shape></wire>
<wire>
<ID>3548</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359.5,285,361.5,285</points>
<connection>
<GID>4987</GID>
<name>OUT</name></connection>
<connection>
<GID>4988</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349.5,282,363.5,282</points>
<connection>
<GID>4988</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349.5,282,349.5,294.5</points>
<intersection>282 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349.5,286,353.5,286</points>
<connection>
<GID>4987</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347,294.5,349.5,294.5</points>
<connection>
<GID>4989</GID>
<name>OUT_0</name></connection>
<intersection>349.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3550</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389,285,391,285</points>
<connection>
<GID>4990</GID>
<name>OUT</name></connection>
<connection>
<GID>4991</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,281.5,393,282</points>
<connection>
<GID>4991</GID>
<name>IN_0</name></connection>
<intersection>281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,281.5,393,281.5</points>
<intersection>379 2</intersection>
<intersection>393 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379,281.5,379,294.5</points>
<intersection>281.5 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379,286,383,286</points>
<connection>
<GID>4990</GID>
<name>IN_0</name></connection>
<intersection>379 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377,294.5,379,294.5</points>
<connection>
<GID>4992</GID>
<name>OUT_0</name></connection>
<intersection>379 2</intersection></hsegment></shape></wire>
<wire>
<ID>3552</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420.5,285,422.5,285</points>
<connection>
<GID>4993</GID>
<name>OUT</name></connection>
<connection>
<GID>4994</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3553</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410.5,282,424.5,282</points>
<connection>
<GID>4994</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410.5,282,410.5,294.5</points>
<intersection>282 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410.5,286,414.5,286</points>
<connection>
<GID>4993</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408,294.5,410.5,294.5</points>
<connection>
<GID>4995</GID>
<name>OUT_0</name></connection>
<intersection>410.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3554</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451,285,453,285</points>
<connection>
<GID>4996</GID>
<name>OUT</name></connection>
<connection>
<GID>4997</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,281.5,455,282</points>
<connection>
<GID>4997</GID>
<name>IN_0</name></connection>
<intersection>281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,281.5,455,281.5</points>
<intersection>441 2</intersection>
<intersection>455 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441,281.5,441,294.5</points>
<intersection>281.5 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441,286,445,286</points>
<connection>
<GID>4996</GID>
<name>IN_0</name></connection>
<intersection>441 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439,294.5,441,294.5</points>
<connection>
<GID>4998</GID>
<name>OUT_0</name></connection>
<intersection>441 2</intersection></hsegment></shape></wire>
<wire>
<ID>3556</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482.5,285,484.5,285</points>
<connection>
<GID>4999</GID>
<name>OUT</name></connection>
<connection>
<GID>5000</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472.5,282,486.5,282</points>
<connection>
<GID>5000</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472.5,282,472.5,294.5</points>
<intersection>282 1</intersection>
<intersection>286 4</intersection>
<intersection>294.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472.5,286,476.5,286</points>
<connection>
<GID>4999</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470,294.5,472.5,294.5</points>
<connection>
<GID>5001</GID>
<name>OUT_0</name></connection>
<intersection>472.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3558</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266.5,301,268.5,301</points>
<connection>
<GID>5002</GID>
<name>OUT</name></connection>
<connection>
<GID>5003</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,297.5,270.5,298</points>
<connection>
<GID>5003</GID>
<name>IN_0</name></connection>
<intersection>297.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,297.5,270.5,297.5</points>
<intersection>256.5 2</intersection>
<intersection>270.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256.5,297.5,256.5,310.5</points>
<intersection>297.5 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256.5,302,260.5,302</points>
<connection>
<GID>5002</GID>
<name>IN_0</name></connection>
<intersection>256.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254.5,310.5,256.5,310.5</points>
<connection>
<GID>5004</GID>
<name>OUT_0</name></connection>
<intersection>256.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3560</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,301,300,301</points>
<connection>
<GID>5005</GID>
<name>OUT</name></connection>
<connection>
<GID>5006</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,298,302,298</points>
<connection>
<GID>5006</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288,298,288,310.5</points>
<intersection>298 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,302,292,302</points>
<connection>
<GID>5005</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285.5,310.5,288,310.5</points>
<connection>
<GID>5007</GID>
<name>OUT_0</name></connection>
<intersection>288 2</intersection></hsegment></shape></wire>
<wire>
<ID>3562</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328.5,301,330.5,301</points>
<connection>
<GID>5008</GID>
<name>OUT</name></connection>
<connection>
<GID>5009</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,297.5,332.5,298</points>
<connection>
<GID>5009</GID>
<name>IN_0</name></connection>
<intersection>297.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,297.5,332.5,297.5</points>
<intersection>318.5 2</intersection>
<intersection>332.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318.5,297.5,318.5,310.5</points>
<intersection>297.5 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318.5,302,322.5,302</points>
<connection>
<GID>5008</GID>
<name>IN_0</name></connection>
<intersection>318.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316.5,310.5,318.5,310.5</points>
<connection>
<GID>5010</GID>
<name>OUT_0</name></connection>
<intersection>318.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3564</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360,301,362,301</points>
<connection>
<GID>5011</GID>
<name>OUT</name></connection>
<connection>
<GID>5012</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,298,364,298</points>
<connection>
<GID>5012</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,298,350,310.5</points>
<intersection>298 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350,302,354,302</points>
<connection>
<GID>5011</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347.5,310.5,350,310.5</points>
<connection>
<GID>5013</GID>
<name>OUT_0</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>3566</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389.5,301,391.5,301</points>
<connection>
<GID>5014</GID>
<name>OUT</name></connection>
<connection>
<GID>5015</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,297.5,393.5,298</points>
<connection>
<GID>5015</GID>
<name>IN_0</name></connection>
<intersection>297.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,297.5,393.5,297.5</points>
<intersection>379.5 2</intersection>
<intersection>393.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379.5,297.5,379.5,310.5</points>
<intersection>297.5 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379.5,302,383.5,302</points>
<connection>
<GID>5014</GID>
<name>IN_0</name></connection>
<intersection>379.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377.5,310.5,379.5,310.5</points>
<connection>
<GID>5016</GID>
<name>OUT_0</name></connection>
<intersection>379.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3568</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421,301,423,301</points>
<connection>
<GID>5017</GID>
<name>OUT</name></connection>
<connection>
<GID>5018</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3569</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411,298,425,298</points>
<connection>
<GID>5018</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411,298,411,310.5</points>
<intersection>298 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411,302,415,302</points>
<connection>
<GID>5017</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408.5,310.5,411,310.5</points>
<connection>
<GID>5019</GID>
<name>OUT_0</name></connection>
<intersection>411 2</intersection></hsegment></shape></wire>
<wire>
<ID>3570</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451.5,301,453.5,301</points>
<connection>
<GID>5020</GID>
<name>OUT</name></connection>
<connection>
<GID>5021</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,297.5,455.5,298</points>
<connection>
<GID>5021</GID>
<name>IN_0</name></connection>
<intersection>297.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,297.5,455.5,297.5</points>
<intersection>441.5 2</intersection>
<intersection>455.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441.5,297.5,441.5,310.5</points>
<intersection>297.5 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441.5,302,445.5,302</points>
<connection>
<GID>5020</GID>
<name>IN_0</name></connection>
<intersection>441.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439.5,310.5,441.5,310.5</points>
<connection>
<GID>5022</GID>
<name>OUT_0</name></connection>
<intersection>441.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3572</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483,301,485,301</points>
<connection>
<GID>5023</GID>
<name>OUT</name></connection>
<connection>
<GID>5024</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473,298,487,298</points>
<connection>
<GID>5024</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473,298,473,310.5</points>
<intersection>298 1</intersection>
<intersection>302 4</intersection>
<intersection>310.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473,302,477,302</points>
<connection>
<GID>5023</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470.5,310.5,473,310.5</points>
<connection>
<GID>5025</GID>
<name>OUT_0</name></connection>
<intersection>473 2</intersection></hsegment></shape></wire>
<wire>
<ID>3574</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267,316.5,269,316.5</points>
<connection>
<GID>5026</GID>
<name>OUT</name></connection>
<connection>
<GID>5027</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,313,271,313.5</points>
<connection>
<GID>5027</GID>
<name>IN_0</name></connection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,313,271,313</points>
<intersection>257 2</intersection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257,313,257,326</points>
<intersection>313 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,317.5,261,317.5</points>
<connection>
<GID>5026</GID>
<name>IN_0</name></connection>
<intersection>257 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255,326,257,326</points>
<connection>
<GID>5028</GID>
<name>OUT_0</name></connection>
<intersection>257 2</intersection></hsegment></shape></wire>
<wire>
<ID>3576</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,316.5,300.5,316.5</points>
<connection>
<GID>5029</GID>
<name>OUT</name></connection>
<connection>
<GID>5030</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288.5,313.5,302.5,313.5</points>
<connection>
<GID>5030</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288.5,313.5,288.5,326</points>
<intersection>313.5 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,317.5,292.5,317.5</points>
<connection>
<GID>5029</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,326,288.5,326</points>
<connection>
<GID>5031</GID>
<name>OUT_0</name></connection>
<intersection>288.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3578</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329,316.5,331,316.5</points>
<connection>
<GID>5032</GID>
<name>OUT</name></connection>
<connection>
<GID>5033</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,313,333,313.5</points>
<connection>
<GID>5033</GID>
<name>IN_0</name></connection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,313,333,313</points>
<intersection>319 2</intersection>
<intersection>333 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319,313,319,326</points>
<intersection>313 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,317.5,323,317.5</points>
<connection>
<GID>5032</GID>
<name>IN_0</name></connection>
<intersection>319 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317,326,319,326</points>
<connection>
<GID>5034</GID>
<name>OUT_0</name></connection>
<intersection>319 2</intersection></hsegment></shape></wire>
<wire>
<ID>3580</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360.5,316.5,362.5,316.5</points>
<connection>
<GID>5035</GID>
<name>OUT</name></connection>
<connection>
<GID>5036</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350.5,313.5,364.5,313.5</points>
<connection>
<GID>5036</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,313.5,350.5,326</points>
<intersection>313.5 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350.5,317.5,354.5,317.5</points>
<connection>
<GID>5035</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348,326,350.5,326</points>
<connection>
<GID>5037</GID>
<name>OUT_0</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3582</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390,316.5,392,316.5</points>
<connection>
<GID>5038</GID>
<name>OUT</name></connection>
<connection>
<GID>5039</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,313,394,313.5</points>
<connection>
<GID>5039</GID>
<name>IN_0</name></connection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,313,394,313</points>
<intersection>380 2</intersection>
<intersection>394 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380,313,380,326</points>
<intersection>313 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,317.5,384,317.5</points>
<connection>
<GID>5038</GID>
<name>IN_0</name></connection>
<intersection>380 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378,326,380,326</points>
<connection>
<GID>5040</GID>
<name>OUT_0</name></connection>
<intersection>380 2</intersection></hsegment></shape></wire>
<wire>
<ID>3584</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421.5,316.5,423.5,316.5</points>
<connection>
<GID>5041</GID>
<name>OUT</name></connection>
<connection>
<GID>5042</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411.5,313.5,425.5,313.5</points>
<connection>
<GID>5042</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411.5,313.5,411.5,326</points>
<intersection>313.5 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411.5,317.5,415.5,317.5</points>
<connection>
<GID>5041</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409,326,411.5,326</points>
<connection>
<GID>5043</GID>
<name>OUT_0</name></connection>
<intersection>411.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3586</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452,316.5,454,316.5</points>
<connection>
<GID>5044</GID>
<name>OUT</name></connection>
<connection>
<GID>5045</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,313,456,313.5</points>
<connection>
<GID>5045</GID>
<name>IN_0</name></connection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,313,456,313</points>
<intersection>442 2</intersection>
<intersection>456 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442,313,442,326</points>
<intersection>313 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442,317.5,446,317.5</points>
<connection>
<GID>5044</GID>
<name>IN_0</name></connection>
<intersection>442 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,326,442,326</points>
<connection>
<GID>5046</GID>
<name>OUT_0</name></connection>
<intersection>442 2</intersection></hsegment></shape></wire>
<wire>
<ID>3588</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483.5,316.5,485.5,316.5</points>
<connection>
<GID>5047</GID>
<name>OUT</name></connection>
<connection>
<GID>5048</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3589</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473.5,313.5,487.5,313.5</points>
<connection>
<GID>5048</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473.5,313.5,473.5,326</points>
<intersection>313.5 1</intersection>
<intersection>317.5 4</intersection>
<intersection>326 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473.5,317.5,477.5,317.5</points>
<connection>
<GID>5047</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471,326,473.5,326</points>
<connection>
<GID>5049</GID>
<name>OUT_0</name></connection>
<intersection>473.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,193,245.5,332.5</points>
<connection>
<GID>4821</GID>
<name>N_in0</name></connection>
<connection>
<GID>4813</GID>
<name>N_in1</name></connection>
<intersection>212.5 14</intersection>
<intersection>229.5 12</intersection>
<intersection>245.5 10</intersection>
<intersection>261 8</intersection>
<intersection>277.5 6</intersection>
<intersection>294.5 4</intersection>
<intersection>310.5 2</intersection>
<intersection>326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,326,249,326</points>
<connection>
<GID>5028</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>245.5,310.5,248.5,310.5</points>
<connection>
<GID>5004</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>245.5,294.5,248,294.5</points>
<connection>
<GID>4980</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>245.5,277.5,247.5,277.5</points>
<connection>
<GID>4948</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>245.5,261,248,261</points>
<connection>
<GID>4895</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>245.5,245.5,247.5,245.5</points>
<connection>
<GID>4871</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>245.5,229.5,247,229.5</points>
<connection>
<GID>4847</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>245.5,212.5,246.5,212.5</points>
<connection>
<GID>4812</GID>
<name>IN_0</name></connection>
<intersection>245.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3591</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,315.5,477.5,315.5</points>
<connection>
<GID>5026</GID>
<name>IN_1</name></connection>
<connection>
<GID>5029</GID>
<name>IN_1</name></connection>
<connection>
<GID>5032</GID>
<name>IN_1</name></connection>
<connection>
<GID>5035</GID>
<name>IN_1</name></connection>
<connection>
<GID>5038</GID>
<name>IN_1</name></connection>
<connection>
<GID>5041</GID>
<name>IN_1</name></connection>
<connection>
<GID>5044</GID>
<name>IN_1</name></connection>
<connection>
<GID>5047</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,315.5,241,318.5</points>
<connection>
<GID>4949</GID>
<name>OUT_0</name></connection>
<intersection>315.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3592</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,323,465,323</points>
<connection>
<GID>4950</GID>
<name>OUT</name></connection>
<connection>
<GID>5028</GID>
<name>clock</name></connection>
<connection>
<GID>5031</GID>
<name>clock</name></connection>
<connection>
<GID>5034</GID>
<name>clock</name></connection>
<connection>
<GID>5037</GID>
<name>clock</name></connection>
<connection>
<GID>5040</GID>
<name>clock</name></connection>
<connection>
<GID>5043</GID>
<name>clock</name></connection>
<connection>
<GID>5046</GID>
<name>clock</name></connection>
<connection>
<GID>5049</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3761</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>260.5,-891,262.5,-891</points>
<connection>
<GID>5290</GID>
<name>OUT</name></connection>
<connection>
<GID>5291</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-894.5,264.5,-894</points>
<connection>
<GID>5291</GID>
<name>IN_0</name></connection>
<intersection>-894.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-894.5,264.5,-894.5</points>
<intersection>250.5 2</intersection>
<intersection>264.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>250.5,-894.5,250.5,-881.5</points>
<intersection>-894.5 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>250.5,-890,254.5,-890</points>
<connection>
<GID>5290</GID>
<name>IN_0</name></connection>
<intersection>250.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>248.5,-881.5,250.5,-881.5</points>
<connection>
<GID>5292</GID>
<name>OUT_0</name></connection>
<intersection>250.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3763</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237,-794,473,-794</points>
<connection>
<GID>5482</GID>
<name>IN_1</name></connection>
<connection>
<GID>5485</GID>
<name>IN_1</name></connection>
<connection>
<GID>5488</GID>
<name>IN_1</name></connection>
<connection>
<GID>5491</GID>
<name>IN_1</name></connection>
<connection>
<GID>5494</GID>
<name>IN_1</name></connection>
<connection>
<GID>5497</GID>
<name>IN_1</name></connection>
<connection>
<GID>5500</GID>
<name>IN_1</name></connection>
<connection>
<GID>5503</GID>
<name>IN_1</name></connection>
<intersection>237 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>237,-794,237,-791.5</points>
<connection>
<GID>5431</GID>
<name>OUT_0</name></connection>
<intersection>-794 1</intersection></vsegment></shape></wire>
<wire>
<ID>3764</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-786.5,460.5,-786.5</points>
<connection>
<GID>5433</GID>
<name>OUT</name></connection>
<connection>
<GID>5484</GID>
<name>clock</name></connection>
<connection>
<GID>5487</GID>
<name>clock</name></connection>
<connection>
<GID>5490</GID>
<name>clock</name></connection>
<connection>
<GID>5493</GID>
<name>clock</name></connection>
<connection>
<GID>5496</GID>
<name>clock</name></connection>
<connection>
<GID>5499</GID>
<name>clock</name></connection>
<connection>
<GID>5502</GID>
<name>clock</name></connection>
<connection>
<GID>5505</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3765</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237,-810,472.5,-810</points>
<connection>
<GID>5458</GID>
<name>IN_1</name></connection>
<connection>
<GID>5461</GID>
<name>IN_1</name></connection>
<connection>
<GID>5464</GID>
<name>IN_1</name></connection>
<connection>
<GID>5467</GID>
<name>IN_1</name></connection>
<connection>
<GID>5470</GID>
<name>IN_1</name></connection>
<connection>
<GID>5473</GID>
<name>IN_1</name></connection>
<connection>
<GID>5476</GID>
<name>IN_1</name></connection>
<connection>
<GID>5479</GID>
<name>IN_1</name></connection>
<intersection>237 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>237,-810,237,-807.5</points>
<connection>
<GID>5435</GID>
<name>OUT_0</name></connection>
<intersection>-810 1</intersection></vsegment></shape></wire>
<wire>
<ID>3766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-802.5,460,-802.5</points>
<connection>
<GID>5437</GID>
<name>OUT</name></connection>
<connection>
<GID>5460</GID>
<name>clock</name></connection>
<connection>
<GID>5463</GID>
<name>clock</name></connection>
<connection>
<GID>5466</GID>
<name>clock</name></connection>
<connection>
<GID>5469</GID>
<name>clock</name></connection>
<connection>
<GID>5472</GID>
<name>clock</name></connection>
<connection>
<GID>5475</GID>
<name>clock</name></connection>
<connection>
<GID>5478</GID>
<name>clock</name></connection>
<connection>
<GID>5481</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3767</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-819.5,459.5,-819.5</points>
<connection>
<GID>5457</GID>
<name>clock</name></connection>
<connection>
<GID>5454</GID>
<name>clock</name></connection>
<connection>
<GID>5451</GID>
<name>clock</name></connection>
<connection>
<GID>5448</GID>
<name>clock</name></connection>
<connection>
<GID>5445</GID>
<name>clock</name></connection>
<connection>
<GID>5442</GID>
<name>clock</name></connection>
<connection>
<GID>5441</GID>
<name>OUT</name></connection>
<connection>
<GID>5436</GID>
<name>clock</name></connection>
<connection>
<GID>5428</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3768</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237,-827,472,-827</points>
<connection>
<GID>5426</GID>
<name>IN_1</name></connection>
<connection>
<GID>5432</GID>
<name>IN_1</name></connection>
<connection>
<GID>5438</GID>
<name>IN_1</name></connection>
<connection>
<GID>5443</GID>
<name>IN_1</name></connection>
<connection>
<GID>5446</GID>
<name>IN_1</name></connection>
<connection>
<GID>5449</GID>
<name>IN_1</name></connection>
<connection>
<GID>5452</GID>
<name>IN_1</name></connection>
<connection>
<GID>5455</GID>
<name>IN_1</name></connection>
<intersection>237 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>237,-827,237,-824.5</points>
<connection>
<GID>5439</GID>
<name>OUT_0</name></connection>
<intersection>-827 1</intersection></vsegment></shape></wire>
<wire>
<ID>3769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-836,460,-836</points>
<connection>
<GID>5419</GID>
<name>OUT</name></connection>
<connection>
<GID>5396</GID>
<name>clock</name></connection>
<connection>
<GID>5393</GID>
<name>clock</name></connection>
<connection>
<GID>5390</GID>
<name>clock</name></connection>
<connection>
<GID>5387</GID>
<name>clock</name></connection>
<connection>
<GID>5384</GID>
<name>clock</name></connection>
<connection>
<GID>5381</GID>
<name>clock</name></connection>
<connection>
<GID>5378</GID>
<name>clock</name></connection>
<connection>
<GID>5375</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,-843.5,472.5,-843.5</points>
<connection>
<GID>5373</GID>
<name>IN_1</name></connection>
<connection>
<GID>5376</GID>
<name>IN_1</name></connection>
<connection>
<GID>5379</GID>
<name>IN_1</name></connection>
<connection>
<GID>5382</GID>
<name>IN_1</name></connection>
<connection>
<GID>5385</GID>
<name>IN_1</name></connection>
<connection>
<GID>5388</GID>
<name>IN_1</name></connection>
<connection>
<GID>5391</GID>
<name>IN_1</name></connection>
<connection>
<GID>5394</GID>
<name>IN_1</name></connection>
<intersection>236 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>236,-843.5,236,-840.5</points>
<connection>
<GID>5418</GID>
<name>OUT_0</name></connection>
<intersection>-843.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3771</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-851.5,459.5,-851.5</points>
<connection>
<GID>5421</GID>
<name>OUT</name></connection>
<connection>
<GID>5372</GID>
<name>clock</name></connection>
<connection>
<GID>5369</GID>
<name>clock</name></connection>
<connection>
<GID>5366</GID>
<name>clock</name></connection>
<connection>
<GID>5363</GID>
<name>clock</name></connection>
<connection>
<GID>5360</GID>
<name>clock</name></connection>
<connection>
<GID>5357</GID>
<name>clock</name></connection>
<connection>
<GID>5354</GID>
<name>clock</name></connection>
<connection>
<GID>5351</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3772</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,-859,472,-859</points>
<connection>
<GID>5349</GID>
<name>IN_1</name></connection>
<connection>
<GID>5352</GID>
<name>IN_1</name></connection>
<connection>
<GID>5355</GID>
<name>IN_1</name></connection>
<connection>
<GID>5358</GID>
<name>IN_1</name></connection>
<connection>
<GID>5361</GID>
<name>IN_1</name></connection>
<connection>
<GID>5364</GID>
<name>IN_1</name></connection>
<connection>
<GID>5367</GID>
<name>IN_1</name></connection>
<connection>
<GID>5370</GID>
<name>IN_1</name></connection>
<intersection>236 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>236,-859,236,-856.5</points>
<connection>
<GID>5420</GID>
<name>OUT_0</name></connection>
<intersection>-859 1</intersection></vsegment></shape></wire>
<wire>
<ID>3773</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>292,-891,294,-891</points>
<connection>
<GID>5304</GID>
<name>OUT</name></connection>
<connection>
<GID>5305</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3774</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>282,-894,296,-894</points>
<connection>
<GID>5305</GID>
<name>IN_0</name></connection>
<intersection>282 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282,-894,282,-881.5</points>
<intersection>-894 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>282,-890,286,-890</points>
<connection>
<GID>5304</GID>
<name>IN_0</name></connection>
<intersection>282 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>279.5,-881.5,282,-881.5</points>
<connection>
<GID>5306</GID>
<name>OUT_0</name></connection>
<intersection>282 2</intersection></hsegment></shape></wire>
<wire>
<ID>3775</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>322.5,-891,324.5,-891</points>
<connection>
<GID>5307</GID>
<name>OUT</name></connection>
<connection>
<GID>5308</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-894.5,326.5,-894</points>
<connection>
<GID>5308</GID>
<name>IN_0</name></connection>
<intersection>-894.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-894.5,326.5,-894.5</points>
<intersection>312.5 2</intersection>
<intersection>326.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>312.5,-894.5,312.5,-881.5</points>
<intersection>-894.5 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>312.5,-890,316.5,-890</points>
<connection>
<GID>5307</GID>
<name>IN_0</name></connection>
<intersection>312.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>310.5,-881.5,312.5,-881.5</points>
<connection>
<GID>5309</GID>
<name>OUT_0</name></connection>
<intersection>312.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3777</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>354,-891,356,-891</points>
<connection>
<GID>5310</GID>
<name>OUT</name></connection>
<connection>
<GID>5311</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3778</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>344,-894,358,-894</points>
<connection>
<GID>5311</GID>
<name>IN_0</name></connection>
<intersection>344 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>344,-894,344,-881.5</points>
<intersection>-894 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>344,-890,348,-890</points>
<connection>
<GID>5310</GID>
<name>IN_0</name></connection>
<intersection>344 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>341.5,-881.5,344,-881.5</points>
<connection>
<GID>5312</GID>
<name>OUT_0</name></connection>
<intersection>344 2</intersection></hsegment></shape></wire>
<wire>
<ID>3779</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>383.5,-891,385.5,-891</points>
<connection>
<GID>5313</GID>
<name>OUT</name></connection>
<connection>
<GID>5314</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387.5,-894.5,387.5,-894</points>
<connection>
<GID>5314</GID>
<name>IN_0</name></connection>
<intersection>-894.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373.5,-894.5,387.5,-894.5</points>
<intersection>373.5 2</intersection>
<intersection>387.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>373.5,-894.5,373.5,-881.5</points>
<intersection>-894.5 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>373.5,-890,377.5,-890</points>
<connection>
<GID>5313</GID>
<name>IN_0</name></connection>
<intersection>373.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>371.5,-881.5,373.5,-881.5</points>
<connection>
<GID>5315</GID>
<name>OUT_0</name></connection>
<intersection>373.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3781</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>415,-891,417,-891</points>
<connection>
<GID>5316</GID>
<name>OUT</name></connection>
<connection>
<GID>5317</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3782</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>405,-894,419,-894</points>
<connection>
<GID>5317</GID>
<name>IN_0</name></connection>
<intersection>405 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>405,-894,405,-881.5</points>
<intersection>-894 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>405,-890,409,-890</points>
<connection>
<GID>5316</GID>
<name>IN_0</name></connection>
<intersection>405 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>402.5,-881.5,405,-881.5</points>
<connection>
<GID>5318</GID>
<name>OUT_0</name></connection>
<intersection>405 2</intersection></hsegment></shape></wire>
<wire>
<ID>3783</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>445.5,-891,447.5,-891</points>
<connection>
<GID>5319</GID>
<name>OUT</name></connection>
<connection>
<GID>5320</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-894.5,449.5,-894</points>
<connection>
<GID>5320</GID>
<name>IN_0</name></connection>
<intersection>-894.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435.5,-894.5,449.5,-894.5</points>
<intersection>435.5 2</intersection>
<intersection>449.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>435.5,-894.5,435.5,-881.5</points>
<intersection>-894.5 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>435.5,-890,439.5,-890</points>
<connection>
<GID>5319</GID>
<name>IN_0</name></connection>
<intersection>435.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>433.5,-881.5,435.5,-881.5</points>
<connection>
<GID>5321</GID>
<name>OUT_0</name></connection>
<intersection>435.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3785</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>477,-891,479,-891</points>
<connection>
<GID>5322</GID>
<name>OUT</name></connection>
<connection>
<GID>5323</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3786</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>467,-894,481,-894</points>
<connection>
<GID>5323</GID>
<name>IN_0</name></connection>
<intersection>467 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>467,-894,467,-881.5</points>
<intersection>-894 1</intersection>
<intersection>-890 4</intersection>
<intersection>-881.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>467,-890,471,-890</points>
<connection>
<GID>5322</GID>
<name>IN_0</name></connection>
<intersection>467 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>464.5,-881.5,467,-881.5</points>
<connection>
<GID>5324</GID>
<name>OUT_0</name></connection>
<intersection>467 2</intersection></hsegment></shape></wire>
<wire>
<ID>3787</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>261,-874,263,-874</points>
<connection>
<GID>5325</GID>
<name>OUT</name></connection>
<connection>
<GID>5326</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265,-877.5,265,-877</points>
<connection>
<GID>5326</GID>
<name>IN_0</name></connection>
<intersection>-877.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251,-877.5,265,-877.5</points>
<intersection>251 2</intersection>
<intersection>265 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>251,-877.5,251,-864.5</points>
<intersection>-877.5 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>251,-873,255,-873</points>
<connection>
<GID>5325</GID>
<name>IN_0</name></connection>
<intersection>251 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>249,-864.5,251,-864.5</points>
<connection>
<GID>5327</GID>
<name>OUT_0</name></connection>
<intersection>251 2</intersection></hsegment></shape></wire>
<wire>
<ID>3789</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>292.5,-874,294.5,-874</points>
<connection>
<GID>5328</GID>
<name>OUT</name></connection>
<connection>
<GID>5329</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3790</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>282.5,-877,296.5,-877</points>
<connection>
<GID>5329</GID>
<name>IN_0</name></connection>
<intersection>282.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>282.5,-877,282.5,-864.5</points>
<intersection>-877 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>282.5,-873,286.5,-873</points>
<connection>
<GID>5328</GID>
<name>IN_0</name></connection>
<intersection>282.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>280,-864.5,282.5,-864.5</points>
<connection>
<GID>5330</GID>
<name>OUT_0</name></connection>
<intersection>282.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3791</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>323,-874,325,-874</points>
<connection>
<GID>5331</GID>
<name>OUT</name></connection>
<connection>
<GID>5332</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327,-877.5,327,-877</points>
<connection>
<GID>5332</GID>
<name>IN_0</name></connection>
<intersection>-877.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-877.5,327,-877.5</points>
<intersection>313 2</intersection>
<intersection>327 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>313,-877.5,313,-864.5</points>
<intersection>-877.5 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>313,-873,317,-873</points>
<connection>
<GID>5331</GID>
<name>IN_0</name></connection>
<intersection>313 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>311,-864.5,313,-864.5</points>
<connection>
<GID>5333</GID>
<name>OUT_0</name></connection>
<intersection>313 2</intersection></hsegment></shape></wire>
<wire>
<ID>2249</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266.5,-358,268.5,-358</points>
<connection>
<GID>3130</GID>
<name>OUT</name></connection>
<connection>
<GID>3131</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3793</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>354.5,-874,356.5,-874</points>
<connection>
<GID>5334</GID>
<name>OUT</name></connection>
<connection>
<GID>5335</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-361.5,270.5,-361</points>
<connection>
<GID>3131</GID>
<name>IN_0</name></connection>
<intersection>-361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,-361.5,270.5,-361.5</points>
<intersection>256.5 2</intersection>
<intersection>270.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256.5,-361.5,256.5,-348.5</points>
<intersection>-361.5 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256.5,-357,260.5,-357</points>
<connection>
<GID>3130</GID>
<name>IN_0</name></connection>
<intersection>256.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254.5,-348.5,256.5,-348.5</points>
<connection>
<GID>3132</GID>
<name>OUT_0</name></connection>
<intersection>256.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3794</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>344.5,-877,358.5,-877</points>
<connection>
<GID>5335</GID>
<name>IN_0</name></connection>
<intersection>344.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>344.5,-877,344.5,-864.5</points>
<intersection>-877 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>344.5,-873,348.5,-873</points>
<connection>
<GID>5334</GID>
<name>IN_0</name></connection>
<intersection>344.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>342,-864.5,344.5,-864.5</points>
<connection>
<GID>5336</GID>
<name>OUT_0</name></connection>
<intersection>344.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-261,479,-261</points>
<connection>
<GID>3322</GID>
<name>IN_1</name></connection>
<connection>
<GID>3325</GID>
<name>IN_1</name></connection>
<connection>
<GID>3328</GID>
<name>IN_1</name></connection>
<connection>
<GID>3331</GID>
<name>IN_1</name></connection>
<connection>
<GID>3334</GID>
<name>IN_1</name></connection>
<connection>
<GID>3337</GID>
<name>IN_1</name></connection>
<connection>
<GID>3340</GID>
<name>IN_1</name></connection>
<connection>
<GID>3343</GID>
<name>IN_1</name></connection>
<intersection>243 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243,-261,243,-258.5</points>
<connection>
<GID>3271</GID>
<name>OUT_0</name></connection>
<intersection>-261 1</intersection></vsegment></shape></wire>
<wire>
<ID>3795</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>384,-874,386,-874</points>
<connection>
<GID>5337</GID>
<name>OUT</name></connection>
<connection>
<GID>5338</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-253.5,466.5,-253.5</points>
<connection>
<GID>3273</GID>
<name>OUT</name></connection>
<connection>
<GID>3324</GID>
<name>clock</name></connection>
<connection>
<GID>3327</GID>
<name>clock</name></connection>
<connection>
<GID>3330</GID>
<name>clock</name></connection>
<connection>
<GID>3333</GID>
<name>clock</name></connection>
<connection>
<GID>3336</GID>
<name>clock</name></connection>
<connection>
<GID>3339</GID>
<name>clock</name></connection>
<connection>
<GID>3342</GID>
<name>clock</name></connection>
<connection>
<GID>3345</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388,-877.5,388,-877</points>
<connection>
<GID>5338</GID>
<name>IN_0</name></connection>
<intersection>-877.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374,-877.5,388,-877.5</points>
<intersection>374 2</intersection>
<intersection>388 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>374,-877.5,374,-864.5</points>
<intersection>-877.5 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>374,-873,378,-873</points>
<connection>
<GID>5337</GID>
<name>IN_0</name></connection>
<intersection>374 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>372,-864.5,374,-864.5</points>
<connection>
<GID>5339</GID>
<name>OUT_0</name></connection>
<intersection>374 2</intersection></hsegment></shape></wire>
<wire>
<ID>2253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-277,478.5,-277</points>
<connection>
<GID>3298</GID>
<name>IN_1</name></connection>
<connection>
<GID>3301</GID>
<name>IN_1</name></connection>
<connection>
<GID>3304</GID>
<name>IN_1</name></connection>
<connection>
<GID>3307</GID>
<name>IN_1</name></connection>
<connection>
<GID>3310</GID>
<name>IN_1</name></connection>
<connection>
<GID>3313</GID>
<name>IN_1</name></connection>
<connection>
<GID>3316</GID>
<name>IN_1</name></connection>
<connection>
<GID>3319</GID>
<name>IN_1</name></connection>
<intersection>243 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243,-277,243,-274.5</points>
<connection>
<GID>3275</GID>
<name>OUT_0</name></connection>
<intersection>-277 1</intersection></vsegment></shape></wire>
<wire>
<ID>3797</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>415.5,-874,417.5,-874</points>
<connection>
<GID>5340</GID>
<name>OUT</name></connection>
<connection>
<GID>5341</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-269.5,466,-269.5</points>
<connection>
<GID>3277</GID>
<name>OUT</name></connection>
<connection>
<GID>3300</GID>
<name>clock</name></connection>
<connection>
<GID>3303</GID>
<name>clock</name></connection>
<connection>
<GID>3306</GID>
<name>clock</name></connection>
<connection>
<GID>3309</GID>
<name>clock</name></connection>
<connection>
<GID>3312</GID>
<name>clock</name></connection>
<connection>
<GID>3315</GID>
<name>clock</name></connection>
<connection>
<GID>3318</GID>
<name>clock</name></connection>
<connection>
<GID>3321</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3798</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>405.5,-877,419.5,-877</points>
<connection>
<GID>5341</GID>
<name>IN_0</name></connection>
<intersection>405.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>405.5,-877,405.5,-864.5</points>
<intersection>-877 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>405.5,-873,409.5,-873</points>
<connection>
<GID>5340</GID>
<name>IN_0</name></connection>
<intersection>405.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>403,-864.5,405.5,-864.5</points>
<connection>
<GID>5342</GID>
<name>OUT_0</name></connection>
<intersection>405.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-286.5,465.5,-286.5</points>
<connection>
<GID>3297</GID>
<name>clock</name></connection>
<connection>
<GID>3294</GID>
<name>clock</name></connection>
<connection>
<GID>3291</GID>
<name>clock</name></connection>
<connection>
<GID>3288</GID>
<name>clock</name></connection>
<connection>
<GID>3285</GID>
<name>clock</name></connection>
<connection>
<GID>3282</GID>
<name>clock</name></connection>
<connection>
<GID>3281</GID>
<name>OUT</name></connection>
<connection>
<GID>3276</GID>
<name>clock</name></connection>
<connection>
<GID>3268</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3799</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>446,-874,448,-874</points>
<connection>
<GID>5343</GID>
<name>OUT</name></connection>
<connection>
<GID>5344</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-294,478,-294</points>
<connection>
<GID>3266</GID>
<name>IN_1</name></connection>
<connection>
<GID>3272</GID>
<name>IN_1</name></connection>
<connection>
<GID>3278</GID>
<name>IN_1</name></connection>
<connection>
<GID>3283</GID>
<name>IN_1</name></connection>
<connection>
<GID>3286</GID>
<name>IN_1</name></connection>
<connection>
<GID>3289</GID>
<name>IN_1</name></connection>
<connection>
<GID>3292</GID>
<name>IN_1</name></connection>
<connection>
<GID>3295</GID>
<name>IN_1</name></connection>
<intersection>243 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243,-294,243,-291.5</points>
<connection>
<GID>3279</GID>
<name>OUT_0</name></connection>
<intersection>-294 1</intersection></vsegment></shape></wire>
<wire>
<ID>3800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,-877.5,450,-877</points>
<connection>
<GID>5344</GID>
<name>IN_0</name></connection>
<intersection>-877.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436,-877.5,450,-877.5</points>
<intersection>436 2</intersection>
<intersection>450 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>436,-877.5,436,-864.5</points>
<intersection>-877.5 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>436,-873,440,-873</points>
<connection>
<GID>5343</GID>
<name>IN_0</name></connection>
<intersection>436 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>434,-864.5,436,-864.5</points>
<connection>
<GID>5345</GID>
<name>OUT_0</name></connection>
<intersection>436 2</intersection></hsegment></shape></wire>
<wire>
<ID>2257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-303,466,-303</points>
<connection>
<GID>3259</GID>
<name>OUT</name></connection>
<connection>
<GID>3236</GID>
<name>clock</name></connection>
<connection>
<GID>3233</GID>
<name>clock</name></connection>
<connection>
<GID>3230</GID>
<name>clock</name></connection>
<connection>
<GID>3227</GID>
<name>clock</name></connection>
<connection>
<GID>3224</GID>
<name>clock</name></connection>
<connection>
<GID>3221</GID>
<name>clock</name></connection>
<connection>
<GID>3218</GID>
<name>clock</name></connection>
<connection>
<GID>3215</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3801</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>477.5,-874,479.5,-874</points>
<connection>
<GID>5346</GID>
<name>OUT</name></connection>
<connection>
<GID>5347</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-310.5,478.5,-310.5</points>
<connection>
<GID>3213</GID>
<name>IN_1</name></connection>
<connection>
<GID>3216</GID>
<name>IN_1</name></connection>
<connection>
<GID>3219</GID>
<name>IN_1</name></connection>
<connection>
<GID>3222</GID>
<name>IN_1</name></connection>
<connection>
<GID>3225</GID>
<name>IN_1</name></connection>
<connection>
<GID>3228</GID>
<name>IN_1</name></connection>
<connection>
<GID>3231</GID>
<name>IN_1</name></connection>
<connection>
<GID>3234</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-310.5,242,-307.5</points>
<connection>
<GID>3258</GID>
<name>OUT_0</name></connection>
<intersection>-310.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3802</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>467.5,-877,481.5,-877</points>
<connection>
<GID>5347</GID>
<name>IN_0</name></connection>
<intersection>467.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>467.5,-877,467.5,-864.5</points>
<intersection>-877 1</intersection>
<intersection>-873 4</intersection>
<intersection>-864.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>467.5,-873,471.5,-873</points>
<connection>
<GID>5346</GID>
<name>IN_0</name></connection>
<intersection>467.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>465,-864.5,467.5,-864.5</points>
<connection>
<GID>5348</GID>
<name>OUT_0</name></connection>
<intersection>467.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-318.5,465.5,-318.5</points>
<connection>
<GID>3261</GID>
<name>OUT</name></connection>
<connection>
<GID>3212</GID>
<name>clock</name></connection>
<connection>
<GID>3209</GID>
<name>clock</name></connection>
<connection>
<GID>3206</GID>
<name>clock</name></connection>
<connection>
<GID>3203</GID>
<name>clock</name></connection>
<connection>
<GID>3200</GID>
<name>clock</name></connection>
<connection>
<GID>3197</GID>
<name>clock</name></connection>
<connection>
<GID>3194</GID>
<name>clock</name></connection>
<connection>
<GID>3191</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3803</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>261.5,-858,263.5,-858</points>
<connection>
<GID>5349</GID>
<name>OUT</name></connection>
<connection>
<GID>5350</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-326,478,-326</points>
<connection>
<GID>3189</GID>
<name>IN_1</name></connection>
<connection>
<GID>3192</GID>
<name>IN_1</name></connection>
<connection>
<GID>3195</GID>
<name>IN_1</name></connection>
<connection>
<GID>3198</GID>
<name>IN_1</name></connection>
<connection>
<GID>3201</GID>
<name>IN_1</name></connection>
<connection>
<GID>3204</GID>
<name>IN_1</name></connection>
<connection>
<GID>3207</GID>
<name>IN_1</name></connection>
<connection>
<GID>3210</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-326,242,-323.5</points>
<connection>
<GID>3260</GID>
<name>OUT_0</name></connection>
<intersection>-326 1</intersection></vsegment></shape></wire>
<wire>
<ID>3804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-861.5,265.5,-861</points>
<connection>
<GID>5350</GID>
<name>IN_0</name></connection>
<intersection>-861.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251.5,-861.5,265.5,-861.5</points>
<intersection>251.5 2</intersection>
<intersection>265.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>251.5,-861.5,251.5,-848.5</points>
<intersection>-861.5 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>251.5,-857,255.5,-857</points>
<connection>
<GID>5349</GID>
<name>IN_0</name></connection>
<intersection>251.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>249.5,-848.5,251.5,-848.5</points>
<connection>
<GID>5351</GID>
<name>OUT_0</name></connection>
<intersection>251.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2261</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,-358,300,-358</points>
<connection>
<GID>3144</GID>
<name>OUT</name></connection>
<connection>
<GID>3145</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3805</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>293,-858,295,-858</points>
<connection>
<GID>5352</GID>
<name>OUT</name></connection>
<connection>
<GID>5353</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,-361,302,-361</points>
<connection>
<GID>3145</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288,-361,288,-348.5</points>
<intersection>-361 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,-357,292,-357</points>
<connection>
<GID>3144</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285.5,-348.5,288,-348.5</points>
<connection>
<GID>3146</GID>
<name>OUT_0</name></connection>
<intersection>288 2</intersection></hsegment></shape></wire>
<wire>
<ID>3806</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,-861,297,-861</points>
<connection>
<GID>5353</GID>
<name>IN_0</name></connection>
<intersection>283 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283,-861,283,-848.5</points>
<intersection>-861 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>283,-857,287,-857</points>
<connection>
<GID>5352</GID>
<name>IN_0</name></connection>
<intersection>283 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>280.5,-848.5,283,-848.5</points>
<connection>
<GID>5354</GID>
<name>OUT_0</name></connection>
<intersection>283 2</intersection></hsegment></shape></wire>
<wire>
<ID>2263</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328.5,-358,330.5,-358</points>
<connection>
<GID>3147</GID>
<name>OUT</name></connection>
<connection>
<GID>3148</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3807</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>323.5,-858,325.5,-858</points>
<connection>
<GID>5355</GID>
<name>OUT</name></connection>
<connection>
<GID>5356</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-361.5,332.5,-361</points>
<connection>
<GID>3148</GID>
<name>IN_0</name></connection>
<intersection>-361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-361.5,332.5,-361.5</points>
<intersection>318.5 2</intersection>
<intersection>332.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318.5,-361.5,318.5,-348.5</points>
<intersection>-361.5 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318.5,-357,322.5,-357</points>
<connection>
<GID>3147</GID>
<name>IN_0</name></connection>
<intersection>318.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316.5,-348.5,318.5,-348.5</points>
<connection>
<GID>3149</GID>
<name>OUT_0</name></connection>
<intersection>318.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-861.5,327.5,-861</points>
<connection>
<GID>5356</GID>
<name>IN_0</name></connection>
<intersection>-861.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,-861.5,327.5,-861.5</points>
<intersection>313.5 2</intersection>
<intersection>327.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>313.5,-861.5,313.5,-848.5</points>
<intersection>-861.5 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>313.5,-857,317.5,-857</points>
<connection>
<GID>5355</GID>
<name>IN_0</name></connection>
<intersection>313.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>311.5,-848.5,313.5,-848.5</points>
<connection>
<GID>5357</GID>
<name>OUT_0</name></connection>
<intersection>313.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2265</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360,-358,362,-358</points>
<connection>
<GID>3150</GID>
<name>OUT</name></connection>
<connection>
<GID>3151</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3809</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>355,-858,357,-858</points>
<connection>
<GID>5358</GID>
<name>OUT</name></connection>
<connection>
<GID>5359</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-361,364,-361</points>
<connection>
<GID>3151</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,-361,350,-348.5</points>
<intersection>-361 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350,-357,354,-357</points>
<connection>
<GID>3150</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347.5,-348.5,350,-348.5</points>
<connection>
<GID>3152</GID>
<name>OUT_0</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>3810</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>345,-861,359,-861</points>
<connection>
<GID>5359</GID>
<name>IN_0</name></connection>
<intersection>345 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>345,-861,345,-848.5</points>
<intersection>-861 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>345,-857,349,-857</points>
<connection>
<GID>5358</GID>
<name>IN_0</name></connection>
<intersection>345 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>342.5,-848.5,345,-848.5</points>
<connection>
<GID>5360</GID>
<name>OUT_0</name></connection>
<intersection>345 2</intersection></hsegment></shape></wire>
<wire>
<ID>2267</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389.5,-358,391.5,-358</points>
<connection>
<GID>3153</GID>
<name>OUT</name></connection>
<connection>
<GID>3154</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3811</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>384.5,-858,386.5,-858</points>
<connection>
<GID>5361</GID>
<name>OUT</name></connection>
<connection>
<GID>5362</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,-361.5,393.5,-361</points>
<connection>
<GID>3154</GID>
<name>IN_0</name></connection>
<intersection>-361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-361.5,393.5,-361.5</points>
<intersection>379.5 2</intersection>
<intersection>393.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379.5,-361.5,379.5,-348.5</points>
<intersection>-361.5 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379.5,-357,383.5,-357</points>
<connection>
<GID>3153</GID>
<name>IN_0</name></connection>
<intersection>379.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377.5,-348.5,379.5,-348.5</points>
<connection>
<GID>3155</GID>
<name>OUT_0</name></connection>
<intersection>379.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,-861.5,388.5,-861</points>
<connection>
<GID>5362</GID>
<name>IN_0</name></connection>
<intersection>-861.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-861.5,388.5,-861.5</points>
<intersection>374.5 2</intersection>
<intersection>388.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>374.5,-861.5,374.5,-848.5</points>
<intersection>-861.5 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>374.5,-857,378.5,-857</points>
<connection>
<GID>5361</GID>
<name>IN_0</name></connection>
<intersection>374.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>372.5,-848.5,374.5,-848.5</points>
<connection>
<GID>5363</GID>
<name>OUT_0</name></connection>
<intersection>374.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2269</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421,-358,423,-358</points>
<connection>
<GID>3156</GID>
<name>OUT</name></connection>
<connection>
<GID>3157</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3813</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>416,-858,418,-858</points>
<connection>
<GID>5364</GID>
<name>OUT</name></connection>
<connection>
<GID>5365</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411,-361,425,-361</points>
<connection>
<GID>3157</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411,-361,411,-348.5</points>
<intersection>-361 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411,-357,415,-357</points>
<connection>
<GID>3156</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408.5,-348.5,411,-348.5</points>
<connection>
<GID>3158</GID>
<name>OUT_0</name></connection>
<intersection>411 2</intersection></hsegment></shape></wire>
<wire>
<ID>3814</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406,-861,420,-861</points>
<connection>
<GID>5365</GID>
<name>IN_0</name></connection>
<intersection>406 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>406,-861,406,-848.5</points>
<intersection>-861 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>406,-857,410,-857</points>
<connection>
<GID>5364</GID>
<name>IN_0</name></connection>
<intersection>406 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>403.5,-848.5,406,-848.5</points>
<connection>
<GID>5366</GID>
<name>OUT_0</name></connection>
<intersection>406 2</intersection></hsegment></shape></wire>
<wire>
<ID>2271</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451.5,-358,453.5,-358</points>
<connection>
<GID>3159</GID>
<name>OUT</name></connection>
<connection>
<GID>3160</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3815</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>446.5,-858,448.5,-858</points>
<connection>
<GID>5367</GID>
<name>OUT</name></connection>
<connection>
<GID>5368</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-361.5,455.5,-361</points>
<connection>
<GID>3160</GID>
<name>IN_0</name></connection>
<intersection>-361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,-361.5,455.5,-361.5</points>
<intersection>441.5 2</intersection>
<intersection>455.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441.5,-361.5,441.5,-348.5</points>
<intersection>-361.5 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441.5,-357,445.5,-357</points>
<connection>
<GID>3159</GID>
<name>IN_0</name></connection>
<intersection>441.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439.5,-348.5,441.5,-348.5</points>
<connection>
<GID>3161</GID>
<name>OUT_0</name></connection>
<intersection>441.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3816</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450.5,-861.5,450.5,-861</points>
<connection>
<GID>5368</GID>
<name>IN_0</name></connection>
<intersection>-861.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,-861.5,450.5,-861.5</points>
<intersection>436.5 2</intersection>
<intersection>450.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>436.5,-861.5,436.5,-848.5</points>
<intersection>-861.5 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>436.5,-857,440.5,-857</points>
<connection>
<GID>5367</GID>
<name>IN_0</name></connection>
<intersection>436.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>434.5,-848.5,436.5,-848.5</points>
<connection>
<GID>5369</GID>
<name>OUT_0</name></connection>
<intersection>436.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2273</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483,-358,485,-358</points>
<connection>
<GID>3162</GID>
<name>OUT</name></connection>
<connection>
<GID>3163</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3817</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>478,-858,480,-858</points>
<connection>
<GID>5370</GID>
<name>OUT</name></connection>
<connection>
<GID>5371</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473,-361,487,-361</points>
<connection>
<GID>3163</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473,-361,473,-348.5</points>
<intersection>-361 1</intersection>
<intersection>-357 4</intersection>
<intersection>-348.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473,-357,477,-357</points>
<connection>
<GID>3162</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470.5,-348.5,473,-348.5</points>
<connection>
<GID>3164</GID>
<name>OUT_0</name></connection>
<intersection>473 2</intersection></hsegment></shape></wire>
<wire>
<ID>3818</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>468,-861,482,-861</points>
<connection>
<GID>5371</GID>
<name>IN_0</name></connection>
<intersection>468 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>468,-861,468,-848.5</points>
<intersection>-861 1</intersection>
<intersection>-857 4</intersection>
<intersection>-848.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>468,-857,472,-857</points>
<connection>
<GID>5370</GID>
<name>IN_0</name></connection>
<intersection>468 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>465.5,-848.5,468,-848.5</points>
<connection>
<GID>5372</GID>
<name>OUT_0</name></connection>
<intersection>468 2</intersection></hsegment></shape></wire>
<wire>
<ID>2275</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267,-341,269,-341</points>
<connection>
<GID>3165</GID>
<name>OUT</name></connection>
<connection>
<GID>3166</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3819</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>262,-842.5,264,-842.5</points>
<connection>
<GID>5373</GID>
<name>OUT</name></connection>
<connection>
<GID>5374</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-344.5,271,-344</points>
<connection>
<GID>3166</GID>
<name>IN_0</name></connection>
<intersection>-344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-344.5,271,-344.5</points>
<intersection>257 2</intersection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257,-344.5,257,-331.5</points>
<intersection>-344.5 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,-340,261,-340</points>
<connection>
<GID>3165</GID>
<name>IN_0</name></connection>
<intersection>257 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255,-331.5,257,-331.5</points>
<connection>
<GID>3167</GID>
<name>OUT_0</name></connection>
<intersection>257 2</intersection></hsegment></shape></wire>
<wire>
<ID>3820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-846,266,-845.5</points>
<connection>
<GID>5374</GID>
<name>IN_0</name></connection>
<intersection>-846 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252,-846,266,-846</points>
<intersection>252 2</intersection>
<intersection>266 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,-846,252,-833</points>
<intersection>-846 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>252,-841.5,256,-841.5</points>
<connection>
<GID>5373</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>250,-833,252,-833</points>
<connection>
<GID>5375</GID>
<name>OUT_0</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>2277</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,-341,300.5,-341</points>
<connection>
<GID>3168</GID>
<name>OUT</name></connection>
<connection>
<GID>3169</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3821</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>293.5,-842.5,295.5,-842.5</points>
<connection>
<GID>5376</GID>
<name>OUT</name></connection>
<connection>
<GID>5377</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288.5,-344,302.5,-344</points>
<connection>
<GID>3169</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288.5,-344,288.5,-331.5</points>
<intersection>-344 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,-340,292.5,-340</points>
<connection>
<GID>3168</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,-331.5,288.5,-331.5</points>
<connection>
<GID>3170</GID>
<name>OUT_0</name></connection>
<intersection>288.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3822</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283.5,-845.5,297.5,-845.5</points>
<connection>
<GID>5377</GID>
<name>IN_0</name></connection>
<intersection>283.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283.5,-845.5,283.5,-833</points>
<intersection>-845.5 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>283.5,-841.5,287.5,-841.5</points>
<connection>
<GID>5376</GID>
<name>IN_0</name></connection>
<intersection>283.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>281,-833,283.5,-833</points>
<connection>
<GID>5378</GID>
<name>OUT_0</name></connection>
<intersection>283.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2279</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329,-341,331,-341</points>
<connection>
<GID>3171</GID>
<name>OUT</name></connection>
<connection>
<GID>3172</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3823</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>324,-842.5,326,-842.5</points>
<connection>
<GID>5379</GID>
<name>OUT</name></connection>
<connection>
<GID>5380</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,-344.5,333,-344</points>
<connection>
<GID>3172</GID>
<name>IN_0</name></connection>
<intersection>-344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-344.5,333,-344.5</points>
<intersection>319 2</intersection>
<intersection>333 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319,-344.5,319,-331.5</points>
<intersection>-344.5 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,-340,323,-340</points>
<connection>
<GID>3171</GID>
<name>IN_0</name></connection>
<intersection>319 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317,-331.5,319,-331.5</points>
<connection>
<GID>3173</GID>
<name>OUT_0</name></connection>
<intersection>319 2</intersection></hsegment></shape></wire>
<wire>
<ID>3824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328,-846,328,-845.5</points>
<connection>
<GID>5380</GID>
<name>IN_0</name></connection>
<intersection>-846 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-846,328,-846</points>
<intersection>314 2</intersection>
<intersection>328 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>314,-846,314,-833</points>
<intersection>-846 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>314,-841.5,318,-841.5</points>
<connection>
<GID>5379</GID>
<name>IN_0</name></connection>
<intersection>314 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>312,-833,314,-833</points>
<connection>
<GID>5381</GID>
<name>OUT_0</name></connection>
<intersection>314 2</intersection></hsegment></shape></wire>
<wire>
<ID>2281</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360.5,-341,362.5,-341</points>
<connection>
<GID>3174</GID>
<name>OUT</name></connection>
<connection>
<GID>3175</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3825</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>355.5,-842.5,357.5,-842.5</points>
<connection>
<GID>5382</GID>
<name>OUT</name></connection>
<connection>
<GID>5383</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350.5,-344,364.5,-344</points>
<connection>
<GID>3175</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,-344,350.5,-331.5</points>
<intersection>-344 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350.5,-340,354.5,-340</points>
<connection>
<GID>3174</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348,-331.5,350.5,-331.5</points>
<connection>
<GID>3176</GID>
<name>OUT_0</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>345.5,-845.5,359.5,-845.5</points>
<connection>
<GID>5383</GID>
<name>IN_0</name></connection>
<intersection>345.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>345.5,-845.5,345.5,-833</points>
<intersection>-845.5 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>345.5,-841.5,349.5,-841.5</points>
<connection>
<GID>5382</GID>
<name>IN_0</name></connection>
<intersection>345.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>343,-833,345.5,-833</points>
<connection>
<GID>5384</GID>
<name>OUT_0</name></connection>
<intersection>345.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2283</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390,-341,392,-341</points>
<connection>
<GID>3177</GID>
<name>OUT</name></connection>
<connection>
<GID>3178</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3827</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>385,-842.5,387,-842.5</points>
<connection>
<GID>5385</GID>
<name>OUT</name></connection>
<connection>
<GID>5386</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,-344.5,394,-344</points>
<connection>
<GID>3178</GID>
<name>IN_0</name></connection>
<intersection>-344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-344.5,394,-344.5</points>
<intersection>380 2</intersection>
<intersection>394 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380,-344.5,380,-331.5</points>
<intersection>-344.5 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,-340,384,-340</points>
<connection>
<GID>3177</GID>
<name>IN_0</name></connection>
<intersection>380 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378,-331.5,380,-331.5</points>
<connection>
<GID>3179</GID>
<name>OUT_0</name></connection>
<intersection>380 2</intersection></hsegment></shape></wire>
<wire>
<ID>3828</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389,-846,389,-845.5</points>
<connection>
<GID>5386</GID>
<name>IN_0</name></connection>
<intersection>-846 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375,-846,389,-846</points>
<intersection>375 2</intersection>
<intersection>389 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>375,-846,375,-833</points>
<intersection>-846 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>375,-841.5,379,-841.5</points>
<connection>
<GID>5385</GID>
<name>IN_0</name></connection>
<intersection>375 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>373,-833,375,-833</points>
<connection>
<GID>5387</GID>
<name>OUT_0</name></connection>
<intersection>375 2</intersection></hsegment></shape></wire>
<wire>
<ID>2285</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421.5,-341,423.5,-341</points>
<connection>
<GID>3180</GID>
<name>OUT</name></connection>
<connection>
<GID>3181</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3829</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>416.5,-842.5,418.5,-842.5</points>
<connection>
<GID>5388</GID>
<name>OUT</name></connection>
<connection>
<GID>5389</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411.5,-344,425.5,-344</points>
<connection>
<GID>3181</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411.5,-344,411.5,-331.5</points>
<intersection>-344 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411.5,-340,415.5,-340</points>
<connection>
<GID>3180</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409,-331.5,411.5,-331.5</points>
<connection>
<GID>3182</GID>
<name>OUT_0</name></connection>
<intersection>411.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3830</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406.5,-845.5,420.5,-845.5</points>
<connection>
<GID>5389</GID>
<name>IN_0</name></connection>
<intersection>406.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>406.5,-845.5,406.5,-833</points>
<intersection>-845.5 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>406.5,-841.5,410.5,-841.5</points>
<connection>
<GID>5388</GID>
<name>IN_0</name></connection>
<intersection>406.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>404,-833,406.5,-833</points>
<connection>
<GID>5390</GID>
<name>OUT_0</name></connection>
<intersection>406.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2287</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452,-341,454,-341</points>
<connection>
<GID>3183</GID>
<name>OUT</name></connection>
<connection>
<GID>3184</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3831</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>447,-842.5,449,-842.5</points>
<connection>
<GID>5391</GID>
<name>OUT</name></connection>
<connection>
<GID>5392</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-344.5,456,-344</points>
<connection>
<GID>3184</GID>
<name>IN_0</name></connection>
<intersection>-344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,-344.5,456,-344.5</points>
<intersection>442 2</intersection>
<intersection>456 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442,-344.5,442,-331.5</points>
<intersection>-344.5 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442,-340,446,-340</points>
<connection>
<GID>3183</GID>
<name>IN_0</name></connection>
<intersection>442 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,-331.5,442,-331.5</points>
<connection>
<GID>3185</GID>
<name>OUT_0</name></connection>
<intersection>442 2</intersection></hsegment></shape></wire>
<wire>
<ID>3832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451,-846,451,-845.5</points>
<connection>
<GID>5392</GID>
<name>IN_0</name></connection>
<intersection>-846 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437,-846,451,-846</points>
<intersection>437 2</intersection>
<intersection>451 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>437,-846,437,-833</points>
<intersection>-846 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>437,-841.5,441,-841.5</points>
<connection>
<GID>5391</GID>
<name>IN_0</name></connection>
<intersection>437 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>435,-833,437,-833</points>
<connection>
<GID>5393</GID>
<name>OUT_0</name></connection>
<intersection>437 2</intersection></hsegment></shape></wire>
<wire>
<ID>2289</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483.5,-341,485.5,-341</points>
<connection>
<GID>3186</GID>
<name>OUT</name></connection>
<connection>
<GID>3187</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3833</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>478.5,-842.5,480.5,-842.5</points>
<connection>
<GID>5394</GID>
<name>OUT</name></connection>
<connection>
<GID>5395</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473.5,-344,487.5,-344</points>
<connection>
<GID>3187</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473.5,-344,473.5,-331.5</points>
<intersection>-344 1</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473.5,-340,477.5,-340</points>
<connection>
<GID>3186</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471,-331.5,473.5,-331.5</points>
<connection>
<GID>3188</GID>
<name>OUT_0</name></connection>
<intersection>473.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3834</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>468.5,-845.5,482.5,-845.5</points>
<connection>
<GID>5395</GID>
<name>IN_0</name></connection>
<intersection>468.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>468.5,-845.5,468.5,-833</points>
<intersection>-845.5 1</intersection>
<intersection>-841.5 4</intersection>
<intersection>-833 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>468.5,-841.5,472.5,-841.5</points>
<connection>
<GID>5394</GID>
<name>IN_0</name></connection>
<intersection>468.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>466,-833,468.5,-833</points>
<connection>
<GID>5396</GID>
<name>OUT_0</name></connection>
<intersection>468.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2291</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267.5,-325,269.5,-325</points>
<connection>
<GID>3189</GID>
<name>OUT</name></connection>
<connection>
<GID>3190</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3835</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-867.5,459,-867.5</points>
<connection>
<GID>5423</GID>
<name>OUT</name></connection>
<connection>
<GID>5348</GID>
<name>clock</name></connection>
<connection>
<GID>5345</GID>
<name>clock</name></connection>
<connection>
<GID>5342</GID>
<name>clock</name></connection>
<connection>
<GID>5339</GID>
<name>clock</name></connection>
<connection>
<GID>5336</GID>
<name>clock</name></connection>
<connection>
<GID>5333</GID>
<name>clock</name></connection>
<connection>
<GID>5330</GID>
<name>clock</name></connection>
<connection>
<GID>5327</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-328.5,271.5,-328</points>
<connection>
<GID>3190</GID>
<name>IN_0</name></connection>
<intersection>-328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-328.5,271.5,-328.5</points>
<intersection>257.5 2</intersection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257.5,-328.5,257.5,-315.5</points>
<intersection>-328.5 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257.5,-324,261.5,-324</points>
<connection>
<GID>3189</GID>
<name>IN_0</name></connection>
<intersection>257.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255.5,-315.5,257.5,-315.5</points>
<connection>
<GID>3191</GID>
<name>OUT_0</name></connection>
<intersection>257.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3836</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,-875,471.5,-875</points>
<connection>
<GID>5325</GID>
<name>IN_1</name></connection>
<connection>
<GID>5328</GID>
<name>IN_1</name></connection>
<connection>
<GID>5331</GID>
<name>IN_1</name></connection>
<connection>
<GID>5334</GID>
<name>IN_1</name></connection>
<connection>
<GID>5337</GID>
<name>IN_1</name></connection>
<connection>
<GID>5340</GID>
<name>IN_1</name></connection>
<connection>
<GID>5343</GID>
<name>IN_1</name></connection>
<connection>
<GID>5346</GID>
<name>IN_1</name></connection>
<intersection>236 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>236,-875,236,-872.5</points>
<connection>
<GID>5422</GID>
<name>OUT_0</name></connection>
<intersection>-875 1</intersection></vsegment></shape></wire>
<wire>
<ID>2293</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299,-325,301,-325</points>
<connection>
<GID>3192</GID>
<name>OUT</name></connection>
<connection>
<GID>3193</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3837</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-884.5,458.5,-884.5</points>
<connection>
<GID>5425</GID>
<name>OUT</name></connection>
<connection>
<GID>5324</GID>
<name>clock</name></connection>
<connection>
<GID>5321</GID>
<name>clock</name></connection>
<connection>
<GID>5318</GID>
<name>clock</name></connection>
<connection>
<GID>5315</GID>
<name>clock</name></connection>
<connection>
<GID>5312</GID>
<name>clock</name></connection>
<connection>
<GID>5309</GID>
<name>clock</name></connection>
<connection>
<GID>5306</GID>
<name>clock</name></connection>
<connection>
<GID>5292</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2294</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-328,303,-328</points>
<connection>
<GID>3193</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289,-328,289,-315.5</points>
<intersection>-328 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289,-324,293,-324</points>
<connection>
<GID>3192</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286.5,-315.5,289,-315.5</points>
<connection>
<GID>3194</GID>
<name>OUT_0</name></connection>
<intersection>289 2</intersection></hsegment></shape></wire>
<wire>
<ID>3838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-892,237,-889.5</points>
<intersection>-892 2</intersection>
<intersection>-889.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>237,-892,471,-892</points>
<connection>
<GID>5290</GID>
<name>IN_1</name></connection>
<connection>
<GID>5304</GID>
<name>IN_1</name></connection>
<connection>
<GID>5307</GID>
<name>IN_1</name></connection>
<connection>
<GID>5310</GID>
<name>IN_1</name></connection>
<connection>
<GID>5313</GID>
<name>IN_1</name></connection>
<connection>
<GID>5316</GID>
<name>IN_1</name></connection>
<connection>
<GID>5319</GID>
<name>IN_1</name></connection>
<connection>
<GID>5322</GID>
<name>IN_1</name></connection>
<intersection>237 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>236,-889.5,237,-889.5</points>
<connection>
<GID>5424</GID>
<name>OUT_0</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>2295</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329.5,-325,331.5,-325</points>
<connection>
<GID>3195</GID>
<name>OUT</name></connection>
<connection>
<GID>3196</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-901.5,272.5,-761.5</points>
<connection>
<GID>5302</GID>
<name>N_in0</name></connection>
<connection>
<GID>5294</GID>
<name>N_in1</name></connection>
<intersection>-881.5 1</intersection>
<intersection>-864.5 3</intersection>
<intersection>-848.5 4</intersection>
<intersection>-833 5</intersection>
<intersection>-816.5 6</intersection>
<intersection>-799.5 7</intersection>
<intersection>-783.5 8</intersection>
<intersection>-768 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272.5,-881.5,273.5,-881.5</points>
<connection>
<GID>5306</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>272.5,-768,276,-768</points>
<connection>
<GID>5511</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>272.5,-864.5,274,-864.5</points>
<connection>
<GID>5330</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>272.5,-848.5,274.5,-848.5</points>
<connection>
<GID>5354</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>272.5,-833,275,-833</points>
<connection>
<GID>5378</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>272.5,-816.5,274.5,-816.5</points>
<connection>
<GID>5436</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>272.5,-799.5,275,-799.5</points>
<connection>
<GID>5463</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>272.5,-783.5,275.5,-783.5</points>
<connection>
<GID>5487</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,-328.5,333.5,-328</points>
<connection>
<GID>3196</GID>
<name>IN_0</name></connection>
<intersection>-328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-328.5,333.5,-328.5</points>
<intersection>319.5 2</intersection>
<intersection>333.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319.5,-328.5,319.5,-315.5</points>
<intersection>-328.5 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319.5,-324,323.5,-324</points>
<connection>
<GID>3195</GID>
<name>IN_0</name></connection>
<intersection>319.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317.5,-315.5,319.5,-315.5</points>
<connection>
<GID>3197</GID>
<name>OUT_0</name></connection>
<intersection>319.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,-901.5,304.5,-761.5</points>
<connection>
<GID>5303</GID>
<name>N_in0</name></connection>
<connection>
<GID>5309</GID>
<name>IN_0</name></connection>
<connection>
<GID>5295</GID>
<name>N_in1</name></connection>
<intersection>-864.5 9</intersection>
<intersection>-848.5 10</intersection>
<intersection>-833 7</intersection>
<intersection>-816.5 11</intersection>
<intersection>-799.5 5</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,-768,307,-768</points>
<connection>
<GID>5514</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-783.5,306.5,-783.5</points>
<connection>
<GID>5490</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>304.5,-799.5,306,-799.5</points>
<connection>
<GID>5466</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>304.5,-833,306,-833</points>
<connection>
<GID>5381</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>304.5,-864.5,305,-864.5</points>
<connection>
<GID>5333</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>304.5,-848.5,305.5,-848.5</points>
<connection>
<GID>5357</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>304.5,-816.5,305.5,-816.5</points>
<connection>
<GID>5442</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2297</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361,-325,363,-325</points>
<connection>
<GID>3198</GID>
<name>OUT</name></connection>
<connection>
<GID>3199</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-900.5,335.5,-761.5</points>
<connection>
<GID>5397</GID>
<name>N_in0</name></connection>
<connection>
<GID>5312</GID>
<name>IN_0</name></connection>
<connection>
<GID>5296</GID>
<name>N_in1</name></connection>
<intersection>-864.5 38</intersection>
<intersection>-848.5 21</intersection>
<intersection>-833 7</intersection>
<intersection>-816.5 20</intersection>
<intersection>-799.5 5</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>335.5,-768,338,-768</points>
<connection>
<GID>5517</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>335.5,-783.5,337.5,-783.5</points>
<connection>
<GID>5493</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>335.5,-799.5,337,-799.5</points>
<connection>
<GID>5469</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>335.5,-833,337,-833</points>
<connection>
<GID>5384</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>335.5,-816.5,336.5,-816.5</points>
<connection>
<GID>5445</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>335.5,-848.5,336.5,-848.5</points>
<connection>
<GID>5360</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>335.5,-864.5,336,-864.5</points>
<connection>
<GID>5336</GID>
<name>IN_0</name></connection>
<intersection>335.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351,-328,365,-328</points>
<connection>
<GID>3199</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351,-328,351,-315.5</points>
<intersection>-328 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351,-324,355,-324</points>
<connection>
<GID>3198</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348.5,-315.5,351,-315.5</points>
<connection>
<GID>3200</GID>
<name>OUT_0</name></connection>
<intersection>351 2</intersection></hsegment></shape></wire>
<wire>
<ID>3842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-864.5,366.5,-762</points>
<connection>
<GID>5448</GID>
<name>IN_0</name></connection>
<connection>
<GID>5363</GID>
<name>IN_0</name></connection>
<connection>
<GID>5398</GID>
<name>N_in0</name></connection>
<intersection>-864.5 9</intersection>
<intersection>-833 7</intersection>
<intersection>-799.5 5</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>366.5,-768,368,-768</points>
<connection>
<GID>5520</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366.5,-783.5,367.5,-783.5</points>
<connection>
<GID>5496</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>366.5,-799.5,367,-799.5</points>
<connection>
<GID>5472</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>366.5,-833,367,-833</points>
<connection>
<GID>5387</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>365.5,-864.5,366.5,-864.5</points>
<connection>
<GID>5339</GID>
<name>IN_0</name></connection>
<intersection>365.5 10</intersection>
<intersection>366.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>365.5,-899.5,365.5,-864.5</points>
<connection>
<GID>5315</GID>
<name>IN_0</name></connection>
<connection>
<GID>5297</GID>
<name>N_in1</name></connection>
<intersection>-864.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>2299</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390.5,-325,392.5,-325</points>
<connection>
<GID>3201</GID>
<name>OUT</name></connection>
<connection>
<GID>3202</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3843</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-899,396.5,-761.5</points>
<connection>
<GID>5399</GID>
<name>N_in0</name></connection>
<connection>
<GID>5318</GID>
<name>IN_0</name></connection>
<connection>
<GID>5298</GID>
<name>N_in1</name></connection>
<intersection>-864.5 13</intersection>
<intersection>-848.5 11</intersection>
<intersection>-833 9</intersection>
<intersection>-816.5 7</intersection>
<intersection>-799.5 5</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>396.5,-768,399,-768</points>
<connection>
<GID>5523</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>396.5,-783.5,398.5,-783.5</points>
<connection>
<GID>5499</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>396.5,-799.5,398,-799.5</points>
<connection>
<GID>5475</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>396.5,-816.5,397.5,-816.5</points>
<connection>
<GID>5451</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>396.5,-833,398,-833</points>
<connection>
<GID>5390</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>396.5,-848.5,397.5,-848.5</points>
<connection>
<GID>5366</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>396.5,-864.5,397,-864.5</points>
<connection>
<GID>5342</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,-328.5,394.5,-328</points>
<connection>
<GID>3202</GID>
<name>IN_0</name></connection>
<intersection>-328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,-328.5,394.5,-328.5</points>
<intersection>380.5 2</intersection>
<intersection>394.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380.5,-328.5,380.5,-315.5</points>
<intersection>-328.5 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380.5,-324,384.5,-324</points>
<connection>
<GID>3201</GID>
<name>IN_0</name></connection>
<intersection>380.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378.5,-315.5,380.5,-315.5</points>
<connection>
<GID>3203</GID>
<name>OUT_0</name></connection>
<intersection>380.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-898,427.5,-761.5</points>
<connection>
<GID>5400</GID>
<name>N_in0</name></connection>
<connection>
<GID>5321</GID>
<name>IN_0</name></connection>
<connection>
<GID>5300</GID>
<name>N_in1</name></connection>
<intersection>-864.5 13</intersection>
<intersection>-848.5 11</intersection>
<intersection>-833 9</intersection>
<intersection>-816.5 7</intersection>
<intersection>-799.5 5</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-768,430,-768</points>
<connection>
<GID>5526</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,-783.5,429.5,-783.5</points>
<connection>
<GID>5502</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>427.5,-799.5,429,-799.5</points>
<connection>
<GID>5478</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>427.5,-816.5,428.5,-816.5</points>
<connection>
<GID>5454</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>427.5,-833,429,-833</points>
<connection>
<GID>5393</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>427.5,-848.5,428.5,-848.5</points>
<connection>
<GID>5369</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>427.5,-864.5,428,-864.5</points>
<connection>
<GID>5345</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2301</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422,-325,424,-325</points>
<connection>
<GID>3204</GID>
<name>OUT</name></connection>
<connection>
<GID>3205</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-900,458.5,-762</points>
<connection>
<GID>5401</GID>
<name>N_in0</name></connection>
<connection>
<GID>5324</GID>
<name>IN_0</name></connection>
<connection>
<GID>5299</GID>
<name>N_in1</name></connection>
<intersection>-864.5 13</intersection>
<intersection>-848.5 10</intersection>
<intersection>-833 8</intersection>
<intersection>-816.5 6</intersection>
<intersection>-799.5 4</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>458.5,-768,461,-768</points>
<connection>
<GID>5529</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>458.5,-783.5,460.5,-783.5</points>
<connection>
<GID>5505</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>458.5,-799.5,460,-799.5</points>
<connection>
<GID>5481</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>458.5,-816.5,459.5,-816.5</points>
<connection>
<GID>5457</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>458.5,-833,460,-833</points>
<connection>
<GID>5396</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>458.5,-848.5,459.5,-848.5</points>
<connection>
<GID>5372</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>458.5,-864.5,459,-864.5</points>
<connection>
<GID>5348</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,-328,426,-328</points>
<connection>
<GID>3205</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412,-328,412,-315.5</points>
<intersection>-328 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412,-324,416,-324</points>
<connection>
<GID>3204</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409.5,-315.5,412,-315.5</points>
<connection>
<GID>3206</GID>
<name>OUT_0</name></connection>
<intersection>412 2</intersection></hsegment></shape></wire>
<wire>
<ID>3846</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-888.5,270.5,-754.5</points>
<connection>
<GID>5402</GID>
<name>N_in0</name></connection>
<intersection>-888.5 13</intersection>
<intersection>-871.5 12</intersection>
<intersection>-855.5 11</intersection>
<intersection>-840 10</intersection>
<intersection>-823.5 9</intersection>
<intersection>-806.5 8</intersection>
<intersection>-790.5 7</intersection>
<intersection>-775 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>267,-775,270.5,-775</points>
<connection>
<GID>5507</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>266.5,-790.5,270.5,-790.5</points>
<connection>
<GID>5483</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>266,-806.5,270.5,-806.5</points>
<connection>
<GID>5459</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>265.5,-823.5,270.5,-823.5</points>
<connection>
<GID>5427</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>266,-840,270.5,-840</points>
<connection>
<GID>5374</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>265.5,-855.5,270.5,-855.5</points>
<connection>
<GID>5350</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>265,-871.5,270.5,-871.5</points>
<connection>
<GID>5326</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>264.5,-888.5,270.5,-888.5</points>
<connection>
<GID>5291</GID>
<name>OUT_0</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2303</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452.5,-325,454.5,-325</points>
<connection>
<GID>3207</GID>
<name>OUT</name></connection>
<connection>
<GID>3208</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-888.5,301.5,-754.5</points>
<connection>
<GID>5416</GID>
<name>N_in0</name></connection>
<intersection>-888.5 13</intersection>
<intersection>-871.5 12</intersection>
<intersection>-855.5 11</intersection>
<intersection>-840 10</intersection>
<intersection>-823.5 9</intersection>
<intersection>-806.5 8</intersection>
<intersection>-790.5 7</intersection>
<intersection>-775 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>298.5,-775,301.5,-775</points>
<connection>
<GID>5510</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>298,-790.5,301.5,-790.5</points>
<connection>
<GID>5486</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>297.5,-806.5,301.5,-806.5</points>
<connection>
<GID>5462</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>297,-823.5,301.5,-823.5</points>
<connection>
<GID>5434</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>297.5,-840,301.5,-840</points>
<connection>
<GID>5377</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>297,-855.5,301.5,-855.5</points>
<connection>
<GID>5353</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>296.5,-871.5,301.5,-871.5</points>
<connection>
<GID>5329</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>296,-888.5,301.5,-888.5</points>
<connection>
<GID>5305</GID>
<name>OUT_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-328.5,456.5,-328</points>
<connection>
<GID>3208</GID>
<name>IN_0</name></connection>
<intersection>-328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,-328.5,456.5,-328.5</points>
<intersection>442.5 2</intersection>
<intersection>456.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442.5,-328.5,442.5,-315.5</points>
<intersection>-328.5 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442.5,-324,446.5,-324</points>
<connection>
<GID>3207</GID>
<name>IN_0</name></connection>
<intersection>442.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,-315.5,442.5,-315.5</points>
<connection>
<GID>3209</GID>
<name>OUT_0</name></connection>
<intersection>442.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,-888.5,333.5,-754.5</points>
<connection>
<GID>5415</GID>
<name>N_in0</name></connection>
<intersection>-888.5 13</intersection>
<intersection>-871.5 12</intersection>
<intersection>-855.5 11</intersection>
<intersection>-840 10</intersection>
<intersection>-823.5 9</intersection>
<intersection>-806.5 8</intersection>
<intersection>-790.5 7</intersection>
<intersection>-775 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>329,-775,333.5,-775</points>
<connection>
<GID>5513</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>328.5,-790.5,333.5,-790.5</points>
<connection>
<GID>5489</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>328,-806.5,333.5,-806.5</points>
<connection>
<GID>5465</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>327.5,-823.5,333.5,-823.5</points>
<connection>
<GID>5440</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>328,-840,333.5,-840</points>
<connection>
<GID>5380</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>327.5,-855.5,333.5,-855.5</points>
<connection>
<GID>5356</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>327,-871.5,333.5,-871.5</points>
<connection>
<GID>5332</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>326.5,-888.5,333.5,-888.5</points>
<connection>
<GID>5308</GID>
<name>OUT_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2305</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484,-325,486,-325</points>
<connection>
<GID>3210</GID>
<name>OUT</name></connection>
<connection>
<GID>3211</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364,-888.5,364,-754.5</points>
<connection>
<GID>5414</GID>
<name>N_in0</name></connection>
<intersection>-888.5 18</intersection>
<intersection>-871.5 17</intersection>
<intersection>-855.5 16</intersection>
<intersection>-840 15</intersection>
<intersection>-823.5 14</intersection>
<intersection>-806.5 13</intersection>
<intersection>-790.5 12</intersection>
<intersection>-775 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>360.5,-775,364,-775</points>
<connection>
<GID>5516</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>360,-790.5,364,-790.5</points>
<connection>
<GID>5492</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>359.5,-806.5,364,-806.5</points>
<connection>
<GID>5468</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>359,-823.5,364,-823.5</points>
<connection>
<GID>5444</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>359.5,-840,364,-840</points>
<connection>
<GID>5383</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>359,-855.5,364,-855.5</points>
<connection>
<GID>5359</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>358.5,-871.5,364,-871.5</points>
<connection>
<GID>5335</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>358,-888.5,364,-888.5</points>
<connection>
<GID>5311</GID>
<name>OUT_0</name></connection>
<intersection>364 0</intersection></hsegment></shape></wire>
<wire>
<ID>2306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474,-328,488,-328</points>
<connection>
<GID>3211</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474,-328,474,-315.5</points>
<intersection>-328 1</intersection>
<intersection>-324 4</intersection>
<intersection>-315.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474,-324,478,-324</points>
<connection>
<GID>3210</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471.5,-315.5,474,-315.5</points>
<connection>
<GID>3212</GID>
<name>OUT_0</name></connection>
<intersection>474 2</intersection></hsegment></shape></wire>
<wire>
<ID>3850</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,-888.5,394.5,-754.5</points>
<connection>
<GID>5413</GID>
<name>N_in0</name></connection>
<intersection>-888.5 9</intersection>
<intersection>-871.5 10</intersection>
<intersection>-855.5 11</intersection>
<intersection>-840 12</intersection>
<intersection>-823.5 13</intersection>
<intersection>-806.5 14</intersection>
<intersection>-790.5 15</intersection>
<intersection>-775 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>387.5,-888.5,394.5,-888.5</points>
<connection>
<GID>5314</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>388,-871.5,394.5,-871.5</points>
<connection>
<GID>5338</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>388.5,-855.5,394.5,-855.5</points>
<connection>
<GID>5362</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>389,-840,394.5,-840</points>
<connection>
<GID>5386</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>388.5,-823.5,394.5,-823.5</points>
<connection>
<GID>5447</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>389,-806.5,394.5,-806.5</points>
<connection>
<GID>5471</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>389.5,-790.5,394.5,-790.5</points>
<connection>
<GID>5495</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>390,-775,394.5,-775</points>
<connection>
<GID>5519</GID>
<name>OUT_0</name></connection>
<intersection>394.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2307</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268,-309.5,270,-309.5</points>
<connection>
<GID>3213</GID>
<name>OUT</name></connection>
<connection>
<GID>3214</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3851</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-888.5,425.5,-754.5</points>
<connection>
<GID>5412</GID>
<name>N_in0</name></connection>
<intersection>-888.5 6</intersection>
<intersection>-871.5 7</intersection>
<intersection>-855.5 8</intersection>
<intersection>-840 9</intersection>
<intersection>-823.5 10</intersection>
<intersection>-806.5 11</intersection>
<intersection>-790.5 12</intersection>
<intersection>-775 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>419,-888.5,425.5,-888.5</points>
<connection>
<GID>5317</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>419.5,-871.5,425.5,-871.5</points>
<connection>
<GID>5341</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>420,-855.5,425.5,-855.5</points>
<connection>
<GID>5365</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>420.5,-840,425.5,-840</points>
<connection>
<GID>5389</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>420,-823.5,425.5,-823.5</points>
<connection>
<GID>5450</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>420.5,-806.5,425.5,-806.5</points>
<connection>
<GID>5474</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>421,-790.5,425.5,-790.5</points>
<connection>
<GID>5498</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>421.5,-775,425.5,-775</points>
<connection>
<GID>5522</GID>
<name>OUT_0</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-313,272,-312.5</points>
<connection>
<GID>3214</GID>
<name>IN_0</name></connection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-313,272,-313</points>
<intersection>258 2</intersection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,-313,258,-300</points>
<intersection>-313 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258,-308.5,262,-308.5</points>
<connection>
<GID>3213</GID>
<name>IN_0</name></connection>
<intersection>258 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256,-300,258,-300</points>
<connection>
<GID>3215</GID>
<name>OUT_0</name></connection>
<intersection>258 2</intersection></hsegment></shape></wire>
<wire>
<ID>3852</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-888.5,456.5,-753.5</points>
<connection>
<GID>5411</GID>
<name>N_in0</name></connection>
<intersection>-888.5 6</intersection>
<intersection>-871.5 7</intersection>
<intersection>-855.5 8</intersection>
<intersection>-840 9</intersection>
<intersection>-823.5 10</intersection>
<intersection>-806.5 11</intersection>
<intersection>-790.5 12</intersection>
<intersection>-775 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>449.5,-888.5,456.5,-888.5</points>
<connection>
<GID>5320</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>450,-871.5,456.5,-871.5</points>
<connection>
<GID>5344</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>450.5,-855.5,456.5,-855.5</points>
<connection>
<GID>5368</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>451,-840,456.5,-840</points>
<connection>
<GID>5392</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>450.5,-823.5,456.5,-823.5</points>
<connection>
<GID>5453</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>451,-806.5,456.5,-806.5</points>
<connection>
<GID>5477</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>451.5,-790.5,456.5,-790.5</points>
<connection>
<GID>5501</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>452,-775,456.5,-775</points>
<connection>
<GID>5525</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2309</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299.5,-309.5,301.5,-309.5</points>
<connection>
<GID>3216</GID>
<name>OUT</name></connection>
<connection>
<GID>3217</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3853</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>487,-888.5,487,-753</points>
<connection>
<GID>5410</GID>
<name>N_in0</name></connection>
<intersection>-888.5 3</intersection>
<intersection>-871.5 4</intersection>
<intersection>-855.5 5</intersection>
<intersection>-840 6</intersection>
<intersection>-823.5 7</intersection>
<intersection>-806.5 8</intersection>
<intersection>-790.5 9</intersection>
<intersection>-775 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>481,-888.5,487,-888.5</points>
<connection>
<GID>5323</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>481.5,-871.5,487,-871.5</points>
<connection>
<GID>5347</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>482,-855.5,487,-855.5</points>
<connection>
<GID>5371</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>482.5,-840,487,-840</points>
<connection>
<GID>5395</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>482,-823.5,487,-823.5</points>
<connection>
<GID>5456</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>482.5,-806.5,487,-806.5</points>
<connection>
<GID>5480</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>483,-790.5,487,-790.5</points>
<connection>
<GID>5504</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>483.5,-775,487,-775</points>
<connection>
<GID>5528</GID>
<name>OUT_0</name></connection>
<intersection>487 0</intersection></hsegment></shape></wire>
<wire>
<ID>2310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,-312.5,303.5,-312.5</points>
<connection>
<GID>3217</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289.5,-312.5,289.5,-300</points>
<intersection>-312.5 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289.5,-308.5,293.5,-308.5</points>
<connection>
<GID>3216</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287,-300,289.5,-300</points>
<connection>
<GID>3218</GID>
<name>OUT_0</name></connection>
<intersection>289.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3854</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-822.5,195.5,-773.5</points>
<intersection>-822.5 2</intersection>
<intersection>-773.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,-773.5,234.5,-773.5</points>
<connection>
<GID>5429</GID>
<name>ENABLE_0</name></connection>
<intersection>195.5 0</intersection>
<intersection>220.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-822.5,195.5,-822.5</points>
<connection>
<GID>5417</GID>
<name>OUT_7</name></connection>
<intersection>195.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>220.5,-773.5,220.5,-770</points>
<intersection>-773.5 1</intersection>
<intersection>-770 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220.5,-770,225,-770</points>
<connection>
<GID>5430</GID>
<name>IN_0</name></connection>
<intersection>220.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2311</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330,-309.5,332,-309.5</points>
<connection>
<GID>3219</GID>
<name>OUT</name></connection>
<connection>
<GID>3220</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3855</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-823.5,197.5,-789</points>
<intersection>-823.5 2</intersection>
<intersection>-789 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197.5,-789,234.5,-789</points>
<intersection>197.5 0</intersection>
<intersection>220.5 4</intersection>
<intersection>234.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-823.5,197.5,-823.5</points>
<connection>
<GID>5417</GID>
<name>OUT_6</name></connection>
<intersection>197.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>234.5,-789.5,234.5,-789</points>
<connection>
<GID>5431</GID>
<name>ENABLE_0</name></connection>
<intersection>-789 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>220.5,-789,220.5,-785.5</points>
<intersection>-789 1</intersection>
<intersection>-785.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220.5,-785.5,224.5,-785.5</points>
<connection>
<GID>5433</GID>
<name>IN_0</name></connection>
<intersection>220.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-313,334,-312.5</points>
<connection>
<GID>3220</GID>
<name>IN_0</name></connection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-313,334,-313</points>
<intersection>320 2</intersection>
<intersection>334 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320,-313,320,-300</points>
<intersection>-313 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320,-308.5,324,-308.5</points>
<connection>
<GID>3219</GID>
<name>IN_0</name></connection>
<intersection>320 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318,-300,320,-300</points>
<connection>
<GID>3221</GID>
<name>OUT_0</name></connection>
<intersection>320 2</intersection></hsegment></shape></wire>
<wire>
<ID>3856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-824.5,199.5,-801.5</points>
<intersection>-824.5 2</intersection>
<intersection>-801.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-801.5,224.5,-801.5</points>
<connection>
<GID>5437</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection>
<intersection>220.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-824.5,199.5,-824.5</points>
<connection>
<GID>5417</GID>
<name>OUT_5</name></connection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>220.5,-805.5,220.5,-801.5</points>
<intersection>-805.5 4</intersection>
<intersection>-801.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>220.5,-805.5,234.5,-805.5</points>
<connection>
<GID>5435</GID>
<name>ENABLE_0</name></connection>
<intersection>220.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2313</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361.5,-309.5,363.5,-309.5</points>
<connection>
<GID>3222</GID>
<name>OUT</name></connection>
<connection>
<GID>3223</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-825.5,201.5,-818.5</points>
<intersection>-825.5 2</intersection>
<intersection>-818.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-818.5,224.5,-818.5</points>
<connection>
<GID>5441</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection>
<intersection>220.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-825.5,201.5,-825.5</points>
<connection>
<GID>5417</GID>
<name>OUT_4</name></connection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>220.5,-822.5,220.5,-818.5</points>
<intersection>-822.5 4</intersection>
<intersection>-818.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>220.5,-822.5,234.5,-822.5</points>
<connection>
<GID>5439</GID>
<name>ENABLE_0</name></connection>
<intersection>220.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351.5,-312.5,365.5,-312.5</points>
<connection>
<GID>3223</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351.5,-312.5,351.5,-300</points>
<intersection>-312.5 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351.5,-308.5,355.5,-308.5</points>
<connection>
<GID>3222</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>349,-300,351.5,-300</points>
<connection>
<GID>3224</GID>
<name>OUT_0</name></connection>
<intersection>351.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3858</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-838.5,201.5,-826.5</points>
<intersection>-838.5 1</intersection>
<intersection>-826.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-838.5,233.5,-838.5</points>
<connection>
<GID>5418</GID>
<name>ENABLE_0</name></connection>
<intersection>201.5 0</intersection>
<intersection>220.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-826.5,201.5,-826.5</points>
<connection>
<GID>5417</GID>
<name>OUT_3</name></connection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>220.5,-838.5,220.5,-835</points>
<intersection>-838.5 1</intersection>
<intersection>-835 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220.5,-835,224.5,-835</points>
<connection>
<GID>5419</GID>
<name>IN_0</name></connection>
<intersection>220.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2315</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391,-309.5,393,-309.5</points>
<connection>
<GID>3225</GID>
<name>OUT</name></connection>
<connection>
<GID>3226</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3859</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-854.5,199.5,-827.5</points>
<intersection>-854.5 1</intersection>
<intersection>-827.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-854.5,233.5,-854.5</points>
<connection>
<GID>5420</GID>
<name>ENABLE_0</name></connection>
<intersection>199.5 0</intersection>
<intersection>220.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-827.5,199.5,-827.5</points>
<connection>
<GID>5417</GID>
<name>OUT_2</name></connection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>220.5,-854.5,220.5,-850.5</points>
<intersection>-854.5 1</intersection>
<intersection>-850.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220.5,-850.5,224.5,-850.5</points>
<connection>
<GID>5421</GID>
<name>IN_0</name></connection>
<intersection>220.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395,-313,395,-312.5</points>
<connection>
<GID>3226</GID>
<name>IN_0</name></connection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-313,395,-313</points>
<intersection>381 2</intersection>
<intersection>395 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381,-313,381,-300</points>
<intersection>-313 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381,-308.5,385,-308.5</points>
<connection>
<GID>3225</GID>
<name>IN_0</name></connection>
<intersection>381 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379,-300,381,-300</points>
<connection>
<GID>3227</GID>
<name>OUT_0</name></connection>
<intersection>381 2</intersection></hsegment></shape></wire>
<wire>
<ID>3860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-870,197.5,-828.5</points>
<intersection>-870 1</intersection>
<intersection>-828.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197.5,-870,233.5,-870</points>
<intersection>197.5 0</intersection>
<intersection>220.5 4</intersection>
<intersection>233.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-828.5,197.5,-828.5</points>
<connection>
<GID>5417</GID>
<name>OUT_1</name></connection>
<intersection>197.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>233.5,-870.5,233.5,-870</points>
<connection>
<GID>5422</GID>
<name>ENABLE_0</name></connection>
<intersection>-870 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>220.5,-870,220.5,-866.5</points>
<intersection>-870 1</intersection>
<intersection>-866.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220.5,-866.5,224.5,-866.5</points>
<connection>
<GID>5423</GID>
<name>IN_0</name></connection>
<intersection>220.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2317</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422.5,-309.5,424.5,-309.5</points>
<connection>
<GID>3228</GID>
<name>OUT</name></connection>
<connection>
<GID>3229</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3861</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-887.5,195.5,-829.5</points>
<intersection>-887.5 1</intersection>
<intersection>-829.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,-887.5,233.5,-887.5</points>
<connection>
<GID>5424</GID>
<name>ENABLE_0</name></connection>
<intersection>195.5 0</intersection>
<intersection>220.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-829.5,195.5,-829.5</points>
<connection>
<GID>5417</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>220.5,-887.5,220.5,-883.5</points>
<intersection>-887.5 1</intersection>
<intersection>-883.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220.5,-883.5,224.5,-883.5</points>
<connection>
<GID>5425</GID>
<name>IN_0</name></connection>
<intersection>220.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,-312.5,426.5,-312.5</points>
<connection>
<GID>3229</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412.5,-312.5,412.5,-300</points>
<intersection>-312.5 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412.5,-308.5,416.5,-308.5</points>
<connection>
<GID>3228</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410,-300,412.5,-300</points>
<connection>
<GID>3230</GID>
<name>OUT_0</name></connection>
<intersection>412.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3862</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>261.5,-826,263.5,-826</points>
<connection>
<GID>5426</GID>
<name>OUT</name></connection>
<connection>
<GID>5427</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2319</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453,-309.5,455,-309.5</points>
<connection>
<GID>3231</GID>
<name>OUT</name></connection>
<connection>
<GID>3232</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3863</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-829.5,265.5,-829</points>
<connection>
<GID>5427</GID>
<name>IN_0</name></connection>
<intersection>-829.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251.5,-829.5,265.5,-829.5</points>
<intersection>251.5 2</intersection>
<intersection>265.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>251.5,-829.5,251.5,-816.5</points>
<intersection>-829.5 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>251.5,-825,255.5,-825</points>
<connection>
<GID>5426</GID>
<name>IN_0</name></connection>
<intersection>251.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>249.5,-816.5,251.5,-816.5</points>
<connection>
<GID>5428</GID>
<name>OUT_0</name></connection>
<intersection>251.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-313,457,-312.5</points>
<connection>
<GID>3232</GID>
<name>IN_0</name></connection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443,-313,457,-313</points>
<intersection>443 2</intersection>
<intersection>457 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443,-313,443,-300</points>
<intersection>-313 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443,-308.5,447,-308.5</points>
<connection>
<GID>3231</GID>
<name>IN_0</name></connection>
<intersection>443 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441,-300,443,-300</points>
<connection>
<GID>3233</GID>
<name>OUT_0</name></connection>
<intersection>443 2</intersection></hsegment></shape></wire>
<wire>
<ID>3864</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>293,-826,295,-826</points>
<connection>
<GID>5432</GID>
<name>OUT</name></connection>
<connection>
<GID>5434</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2321</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484.5,-309.5,486.5,-309.5</points>
<connection>
<GID>3234</GID>
<name>OUT</name></connection>
<connection>
<GID>3235</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3865</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283,-829,297,-829</points>
<connection>
<GID>5434</GID>
<name>IN_0</name></connection>
<intersection>283 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283,-829,283,-816.5</points>
<intersection>-829 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>283,-825,287,-825</points>
<connection>
<GID>5432</GID>
<name>IN_0</name></connection>
<intersection>283 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>280.5,-816.5,283,-816.5</points>
<connection>
<GID>5436</GID>
<name>OUT_0</name></connection>
<intersection>283 2</intersection></hsegment></shape></wire>
<wire>
<ID>2322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474.5,-312.5,488.5,-312.5</points>
<connection>
<GID>3235</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474.5,-312.5,474.5,-300</points>
<intersection>-312.5 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-300 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474.5,-308.5,478.5,-308.5</points>
<connection>
<GID>3234</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472,-300,474.5,-300</points>
<connection>
<GID>3236</GID>
<name>OUT_0</name></connection>
<intersection>474.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3866</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>323.5,-826,325.5,-826</points>
<connection>
<GID>5438</GID>
<name>OUT</name></connection>
<connection>
<GID>5440</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-334.5,465,-334.5</points>
<connection>
<GID>3263</GID>
<name>OUT</name></connection>
<connection>
<GID>3188</GID>
<name>clock</name></connection>
<connection>
<GID>3185</GID>
<name>clock</name></connection>
<connection>
<GID>3182</GID>
<name>clock</name></connection>
<connection>
<GID>3179</GID>
<name>clock</name></connection>
<connection>
<GID>3176</GID>
<name>clock</name></connection>
<connection>
<GID>3173</GID>
<name>clock</name></connection>
<connection>
<GID>3170</GID>
<name>clock</name></connection>
<connection>
<GID>3167</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-829.5,327.5,-829</points>
<connection>
<GID>5440</GID>
<name>IN_0</name></connection>
<intersection>-829.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,-829.5,327.5,-829.5</points>
<intersection>313.5 2</intersection>
<intersection>327.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>313.5,-829.5,313.5,-816.5</points>
<intersection>-829.5 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>313.5,-825,317.5,-825</points>
<connection>
<GID>5438</GID>
<name>IN_0</name></connection>
<intersection>313.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>311.5,-816.5,313.5,-816.5</points>
<connection>
<GID>5442</GID>
<name>OUT_0</name></connection>
<intersection>313.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-342,477.5,-342</points>
<connection>
<GID>3165</GID>
<name>IN_1</name></connection>
<connection>
<GID>3168</GID>
<name>IN_1</name></connection>
<connection>
<GID>3171</GID>
<name>IN_1</name></connection>
<connection>
<GID>3174</GID>
<name>IN_1</name></connection>
<connection>
<GID>3177</GID>
<name>IN_1</name></connection>
<connection>
<GID>3180</GID>
<name>IN_1</name></connection>
<connection>
<GID>3183</GID>
<name>IN_1</name></connection>
<connection>
<GID>3186</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-342,242,-339.5</points>
<connection>
<GID>3262</GID>
<name>OUT_0</name></connection>
<intersection>-342 1</intersection></vsegment></shape></wire>
<wire>
<ID>3868</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>355,-826,357,-826</points>
<connection>
<GID>5443</GID>
<name>OUT</name></connection>
<connection>
<GID>5444</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-351.5,464.5,-351.5</points>
<connection>
<GID>3265</GID>
<name>OUT</name></connection>
<connection>
<GID>3164</GID>
<name>clock</name></connection>
<connection>
<GID>3161</GID>
<name>clock</name></connection>
<connection>
<GID>3158</GID>
<name>clock</name></connection>
<connection>
<GID>3155</GID>
<name>clock</name></connection>
<connection>
<GID>3152</GID>
<name>clock</name></connection>
<connection>
<GID>3149</GID>
<name>clock</name></connection>
<connection>
<GID>3146</GID>
<name>clock</name></connection>
<connection>
<GID>3132</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3869</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>345,-829,359,-829</points>
<connection>
<GID>5444</GID>
<name>IN_0</name></connection>
<intersection>345 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>345,-829,345,-816.5</points>
<intersection>-829 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>345,-825,349,-825</points>
<connection>
<GID>5443</GID>
<name>IN_0</name></connection>
<intersection>345 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>342.5,-816.5,345,-816.5</points>
<connection>
<GID>5445</GID>
<name>OUT_0</name></connection>
<intersection>345 2</intersection></hsegment></shape></wire>
<wire>
<ID>2326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-359,243,-356.5</points>
<intersection>-359 2</intersection>
<intersection>-356.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>243,-359,477,-359</points>
<connection>
<GID>3130</GID>
<name>IN_1</name></connection>
<connection>
<GID>3144</GID>
<name>IN_1</name></connection>
<connection>
<GID>3147</GID>
<name>IN_1</name></connection>
<connection>
<GID>3150</GID>
<name>IN_1</name></connection>
<connection>
<GID>3153</GID>
<name>IN_1</name></connection>
<connection>
<GID>3156</GID>
<name>IN_1</name></connection>
<connection>
<GID>3159</GID>
<name>IN_1</name></connection>
<connection>
<GID>3162</GID>
<name>IN_1</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>242,-356.5,243,-356.5</points>
<connection>
<GID>3264</GID>
<name>OUT_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>3870</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>384.5,-826,386.5,-826</points>
<connection>
<GID>5446</GID>
<name>OUT</name></connection>
<connection>
<GID>5447</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-368.5,278.5,-228.5</points>
<connection>
<GID>3142</GID>
<name>N_in0</name></connection>
<connection>
<GID>3134</GID>
<name>N_in1</name></connection>
<intersection>-348.5 1</intersection>
<intersection>-331.5 3</intersection>
<intersection>-315.5 4</intersection>
<intersection>-300 5</intersection>
<intersection>-283.5 6</intersection>
<intersection>-266.5 7</intersection>
<intersection>-250.5 8</intersection>
<intersection>-235 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278.5,-348.5,279.5,-348.5</points>
<connection>
<GID>3146</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278.5,-235,282,-235</points>
<connection>
<GID>3351</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>278.5,-331.5,280,-331.5</points>
<connection>
<GID>3170</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>278.5,-315.5,280.5,-315.5</points>
<connection>
<GID>3194</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>278.5,-300,281,-300</points>
<connection>
<GID>3218</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>278.5,-283.5,280.5,-283.5</points>
<connection>
<GID>3276</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>278.5,-266.5,281,-266.5</points>
<connection>
<GID>3303</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>278.5,-250.5,281.5,-250.5</points>
<connection>
<GID>3327</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3871</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,-829.5,388.5,-829</points>
<connection>
<GID>5447</GID>
<name>IN_0</name></connection>
<intersection>-829.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-829.5,388.5,-829.5</points>
<intersection>374.5 2</intersection>
<intersection>388.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>374.5,-829.5,374.5,-816.5</points>
<intersection>-829.5 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>374.5,-825,378.5,-825</points>
<connection>
<GID>5446</GID>
<name>IN_0</name></connection>
<intersection>374.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>372.5,-816.5,374.5,-816.5</points>
<connection>
<GID>5448</GID>
<name>OUT_0</name></connection>
<intersection>374.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-368.5,310.5,-228.5</points>
<connection>
<GID>3143</GID>
<name>N_in0</name></connection>
<connection>
<GID>3149</GID>
<name>IN_0</name></connection>
<connection>
<GID>3135</GID>
<name>N_in1</name></connection>
<intersection>-331.5 9</intersection>
<intersection>-315.5 10</intersection>
<intersection>-300 7</intersection>
<intersection>-283.5 11</intersection>
<intersection>-266.5 5</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-235,313,-235</points>
<connection>
<GID>3354</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310.5,-250.5,312.5,-250.5</points>
<connection>
<GID>3330</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>310.5,-266.5,312,-266.5</points>
<connection>
<GID>3306</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>310.5,-300,312,-300</points>
<connection>
<GID>3221</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>310.5,-331.5,311,-331.5</points>
<connection>
<GID>3173</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>310.5,-315.5,311.5,-315.5</points>
<connection>
<GID>3197</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>310.5,-283.5,311.5,-283.5</points>
<connection>
<GID>3282</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3872</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>416,-826,418,-826</points>
<connection>
<GID>5449</GID>
<name>OUT</name></connection>
<connection>
<GID>5450</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-367.5,341.5,-228.5</points>
<connection>
<GID>3237</GID>
<name>N_in0</name></connection>
<connection>
<GID>3152</GID>
<name>IN_0</name></connection>
<connection>
<GID>3136</GID>
<name>N_in1</name></connection>
<intersection>-331.5 38</intersection>
<intersection>-315.5 21</intersection>
<intersection>-300 7</intersection>
<intersection>-283.5 20</intersection>
<intersection>-266.5 5</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>341.5,-235,344,-235</points>
<connection>
<GID>3357</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-250.5,343.5,-250.5</points>
<connection>
<GID>3333</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>341.5,-266.5,343,-266.5</points>
<connection>
<GID>3309</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>341.5,-300,343,-300</points>
<connection>
<GID>3224</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>341.5,-283.5,342.5,-283.5</points>
<connection>
<GID>3285</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>341.5,-315.5,342.5,-315.5</points>
<connection>
<GID>3200</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>341.5,-331.5,342,-331.5</points>
<connection>
<GID>3176</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3873</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406,-829,420,-829</points>
<connection>
<GID>5450</GID>
<name>IN_0</name></connection>
<intersection>406 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>406,-829,406,-816.5</points>
<intersection>-829 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>406,-825,410,-825</points>
<connection>
<GID>5449</GID>
<name>IN_0</name></connection>
<intersection>406 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>403.5,-816.5,406,-816.5</points>
<connection>
<GID>5451</GID>
<name>OUT_0</name></connection>
<intersection>406 2</intersection></hsegment></shape></wire>
<wire>
<ID>2330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372.5,-331.5,372.5,-229</points>
<connection>
<GID>3288</GID>
<name>IN_0</name></connection>
<connection>
<GID>3203</GID>
<name>IN_0</name></connection>
<connection>
<GID>3238</GID>
<name>N_in0</name></connection>
<intersection>-331.5 9</intersection>
<intersection>-300 7</intersection>
<intersection>-266.5 5</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372.5,-235,374,-235</points>
<connection>
<GID>3360</GID>
<name>IN_0</name></connection>
<intersection>372.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-250.5,373.5,-250.5</points>
<connection>
<GID>3336</GID>
<name>IN_0</name></connection>
<intersection>372.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>372.5,-266.5,373,-266.5</points>
<connection>
<GID>3312</GID>
<name>IN_0</name></connection>
<intersection>372.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>372.5,-300,373,-300</points>
<connection>
<GID>3227</GID>
<name>IN_0</name></connection>
<intersection>372.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>371.5,-331.5,372.5,-331.5</points>
<connection>
<GID>3179</GID>
<name>IN_0</name></connection>
<intersection>371.5 10</intersection>
<intersection>372.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>371.5,-366.5,371.5,-331.5</points>
<connection>
<GID>3155</GID>
<name>IN_0</name></connection>
<connection>
<GID>3137</GID>
<name>N_in1</name></connection>
<intersection>-331.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>3874</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>446.5,-826,448.5,-826</points>
<connection>
<GID>5452</GID>
<name>OUT</name></connection>
<connection>
<GID>5453</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-366,402.5,-228.5</points>
<connection>
<GID>3239</GID>
<name>N_in0</name></connection>
<connection>
<GID>3158</GID>
<name>IN_0</name></connection>
<connection>
<GID>3138</GID>
<name>N_in1</name></connection>
<intersection>-331.5 13</intersection>
<intersection>-315.5 11</intersection>
<intersection>-300 9</intersection>
<intersection>-283.5 7</intersection>
<intersection>-266.5 5</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,-235,405,-235</points>
<connection>
<GID>3363</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>402.5,-250.5,404.5,-250.5</points>
<connection>
<GID>3339</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>402.5,-266.5,404,-266.5</points>
<connection>
<GID>3315</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>402.5,-283.5,403.5,-283.5</points>
<connection>
<GID>3291</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>402.5,-300,404,-300</points>
<connection>
<GID>3230</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>402.5,-315.5,403.5,-315.5</points>
<connection>
<GID>3206</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>402.5,-331.5,403,-331.5</points>
<connection>
<GID>3182</GID>
<name>IN_0</name></connection>
<intersection>402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450.5,-829.5,450.5,-829</points>
<connection>
<GID>5453</GID>
<name>IN_0</name></connection>
<intersection>-829.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,-829.5,450.5,-829.5</points>
<intersection>436.5 2</intersection>
<intersection>450.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>436.5,-829.5,436.5,-816.5</points>
<intersection>-829.5 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>436.5,-825,440.5,-825</points>
<connection>
<GID>5452</GID>
<name>IN_0</name></connection>
<intersection>436.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>434.5,-816.5,436.5,-816.5</points>
<connection>
<GID>5454</GID>
<name>OUT_0</name></connection>
<intersection>436.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,-365,433.5,-228.5</points>
<connection>
<GID>3240</GID>
<name>N_in0</name></connection>
<connection>
<GID>3161</GID>
<name>IN_0</name></connection>
<connection>
<GID>3140</GID>
<name>N_in1</name></connection>
<intersection>-331.5 13</intersection>
<intersection>-315.5 11</intersection>
<intersection>-300 9</intersection>
<intersection>-283.5 7</intersection>
<intersection>-266.5 5</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433.5,-235,436,-235</points>
<connection>
<GID>3366</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-250.5,435.5,-250.5</points>
<connection>
<GID>3342</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>433.5,-266.5,435,-266.5</points>
<connection>
<GID>3318</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>433.5,-283.5,434.5,-283.5</points>
<connection>
<GID>3294</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>433.5,-300,435,-300</points>
<connection>
<GID>3233</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>433.5,-315.5,434.5,-315.5</points>
<connection>
<GID>3209</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>433.5,-331.5,434,-331.5</points>
<connection>
<GID>3185</GID>
<name>IN_0</name></connection>
<intersection>433.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3876</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>478,-826,480,-826</points>
<connection>
<GID>5455</GID>
<name>OUT</name></connection>
<connection>
<GID>5456</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,-367,464.5,-229</points>
<connection>
<GID>3241</GID>
<name>N_in0</name></connection>
<connection>
<GID>3164</GID>
<name>IN_0</name></connection>
<connection>
<GID>3139</GID>
<name>N_in1</name></connection>
<intersection>-331.5 13</intersection>
<intersection>-315.5 10</intersection>
<intersection>-300 8</intersection>
<intersection>-283.5 6</intersection>
<intersection>-266.5 4</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>464.5,-235,467,-235</points>
<connection>
<GID>3369</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464.5,-250.5,466.5,-250.5</points>
<connection>
<GID>3345</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>464.5,-266.5,466,-266.5</points>
<connection>
<GID>3321</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>464.5,-283.5,465.5,-283.5</points>
<connection>
<GID>3297</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>464.5,-300,466,-300</points>
<connection>
<GID>3236</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>464.5,-315.5,465.5,-315.5</points>
<connection>
<GID>3212</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>464.5,-331.5,465,-331.5</points>
<connection>
<GID>3188</GID>
<name>IN_0</name></connection>
<intersection>464.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3877</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>468,-829,482,-829</points>
<connection>
<GID>5456</GID>
<name>IN_0</name></connection>
<intersection>468 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>468,-829,468,-816.5</points>
<intersection>-829 1</intersection>
<intersection>-825 4</intersection>
<intersection>-816.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>468,-825,472,-825</points>
<connection>
<GID>5455</GID>
<name>IN_0</name></connection>
<intersection>468 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>465.5,-816.5,468,-816.5</points>
<connection>
<GID>5457</GID>
<name>OUT_0</name></connection>
<intersection>468 2</intersection></hsegment></shape></wire>
<wire>
<ID>2334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,-376.5,276.5,-221.5</points>
<connection>
<GID>3243</GID>
<name>N_in1</name></connection>
<connection>
<GID>3242</GID>
<name>N_in0</name></connection>
<intersection>-355.5 13</intersection>
<intersection>-338.5 12</intersection>
<intersection>-322.5 11</intersection>
<intersection>-307 10</intersection>
<intersection>-290.5 9</intersection>
<intersection>-273.5 8</intersection>
<intersection>-257.5 7</intersection>
<intersection>-242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>273,-242,276.5,-242</points>
<connection>
<GID>3347</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>272.5,-257.5,276.5,-257.5</points>
<connection>
<GID>3323</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>272,-273.5,276.5,-273.5</points>
<connection>
<GID>3299</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>271.5,-290.5,276.5,-290.5</points>
<connection>
<GID>3267</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>272,-307,276.5,-307</points>
<connection>
<GID>3214</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>271.5,-322.5,276.5,-322.5</points>
<connection>
<GID>3190</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>271,-338.5,276.5,-338.5</points>
<connection>
<GID>3166</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>270.5,-355.5,276.5,-355.5</points>
<connection>
<GID>3131</GID>
<name>OUT_0</name></connection>
<intersection>276.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3878</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>262,-809,264,-809</points>
<connection>
<GID>5458</GID>
<name>OUT</name></connection>
<connection>
<GID>5459</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-355.5,307.5,-221.5</points>
<connection>
<GID>3256</GID>
<name>N_in0</name></connection>
<intersection>-355.5 13</intersection>
<intersection>-338.5 12</intersection>
<intersection>-322.5 11</intersection>
<intersection>-307 10</intersection>
<intersection>-290.5 9</intersection>
<intersection>-273.5 8</intersection>
<intersection>-257.5 7</intersection>
<intersection>-242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>304.5,-242,307.5,-242</points>
<connection>
<GID>3350</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>304,-257.5,307.5,-257.5</points>
<connection>
<GID>3326</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>303.5,-273.5,307.5,-273.5</points>
<connection>
<GID>3302</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>303,-290.5,307.5,-290.5</points>
<connection>
<GID>3274</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>303.5,-307,307.5,-307</points>
<connection>
<GID>3217</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>303,-322.5,307.5,-322.5</points>
<connection>
<GID>3193</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>302.5,-338.5,307.5,-338.5</points>
<connection>
<GID>3169</GID>
<name>OUT_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>302,-355.5,307.5,-355.5</points>
<connection>
<GID>3145</GID>
<name>OUT_0</name></connection>
<intersection>303.5 22</intersection>
<intersection>307.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>303.5,-373,303.5,-355.5</points>
<connection>
<GID>5779</GID>
<name>N_in1</name></connection>
<intersection>-355.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-812.5,266,-812</points>
<connection>
<GID>5459</GID>
<name>IN_0</name></connection>
<intersection>-812.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252,-812.5,266,-812.5</points>
<intersection>252 2</intersection>
<intersection>266 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,-812.5,252,-799.5</points>
<intersection>-812.5 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>252,-808,256,-808</points>
<connection>
<GID>5458</GID>
<name>IN_0</name></connection>
<intersection>252 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>250,-799.5,252,-799.5</points>
<connection>
<GID>5460</GID>
<name>OUT_0</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>2336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,-375.5,339.5,-221.5</points>
<connection>
<GID>3255</GID>
<name>N_in0</name></connection>
<connection>
<GID>3244</GID>
<name>N_in1</name></connection>
<intersection>-355.5 13</intersection>
<intersection>-338.5 12</intersection>
<intersection>-322.5 11</intersection>
<intersection>-307 10</intersection>
<intersection>-290.5 9</intersection>
<intersection>-273.5 8</intersection>
<intersection>-257.5 7</intersection>
<intersection>-242 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>335,-242,339.5,-242</points>
<connection>
<GID>3353</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>334.5,-257.5,339.5,-257.5</points>
<connection>
<GID>3329</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>334,-273.5,339.5,-273.5</points>
<connection>
<GID>3305</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>333.5,-290.5,339.5,-290.5</points>
<connection>
<GID>3280</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>334,-307,339.5,-307</points>
<connection>
<GID>3220</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>333.5,-322.5,339.5,-322.5</points>
<connection>
<GID>3196</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>333,-338.5,339.5,-338.5</points>
<connection>
<GID>3172</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>332.5,-355.5,339.5,-355.5</points>
<connection>
<GID>3148</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3880</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>293.5,-809,295.5,-809</points>
<connection>
<GID>5461</GID>
<name>OUT</name></connection>
<connection>
<GID>5462</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,-375,370,-221.5</points>
<connection>
<GID>3254</GID>
<name>N_in0</name></connection>
<connection>
<GID>3245</GID>
<name>N_in1</name></connection>
<intersection>-355.5 18</intersection>
<intersection>-338.5 17</intersection>
<intersection>-322.5 16</intersection>
<intersection>-307 15</intersection>
<intersection>-290.5 14</intersection>
<intersection>-273.5 13</intersection>
<intersection>-257.5 12</intersection>
<intersection>-242 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>366.5,-242,370,-242</points>
<connection>
<GID>3356</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>366,-257.5,370,-257.5</points>
<connection>
<GID>3332</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>365.5,-273.5,370,-273.5</points>
<connection>
<GID>3308</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>365,-290.5,370,-290.5</points>
<connection>
<GID>3284</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>365.5,-307,370,-307</points>
<connection>
<GID>3223</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>365,-322.5,370,-322.5</points>
<connection>
<GID>3199</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>364.5,-338.5,370,-338.5</points>
<connection>
<GID>3175</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>364,-355.5,370,-355.5</points>
<connection>
<GID>3151</GID>
<name>OUT_0</name></connection>
<intersection>370 0</intersection></hsegment></shape></wire>
<wire>
<ID>3881</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>283.5,-812,297.5,-812</points>
<connection>
<GID>5462</GID>
<name>IN_0</name></connection>
<intersection>283.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283.5,-812,283.5,-799.5</points>
<intersection>-812 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>283.5,-808,287.5,-808</points>
<connection>
<GID>5461</GID>
<name>IN_0</name></connection>
<intersection>283.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>281,-799.5,283.5,-799.5</points>
<connection>
<GID>5463</GID>
<name>OUT_0</name></connection>
<intersection>283.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,-375,400.5,-221.5</points>
<connection>
<GID>3253</GID>
<name>N_in0</name></connection>
<connection>
<GID>3246</GID>
<name>N_in1</name></connection>
<intersection>-355.5 9</intersection>
<intersection>-338.5 10</intersection>
<intersection>-322.5 11</intersection>
<intersection>-307 12</intersection>
<intersection>-290.5 13</intersection>
<intersection>-273.5 14</intersection>
<intersection>-257.5 15</intersection>
<intersection>-242 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>393.5,-355.5,400.5,-355.5</points>
<connection>
<GID>3154</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>394,-338.5,400.5,-338.5</points>
<connection>
<GID>3178</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>394.5,-322.5,400.5,-322.5</points>
<connection>
<GID>3202</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>395,-307,400.5,-307</points>
<connection>
<GID>3226</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>394.5,-290.5,400.5,-290.5</points>
<connection>
<GID>3287</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>395,-273.5,400.5,-273.5</points>
<connection>
<GID>3311</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>395.5,-257.5,400.5,-257.5</points>
<connection>
<GID>3335</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>396,-242,400.5,-242</points>
<connection>
<GID>3359</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3882</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>324,-809,326,-809</points>
<connection>
<GID>5464</GID>
<name>OUT</name></connection>
<connection>
<GID>5465</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,-375,431.5,-221.5</points>
<connection>
<GID>3252</GID>
<name>N_in0</name></connection>
<connection>
<GID>3247</GID>
<name>N_in1</name></connection>
<intersection>-355.5 6</intersection>
<intersection>-338.5 7</intersection>
<intersection>-322.5 8</intersection>
<intersection>-307 9</intersection>
<intersection>-290.5 10</intersection>
<intersection>-273.5 11</intersection>
<intersection>-257.5 12</intersection>
<intersection>-242 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>425,-355.5,431.5,-355.5</points>
<connection>
<GID>3157</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>425.5,-338.5,431.5,-338.5</points>
<connection>
<GID>3181</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>426,-322.5,431.5,-322.5</points>
<connection>
<GID>3205</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>426.5,-307,431.5,-307</points>
<connection>
<GID>3229</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>426,-290.5,431.5,-290.5</points>
<connection>
<GID>3290</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>426.5,-273.5,431.5,-273.5</points>
<connection>
<GID>3314</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>427,-257.5,431.5,-257.5</points>
<connection>
<GID>3338</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>427.5,-242,431.5,-242</points>
<connection>
<GID>3362</GID>
<name>OUT_0</name></connection>
<intersection>431.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3883</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328,-812.5,328,-812</points>
<connection>
<GID>5465</GID>
<name>IN_0</name></connection>
<intersection>-812.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-812.5,328,-812.5</points>
<intersection>314 2</intersection>
<intersection>328 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>314,-812.5,314,-799.5</points>
<intersection>-812.5 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>314,-808,318,-808</points>
<connection>
<GID>5464</GID>
<name>IN_0</name></connection>
<intersection>314 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>312,-799.5,314,-799.5</points>
<connection>
<GID>5466</GID>
<name>OUT_0</name></connection>
<intersection>314 2</intersection></hsegment></shape></wire>
<wire>
<ID>2340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,-375.5,462.5,-220.5</points>
<connection>
<GID>3251</GID>
<name>N_in0</name></connection>
<connection>
<GID>3248</GID>
<name>N_in1</name></connection>
<intersection>-355.5 6</intersection>
<intersection>-338.5 7</intersection>
<intersection>-322.5 8</intersection>
<intersection>-307 9</intersection>
<intersection>-290.5 10</intersection>
<intersection>-273.5 11</intersection>
<intersection>-257.5 12</intersection>
<intersection>-242 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>455.5,-355.5,462.5,-355.5</points>
<connection>
<GID>3160</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>456,-338.5,462.5,-338.5</points>
<connection>
<GID>3184</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>456.5,-322.5,462.5,-322.5</points>
<connection>
<GID>3208</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>457,-307,462.5,-307</points>
<connection>
<GID>3232</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>456.5,-290.5,462.5,-290.5</points>
<connection>
<GID>3293</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>457,-273.5,462.5,-273.5</points>
<connection>
<GID>3317</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>457.5,-257.5,462.5,-257.5</points>
<connection>
<GID>3341</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>458,-242,462.5,-242</points>
<connection>
<GID>3365</GID>
<name>OUT_0</name></connection>
<intersection>462.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3884</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>355.5,-809,357.5,-809</points>
<connection>
<GID>5467</GID>
<name>OUT</name></connection>
<connection>
<GID>5468</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493,-375,493,-220</points>
<connection>
<GID>3250</GID>
<name>N_in0</name></connection>
<connection>
<GID>3249</GID>
<name>N_in1</name></connection>
<intersection>-355.5 3</intersection>
<intersection>-338.5 4</intersection>
<intersection>-322.5 5</intersection>
<intersection>-307 6</intersection>
<intersection>-290.5 7</intersection>
<intersection>-273.5 8</intersection>
<intersection>-257.5 9</intersection>
<intersection>-242 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>487,-355.5,493,-355.5</points>
<connection>
<GID>3163</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>487.5,-338.5,493,-338.5</points>
<connection>
<GID>3187</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>488,-322.5,493,-322.5</points>
<connection>
<GID>3211</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>488.5,-307,493,-307</points>
<connection>
<GID>3235</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>488,-290.5,493,-290.5</points>
<connection>
<GID>3296</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>488.5,-273.5,493,-273.5</points>
<connection>
<GID>3320</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>489,-257.5,493,-257.5</points>
<connection>
<GID>3344</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>489.5,-242,493,-242</points>
<connection>
<GID>3368</GID>
<name>OUT_0</name></connection>
<intersection>493 0</intersection></hsegment></shape></wire>
<wire>
<ID>3885</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>345.5,-812,359.5,-812</points>
<connection>
<GID>5468</GID>
<name>IN_0</name></connection>
<intersection>345.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>345.5,-812,345.5,-799.5</points>
<intersection>-812 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>345.5,-808,349.5,-808</points>
<connection>
<GID>5467</GID>
<name>IN_0</name></connection>
<intersection>345.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>343,-799.5,345.5,-799.5</points>
<connection>
<GID>5469</GID>
<name>OUT_0</name></connection>
<intersection>345.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-289.5,201.5,-240.5</points>
<intersection>-289.5 2</intersection>
<intersection>-240.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-240.5,240.5,-240.5</points>
<connection>
<GID>3269</GID>
<name>ENABLE_0</name></connection>
<intersection>201.5 0</intersection>
<intersection>226.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-289.5,201.5,-289.5</points>
<connection>
<GID>3257</GID>
<name>OUT_7</name></connection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226.5,-240.5,226.5,-237</points>
<intersection>-240.5 1</intersection>
<intersection>-237 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-237,231,-237</points>
<connection>
<GID>3270</GID>
<name>IN_0</name></connection>
<intersection>226.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3886</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>385,-809,387,-809</points>
<connection>
<GID>5470</GID>
<name>OUT</name></connection>
<connection>
<GID>5471</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-290.5,203.5,-256</points>
<intersection>-290.5 2</intersection>
<intersection>-256 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-256,240.5,-256</points>
<intersection>203.5 0</intersection>
<intersection>226.5 4</intersection>
<intersection>240.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-290.5,203.5,-290.5</points>
<connection>
<GID>3257</GID>
<name>OUT_6</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240.5,-256.5,240.5,-256</points>
<connection>
<GID>3271</GID>
<name>ENABLE_0</name></connection>
<intersection>-256 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>226.5,-256,226.5,-252.5</points>
<intersection>-256 1</intersection>
<intersection>-252.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-252.5,230.5,-252.5</points>
<connection>
<GID>3273</GID>
<name>IN_0</name></connection>
<intersection>226.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3887</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389,-812.5,389,-812</points>
<connection>
<GID>5471</GID>
<name>IN_0</name></connection>
<intersection>-812.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375,-812.5,389,-812.5</points>
<intersection>375 2</intersection>
<intersection>389 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>375,-812.5,375,-799.5</points>
<intersection>-812.5 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>375,-808,379,-808</points>
<connection>
<GID>5470</GID>
<name>IN_0</name></connection>
<intersection>375 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>373,-799.5,375,-799.5</points>
<connection>
<GID>5472</GID>
<name>OUT_0</name></connection>
<intersection>375 2</intersection></hsegment></shape></wire>
<wire>
<ID>2344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-291.5,205.5,-268.5</points>
<intersection>-291.5 2</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-268.5,230.5,-268.5</points>
<connection>
<GID>3277</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection>
<intersection>226.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-291.5,205.5,-291.5</points>
<connection>
<GID>3257</GID>
<name>OUT_5</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>226.5,-272.5,226.5,-268.5</points>
<intersection>-272.5 4</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-272.5,240.5,-272.5</points>
<connection>
<GID>3275</GID>
<name>ENABLE_0</name></connection>
<intersection>226.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3888</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>416.5,-809,418.5,-809</points>
<connection>
<GID>5473</GID>
<name>OUT</name></connection>
<connection>
<GID>5474</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-292.5,207.5,-285.5</points>
<intersection>-292.5 2</intersection>
<intersection>-285.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-285.5,230.5,-285.5</points>
<connection>
<GID>3281</GID>
<name>IN_0</name></connection>
<intersection>207.5 0</intersection>
<intersection>226.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-292.5,207.5,-292.5</points>
<connection>
<GID>3257</GID>
<name>OUT_4</name></connection>
<intersection>207.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>226.5,-289.5,226.5,-285.5</points>
<intersection>-289.5 4</intersection>
<intersection>-285.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-289.5,240.5,-289.5</points>
<connection>
<GID>3279</GID>
<name>ENABLE_0</name></connection>
<intersection>226.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3889</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406.5,-812,420.5,-812</points>
<connection>
<GID>5474</GID>
<name>IN_0</name></connection>
<intersection>406.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>406.5,-812,406.5,-799.5</points>
<intersection>-812 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>406.5,-808,410.5,-808</points>
<connection>
<GID>5473</GID>
<name>IN_0</name></connection>
<intersection>406.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>404,-799.5,406.5,-799.5</points>
<connection>
<GID>5475</GID>
<name>OUT_0</name></connection>
<intersection>406.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-305.5,207.5,-293.5</points>
<intersection>-305.5 1</intersection>
<intersection>-293.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-305.5,239.5,-305.5</points>
<connection>
<GID>3258</GID>
<name>ENABLE_0</name></connection>
<intersection>207.5 0</intersection>
<intersection>226.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-293.5,207.5,-293.5</points>
<connection>
<GID>3257</GID>
<name>OUT_3</name></connection>
<intersection>207.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226.5,-305.5,226.5,-302</points>
<intersection>-305.5 1</intersection>
<intersection>-302 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-302,230.5,-302</points>
<connection>
<GID>3259</GID>
<name>IN_0</name></connection>
<intersection>226.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3890</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>447,-809,449,-809</points>
<connection>
<GID>5476</GID>
<name>OUT</name></connection>
<connection>
<GID>5477</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-321.5,205.5,-294.5</points>
<intersection>-321.5 1</intersection>
<intersection>-294.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-321.5,239.5,-321.5</points>
<connection>
<GID>3260</GID>
<name>ENABLE_0</name></connection>
<intersection>205.5 0</intersection>
<intersection>226.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-294.5,205.5,-294.5</points>
<connection>
<GID>3257</GID>
<name>OUT_2</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226.5,-321.5,226.5,-317.5</points>
<intersection>-321.5 1</intersection>
<intersection>-317.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-317.5,230.5,-317.5</points>
<connection>
<GID>3261</GID>
<name>IN_0</name></connection>
<intersection>226.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451,-812.5,451,-812</points>
<connection>
<GID>5477</GID>
<name>IN_0</name></connection>
<intersection>-812.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437,-812.5,451,-812.5</points>
<intersection>437 2</intersection>
<intersection>451 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>437,-812.5,437,-799.5</points>
<intersection>-812.5 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>437,-808,441,-808</points>
<connection>
<GID>5476</GID>
<name>IN_0</name></connection>
<intersection>437 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>435,-799.5,437,-799.5</points>
<connection>
<GID>5478</GID>
<name>OUT_0</name></connection>
<intersection>437 2</intersection></hsegment></shape></wire>
<wire>
<ID>2348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-337,203.5,-295.5</points>
<intersection>-337 1</intersection>
<intersection>-295.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-337,239.5,-337</points>
<intersection>203.5 0</intersection>
<intersection>226.5 4</intersection>
<intersection>239.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-295.5,203.5,-295.5</points>
<connection>
<GID>3257</GID>
<name>OUT_1</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239.5,-337.5,239.5,-337</points>
<connection>
<GID>3262</GID>
<name>ENABLE_0</name></connection>
<intersection>-337 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>226.5,-337,226.5,-333.5</points>
<intersection>-337 1</intersection>
<intersection>-333.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-333.5,230.5,-333.5</points>
<connection>
<GID>3263</GID>
<name>IN_0</name></connection>
<intersection>226.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3892</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>478.5,-809,480.5,-809</points>
<connection>
<GID>5479</GID>
<name>OUT</name></connection>
<connection>
<GID>5480</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-354.5,201.5,-296.5</points>
<intersection>-354.5 1</intersection>
<intersection>-296.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-354.5,239.5,-354.5</points>
<connection>
<GID>3264</GID>
<name>ENABLE_0</name></connection>
<intersection>201.5 0</intersection>
<intersection>226.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-296.5,201.5,-296.5</points>
<connection>
<GID>3257</GID>
<name>OUT_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226.5,-354.5,226.5,-350.5</points>
<intersection>-354.5 1</intersection>
<intersection>-350.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-350.5,230.5,-350.5</points>
<connection>
<GID>3265</GID>
<name>IN_0</name></connection>
<intersection>226.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3893</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>468.5,-812,482.5,-812</points>
<connection>
<GID>5480</GID>
<name>IN_0</name></connection>
<intersection>468.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>468.5,-812,468.5,-799.5</points>
<intersection>-812 1</intersection>
<intersection>-808 4</intersection>
<intersection>-799.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>468.5,-808,472.5,-808</points>
<connection>
<GID>5479</GID>
<name>IN_0</name></connection>
<intersection>468.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>466,-799.5,468.5,-799.5</points>
<connection>
<GID>5481</GID>
<name>OUT_0</name></connection>
<intersection>468.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2350</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267.5,-293,269.5,-293</points>
<connection>
<GID>3266</GID>
<name>OUT</name></connection>
<connection>
<GID>3267</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3894</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>262.5,-793,264.5,-793</points>
<connection>
<GID>5482</GID>
<name>OUT</name></connection>
<connection>
<GID>5483</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-296.5,271.5,-296</points>
<connection>
<GID>3267</GID>
<name>IN_0</name></connection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-296.5,271.5,-296.5</points>
<intersection>257.5 2</intersection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257.5,-296.5,257.5,-283.5</points>
<intersection>-296.5 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257.5,-292,261.5,-292</points>
<connection>
<GID>3266</GID>
<name>IN_0</name></connection>
<intersection>257.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255.5,-283.5,257.5,-283.5</points>
<connection>
<GID>3268</GID>
<name>OUT_0</name></connection>
<intersection>257.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3895</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-796.5,266.5,-796</points>
<connection>
<GID>5483</GID>
<name>IN_0</name></connection>
<intersection>-796.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252.5,-796.5,266.5,-796.5</points>
<intersection>252.5 2</intersection>
<intersection>266.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252.5,-796.5,252.5,-783.5</points>
<intersection>-796.5 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>252.5,-792,256.5,-792</points>
<connection>
<GID>5482</GID>
<name>IN_0</name></connection>
<intersection>252.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>250.5,-783.5,252.5,-783.5</points>
<connection>
<GID>5484</GID>
<name>OUT_0</name></connection>
<intersection>252.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2352</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299,-293,301,-293</points>
<connection>
<GID>3272</GID>
<name>OUT</name></connection>
<connection>
<GID>3274</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3896</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>294,-793,296,-793</points>
<connection>
<GID>5485</GID>
<name>OUT</name></connection>
<connection>
<GID>5486</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-296,303,-296</points>
<connection>
<GID>3274</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289,-296,289,-283.5</points>
<intersection>-296 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289,-292,293,-292</points>
<connection>
<GID>3272</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286.5,-283.5,289,-283.5</points>
<connection>
<GID>3276</GID>
<name>OUT_0</name></connection>
<intersection>289 2</intersection></hsegment></shape></wire>
<wire>
<ID>3897</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>284,-796,298,-796</points>
<connection>
<GID>5486</GID>
<name>IN_0</name></connection>
<intersection>284 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>284,-796,284,-783.5</points>
<intersection>-796 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>284,-792,288,-792</points>
<connection>
<GID>5485</GID>
<name>IN_0</name></connection>
<intersection>284 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>281.5,-783.5,284,-783.5</points>
<connection>
<GID>5487</GID>
<name>OUT_0</name></connection>
<intersection>284 2</intersection></hsegment></shape></wire>
<wire>
<ID>2354</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329.5,-293,331.5,-293</points>
<connection>
<GID>3278</GID>
<name>OUT</name></connection>
<connection>
<GID>3280</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3898</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>324.5,-793,326.5,-793</points>
<connection>
<GID>5488</GID>
<name>OUT</name></connection>
<connection>
<GID>5489</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,-296.5,333.5,-296</points>
<connection>
<GID>3280</GID>
<name>IN_0</name></connection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-296.5,333.5,-296.5</points>
<intersection>319.5 2</intersection>
<intersection>333.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319.5,-296.5,319.5,-283.5</points>
<intersection>-296.5 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319.5,-292,323.5,-292</points>
<connection>
<GID>3278</GID>
<name>IN_0</name></connection>
<intersection>319.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317.5,-283.5,319.5,-283.5</points>
<connection>
<GID>3282</GID>
<name>OUT_0</name></connection>
<intersection>319.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3899</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-796.5,328.5,-796</points>
<connection>
<GID>5489</GID>
<name>IN_0</name></connection>
<intersection>-796.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314.5,-796.5,328.5,-796.5</points>
<intersection>314.5 2</intersection>
<intersection>328.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>314.5,-796.5,314.5,-783.5</points>
<intersection>-796.5 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>314.5,-792,318.5,-792</points>
<connection>
<GID>5488</GID>
<name>IN_0</name></connection>
<intersection>314.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>312.5,-783.5,314.5,-783.5</points>
<connection>
<GID>5490</GID>
<name>OUT_0</name></connection>
<intersection>314.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2356</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361,-293,363,-293</points>
<connection>
<GID>3283</GID>
<name>OUT</name></connection>
<connection>
<GID>3284</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3900</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>356,-793,358,-793</points>
<connection>
<GID>5491</GID>
<name>OUT</name></connection>
<connection>
<GID>5492</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351,-296,365,-296</points>
<connection>
<GID>3284</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351,-296,351,-283.5</points>
<intersection>-296 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351,-292,355,-292</points>
<connection>
<GID>3283</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348.5,-283.5,351,-283.5</points>
<connection>
<GID>3285</GID>
<name>OUT_0</name></connection>
<intersection>351 2</intersection></hsegment></shape></wire>
<wire>
<ID>3901</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>346,-796,360,-796</points>
<connection>
<GID>5492</GID>
<name>IN_0</name></connection>
<intersection>346 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>346,-796,346,-783.5</points>
<intersection>-796 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>346,-792,350,-792</points>
<connection>
<GID>5491</GID>
<name>IN_0</name></connection>
<intersection>346 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>343.5,-783.5,346,-783.5</points>
<connection>
<GID>5493</GID>
<name>OUT_0</name></connection>
<intersection>346 2</intersection></hsegment></shape></wire>
<wire>
<ID>2358</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390.5,-293,392.5,-293</points>
<connection>
<GID>3286</GID>
<name>OUT</name></connection>
<connection>
<GID>3287</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3902</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>385.5,-793,387.5,-793</points>
<connection>
<GID>5494</GID>
<name>OUT</name></connection>
<connection>
<GID>5495</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,-296.5,394.5,-296</points>
<connection>
<GID>3287</GID>
<name>IN_0</name></connection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,-296.5,394.5,-296.5</points>
<intersection>380.5 2</intersection>
<intersection>394.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380.5,-296.5,380.5,-283.5</points>
<intersection>-296.5 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380.5,-292,384.5,-292</points>
<connection>
<GID>3286</GID>
<name>IN_0</name></connection>
<intersection>380.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378.5,-283.5,380.5,-283.5</points>
<connection>
<GID>3288</GID>
<name>OUT_0</name></connection>
<intersection>380.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3903</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389.5,-796.5,389.5,-796</points>
<connection>
<GID>5495</GID>
<name>IN_0</name></connection>
<intersection>-796.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-796.5,389.5,-796.5</points>
<intersection>375.5 2</intersection>
<intersection>389.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>375.5,-796.5,375.5,-783.5</points>
<intersection>-796.5 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>375.5,-792,379.5,-792</points>
<connection>
<GID>5494</GID>
<name>IN_0</name></connection>
<intersection>375.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>373.5,-783.5,375.5,-783.5</points>
<connection>
<GID>5496</GID>
<name>OUT_0</name></connection>
<intersection>375.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2360</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422,-293,424,-293</points>
<connection>
<GID>3289</GID>
<name>OUT</name></connection>
<connection>
<GID>3290</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3904</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>417,-793,419,-793</points>
<connection>
<GID>5497</GID>
<name>OUT</name></connection>
<connection>
<GID>5498</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2361</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,-296,426,-296</points>
<connection>
<GID>3290</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412,-296,412,-283.5</points>
<intersection>-296 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412,-292,416,-292</points>
<connection>
<GID>3289</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409.5,-283.5,412,-283.5</points>
<connection>
<GID>3291</GID>
<name>OUT_0</name></connection>
<intersection>412 2</intersection></hsegment></shape></wire>
<wire>
<ID>3905</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>407,-796,421,-796</points>
<connection>
<GID>5498</GID>
<name>IN_0</name></connection>
<intersection>407 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>407,-796,407,-783.5</points>
<intersection>-796 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>407,-792,411,-792</points>
<connection>
<GID>5497</GID>
<name>IN_0</name></connection>
<intersection>407 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>404.5,-783.5,407,-783.5</points>
<connection>
<GID>5499</GID>
<name>OUT_0</name></connection>
<intersection>407 2</intersection></hsegment></shape></wire>
<wire>
<ID>2362</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452.5,-293,454.5,-293</points>
<connection>
<GID>3292</GID>
<name>OUT</name></connection>
<connection>
<GID>3293</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3906</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>447.5,-793,449.5,-793</points>
<connection>
<GID>5500</GID>
<name>OUT</name></connection>
<connection>
<GID>5501</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-296.5,456.5,-296</points>
<connection>
<GID>3293</GID>
<name>IN_0</name></connection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,-296.5,456.5,-296.5</points>
<intersection>442.5 2</intersection>
<intersection>456.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442.5,-296.5,442.5,-283.5</points>
<intersection>-296.5 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442.5,-292,446.5,-292</points>
<connection>
<GID>3292</GID>
<name>IN_0</name></connection>
<intersection>442.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,-283.5,442.5,-283.5</points>
<connection>
<GID>3294</GID>
<name>OUT_0</name></connection>
<intersection>442.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3907</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451.5,-796.5,451.5,-796</points>
<connection>
<GID>5501</GID>
<name>IN_0</name></connection>
<intersection>-796.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437.5,-796.5,451.5,-796.5</points>
<intersection>437.5 2</intersection>
<intersection>451.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>437.5,-796.5,437.5,-783.5</points>
<intersection>-796.5 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>437.5,-792,441.5,-792</points>
<connection>
<GID>5500</GID>
<name>IN_0</name></connection>
<intersection>437.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>435.5,-783.5,437.5,-783.5</points>
<connection>
<GID>5502</GID>
<name>OUT_0</name></connection>
<intersection>437.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2364</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484,-293,486,-293</points>
<connection>
<GID>3295</GID>
<name>OUT</name></connection>
<connection>
<GID>3296</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3908</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>479,-793,481,-793</points>
<connection>
<GID>5503</GID>
<name>OUT</name></connection>
<connection>
<GID>5504</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474,-296,488,-296</points>
<connection>
<GID>3296</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474,-296,474,-283.5</points>
<intersection>-296 1</intersection>
<intersection>-292 4</intersection>
<intersection>-283.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474,-292,478,-292</points>
<connection>
<GID>3295</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471.5,-283.5,474,-283.5</points>
<connection>
<GID>3297</GID>
<name>OUT_0</name></connection>
<intersection>474 2</intersection></hsegment></shape></wire>
<wire>
<ID>3909</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>469,-796,483,-796</points>
<connection>
<GID>5504</GID>
<name>IN_0</name></connection>
<intersection>469 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>469,-796,469,-783.5</points>
<intersection>-796 1</intersection>
<intersection>-792 4</intersection>
<intersection>-783.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>469,-792,473,-792</points>
<connection>
<GID>5503</GID>
<name>IN_0</name></connection>
<intersection>469 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>466.5,-783.5,469,-783.5</points>
<connection>
<GID>5505</GID>
<name>OUT_0</name></connection>
<intersection>469 2</intersection></hsegment></shape></wire>
<wire>
<ID>2366</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268,-276,270,-276</points>
<connection>
<GID>3298</GID>
<name>OUT</name></connection>
<connection>
<GID>3299</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3910</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>263,-777.5,265,-777.5</points>
<connection>
<GID>5506</GID>
<name>OUT</name></connection>
<connection>
<GID>5507</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-279.5,272,-279</points>
<connection>
<GID>3299</GID>
<name>IN_0</name></connection>
<intersection>-279.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-279.5,272,-279.5</points>
<intersection>258 2</intersection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,-279.5,258,-266.5</points>
<intersection>-279.5 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258,-275,262,-275</points>
<connection>
<GID>3298</GID>
<name>IN_0</name></connection>
<intersection>258 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256,-266.5,258,-266.5</points>
<connection>
<GID>3300</GID>
<name>OUT_0</name></connection>
<intersection>258 2</intersection></hsegment></shape></wire>
<wire>
<ID>3911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267,-781,267,-780.5</points>
<connection>
<GID>5507</GID>
<name>IN_0</name></connection>
<intersection>-781 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253,-781,267,-781</points>
<intersection>253 2</intersection>
<intersection>267 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>253,-781,253,-768</points>
<intersection>-781 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>253,-776.5,257,-776.5</points>
<connection>
<GID>5506</GID>
<name>IN_0</name></connection>
<intersection>253 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>251,-768,253,-768</points>
<connection>
<GID>5508</GID>
<name>OUT_0</name></connection>
<intersection>253 2</intersection></hsegment></shape></wire>
<wire>
<ID>2368</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299.5,-276,301.5,-276</points>
<connection>
<GID>3301</GID>
<name>OUT</name></connection>
<connection>
<GID>3302</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3912</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>294.5,-777.5,296.5,-777.5</points>
<connection>
<GID>5509</GID>
<name>OUT</name></connection>
<connection>
<GID>5510</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,-279,303.5,-279</points>
<connection>
<GID>3302</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289.5,-279,289.5,-266.5</points>
<intersection>-279 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289.5,-275,293.5,-275</points>
<connection>
<GID>3301</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287,-266.5,289.5,-266.5</points>
<connection>
<GID>3303</GID>
<name>OUT_0</name></connection>
<intersection>289.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3913</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>284.5,-780.5,298.5,-780.5</points>
<connection>
<GID>5510</GID>
<name>IN_0</name></connection>
<intersection>284.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>284.5,-780.5,284.5,-768</points>
<intersection>-780.5 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>284.5,-776.5,288.5,-776.5</points>
<connection>
<GID>5509</GID>
<name>IN_0</name></connection>
<intersection>284.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>282,-768,284.5,-768</points>
<connection>
<GID>5511</GID>
<name>OUT_0</name></connection>
<intersection>284.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2370</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330,-276,332,-276</points>
<connection>
<GID>3304</GID>
<name>OUT</name></connection>
<connection>
<GID>3305</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3914</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>325,-777.5,327,-777.5</points>
<connection>
<GID>5512</GID>
<name>OUT</name></connection>
<connection>
<GID>5513</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-279.5,334,-279</points>
<connection>
<GID>3305</GID>
<name>IN_0</name></connection>
<intersection>-279.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-279.5,334,-279.5</points>
<intersection>320 2</intersection>
<intersection>334 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320,-279.5,320,-266.5</points>
<intersection>-279.5 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320,-275,324,-275</points>
<connection>
<GID>3304</GID>
<name>IN_0</name></connection>
<intersection>320 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318,-266.5,320,-266.5</points>
<connection>
<GID>3306</GID>
<name>OUT_0</name></connection>
<intersection>320 2</intersection></hsegment></shape></wire>
<wire>
<ID>3915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,-781,329,-780.5</points>
<connection>
<GID>5513</GID>
<name>IN_0</name></connection>
<intersection>-781 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-781,329,-781</points>
<intersection>315 2</intersection>
<intersection>329 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>315,-781,315,-768</points>
<intersection>-781 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>315,-776.5,319,-776.5</points>
<connection>
<GID>5512</GID>
<name>IN_0</name></connection>
<intersection>315 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>313,-768,315,-768</points>
<connection>
<GID>5514</GID>
<name>OUT_0</name></connection>
<intersection>315 2</intersection></hsegment></shape></wire>
<wire>
<ID>2372</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361.5,-276,363.5,-276</points>
<connection>
<GID>3307</GID>
<name>OUT</name></connection>
<connection>
<GID>3308</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3916</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>356.5,-777.5,358.5,-777.5</points>
<connection>
<GID>5515</GID>
<name>OUT</name></connection>
<connection>
<GID>5516</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351.5,-279,365.5,-279</points>
<connection>
<GID>3308</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351.5,-279,351.5,-266.5</points>
<intersection>-279 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351.5,-275,355.5,-275</points>
<connection>
<GID>3307</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>349,-266.5,351.5,-266.5</points>
<connection>
<GID>3309</GID>
<name>OUT_0</name></connection>
<intersection>351.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3917</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>346.5,-780.5,360.5,-780.5</points>
<connection>
<GID>5516</GID>
<name>IN_0</name></connection>
<intersection>346.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>346.5,-780.5,346.5,-768</points>
<intersection>-780.5 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>346.5,-776.5,350.5,-776.5</points>
<connection>
<GID>5515</GID>
<name>IN_0</name></connection>
<intersection>346.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>344,-768,346.5,-768</points>
<connection>
<GID>5517</GID>
<name>OUT_0</name></connection>
<intersection>346.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2374</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391,-276,393,-276</points>
<connection>
<GID>3310</GID>
<name>OUT</name></connection>
<connection>
<GID>3311</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3918</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>386,-777.5,388,-777.5</points>
<connection>
<GID>5518</GID>
<name>OUT</name></connection>
<connection>
<GID>5519</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395,-279.5,395,-279</points>
<connection>
<GID>3311</GID>
<name>IN_0</name></connection>
<intersection>-279.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-279.5,395,-279.5</points>
<intersection>381 2</intersection>
<intersection>395 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381,-279.5,381,-266.5</points>
<intersection>-279.5 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381,-275,385,-275</points>
<connection>
<GID>3310</GID>
<name>IN_0</name></connection>
<intersection>381 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379,-266.5,381,-266.5</points>
<connection>
<GID>3312</GID>
<name>OUT_0</name></connection>
<intersection>381 2</intersection></hsegment></shape></wire>
<wire>
<ID>3919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>390,-781,390,-780.5</points>
<connection>
<GID>5519</GID>
<name>IN_0</name></connection>
<intersection>-781 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>376,-781,390,-781</points>
<intersection>376 2</intersection>
<intersection>390 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>376,-781,376,-768</points>
<intersection>-781 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>376,-776.5,380,-776.5</points>
<connection>
<GID>5518</GID>
<name>IN_0</name></connection>
<intersection>376 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>374,-768,376,-768</points>
<connection>
<GID>5520</GID>
<name>OUT_0</name></connection>
<intersection>376 2</intersection></hsegment></shape></wire>
<wire>
<ID>2376</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422.5,-276,424.5,-276</points>
<connection>
<GID>3313</GID>
<name>OUT</name></connection>
<connection>
<GID>3314</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3920</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>417.5,-777.5,419.5,-777.5</points>
<connection>
<GID>5521</GID>
<name>OUT</name></connection>
<connection>
<GID>5522</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,-279,426.5,-279</points>
<connection>
<GID>3314</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412.5,-279,412.5,-266.5</points>
<intersection>-279 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412.5,-275,416.5,-275</points>
<connection>
<GID>3313</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410,-266.5,412.5,-266.5</points>
<connection>
<GID>3315</GID>
<name>OUT_0</name></connection>
<intersection>412.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3921</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>407.5,-780.5,421.5,-780.5</points>
<connection>
<GID>5522</GID>
<name>IN_0</name></connection>
<intersection>407.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>407.5,-780.5,407.5,-768</points>
<intersection>-780.5 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>407.5,-776.5,411.5,-776.5</points>
<connection>
<GID>5521</GID>
<name>IN_0</name></connection>
<intersection>407.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>405,-768,407.5,-768</points>
<connection>
<GID>5523</GID>
<name>OUT_0</name></connection>
<intersection>407.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2378</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453,-276,455,-276</points>
<connection>
<GID>3316</GID>
<name>OUT</name></connection>
<connection>
<GID>3317</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3922</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>448,-777.5,450,-777.5</points>
<connection>
<GID>5524</GID>
<name>OUT</name></connection>
<connection>
<GID>5525</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-279.5,457,-279</points>
<connection>
<GID>3317</GID>
<name>IN_0</name></connection>
<intersection>-279.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443,-279.5,457,-279.5</points>
<intersection>443 2</intersection>
<intersection>457 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443,-279.5,443,-266.5</points>
<intersection>-279.5 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443,-275,447,-275</points>
<connection>
<GID>3316</GID>
<name>IN_0</name></connection>
<intersection>443 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441,-266.5,443,-266.5</points>
<connection>
<GID>3318</GID>
<name>OUT_0</name></connection>
<intersection>443 2</intersection></hsegment></shape></wire>
<wire>
<ID>3923</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-781,452,-780.5</points>
<connection>
<GID>5525</GID>
<name>IN_0</name></connection>
<intersection>-781 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,-781,452,-781</points>
<intersection>438 2</intersection>
<intersection>452 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>438,-781,438,-768</points>
<intersection>-781 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>438,-776.5,442,-776.5</points>
<connection>
<GID>5524</GID>
<name>IN_0</name></connection>
<intersection>438 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>436,-768,438,-768</points>
<connection>
<GID>5526</GID>
<name>OUT_0</name></connection>
<intersection>438 2</intersection></hsegment></shape></wire>
<wire>
<ID>2380</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484.5,-276,486.5,-276</points>
<connection>
<GID>3319</GID>
<name>OUT</name></connection>
<connection>
<GID>3320</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3924</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>479.5,-777.5,481.5,-777.5</points>
<connection>
<GID>5527</GID>
<name>OUT</name></connection>
<connection>
<GID>5528</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2381</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474.5,-279,488.5,-279</points>
<connection>
<GID>3320</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474.5,-279,474.5,-266.5</points>
<intersection>-279 1</intersection>
<intersection>-275 4</intersection>
<intersection>-266.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474.5,-275,478.5,-275</points>
<connection>
<GID>3319</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472,-266.5,474.5,-266.5</points>
<connection>
<GID>3321</GID>
<name>OUT_0</name></connection>
<intersection>474.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3925</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>469.5,-780.5,483.5,-780.5</points>
<connection>
<GID>5528</GID>
<name>IN_0</name></connection>
<intersection>469.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>469.5,-780.5,469.5,-768</points>
<intersection>-780.5 1</intersection>
<intersection>-776.5 4</intersection>
<intersection>-768 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>469.5,-776.5,473.5,-776.5</points>
<connection>
<GID>5527</GID>
<name>IN_0</name></connection>
<intersection>469.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>467,-768,469.5,-768</points>
<connection>
<GID>5529</GID>
<name>OUT_0</name></connection>
<intersection>469.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2382</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268.5,-260,270.5,-260</points>
<connection>
<GID>3322</GID>
<name>OUT</name></connection>
<connection>
<GID>3323</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3926</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-901,241.5,-761.5</points>
<connection>
<GID>5301</GID>
<name>N_in0</name></connection>
<connection>
<GID>5293</GID>
<name>N_in1</name></connection>
<intersection>-881.5 14</intersection>
<intersection>-864.5 12</intersection>
<intersection>-848.5 10</intersection>
<intersection>-833 8</intersection>
<intersection>-816.5 6</intersection>
<intersection>-799.5 4</intersection>
<intersection>-783.5 2</intersection>
<intersection>-768 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241.5,-768,245,-768</points>
<connection>
<GID>5508</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>241.5,-783.5,244.5,-783.5</points>
<connection>
<GID>5484</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>241.5,-799.5,244,-799.5</points>
<connection>
<GID>5460</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>241.5,-816.5,243.5,-816.5</points>
<connection>
<GID>5428</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>241.5,-833,244,-833</points>
<connection>
<GID>5375</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>241.5,-848.5,243.5,-848.5</points>
<connection>
<GID>5351</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>241.5,-864.5,243,-864.5</points>
<connection>
<GID>5327</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>241.5,-881.5,242.5,-881.5</points>
<connection>
<GID>5292</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-263.5,272.5,-263</points>
<connection>
<GID>3323</GID>
<name>IN_0</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,-263.5,272.5,-263.5</points>
<intersection>258.5 2</intersection>
<intersection>272.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258.5,-263.5,258.5,-250.5</points>
<intersection>-263.5 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258.5,-259,262.5,-259</points>
<connection>
<GID>3322</GID>
<name>IN_0</name></connection>
<intersection>258.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256.5,-250.5,258.5,-250.5</points>
<connection>
<GID>3324</GID>
<name>OUT_0</name></connection>
<intersection>258.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3927</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237,-778.5,473.5,-778.5</points>
<connection>
<GID>5506</GID>
<name>IN_1</name></connection>
<connection>
<GID>5509</GID>
<name>IN_1</name></connection>
<connection>
<GID>5512</GID>
<name>IN_1</name></connection>
<connection>
<GID>5515</GID>
<name>IN_1</name></connection>
<connection>
<GID>5518</GID>
<name>IN_1</name></connection>
<connection>
<GID>5521</GID>
<name>IN_1</name></connection>
<connection>
<GID>5524</GID>
<name>IN_1</name></connection>
<connection>
<GID>5527</GID>
<name>IN_1</name></connection>
<intersection>237 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>237,-778.5,237,-775.5</points>
<connection>
<GID>5429</GID>
<name>OUT_0</name></connection>
<intersection>-778.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2384</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>300,-260,302,-260</points>
<connection>
<GID>3325</GID>
<name>OUT</name></connection>
<connection>
<GID>3326</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>231,-771,461,-771</points>
<connection>
<GID>5430</GID>
<name>OUT</name></connection>
<connection>
<GID>5508</GID>
<name>clock</name></connection>
<connection>
<GID>5511</GID>
<name>clock</name></connection>
<connection>
<GID>5514</GID>
<name>clock</name></connection>
<connection>
<GID>5517</GID>
<name>clock</name></connection>
<connection>
<GID>5520</GID>
<name>clock</name></connection>
<connection>
<GID>5523</GID>
<name>clock</name></connection>
<connection>
<GID>5526</GID>
<name>clock</name></connection>
<connection>
<GID>5529</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-263,304,-263</points>
<connection>
<GID>3326</GID>
<name>IN_0</name></connection>
<intersection>290 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>290,-263,290,-250.5</points>
<intersection>-263 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>290,-259,294,-259</points>
<connection>
<GID>3325</GID>
<name>IN_0</name></connection>
<intersection>290 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287.5,-250.5,290,-250.5</points>
<connection>
<GID>3327</GID>
<name>OUT_0</name></connection>
<intersection>290 2</intersection></hsegment></shape></wire>
<wire>
<ID>3929</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266,386.5,268,386.5</points>
<connection>
<GID>5531</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5530</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2386</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330.5,-260,332.5,-260</points>
<connection>
<GID>3328</GID>
<name>OUT</name></connection>
<connection>
<GID>3329</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,383,270,383.5</points>
<connection>
<GID>5531</GID>
<name>IN_0</name></connection>
<intersection>383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,383,270,383</points>
<intersection>256 2</intersection>
<intersection>270 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256,383,256,396</points>
<intersection>383 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256,387.5,260,387.5</points>
<connection>
<GID>5530</GID>
<name>IN_0</name></connection>
<intersection>256 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254,396,256,396</points>
<connection>
<GID>5532</GID>
<name>OUT_0</name></connection>
<intersection>256 2</intersection></hsegment></shape></wire>
<wire>
<ID>2387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,-263.5,334.5,-263</points>
<connection>
<GID>3329</GID>
<name>IN_0</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-263.5,334.5,-263.5</points>
<intersection>320.5 2</intersection>
<intersection>334.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320.5,-263.5,320.5,-250.5</points>
<intersection>-263.5 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320.5,-259,324.5,-259</points>
<connection>
<GID>3328</GID>
<name>IN_0</name></connection>
<intersection>320.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318.5,-250.5,320.5,-250.5</points>
<connection>
<GID>3330</GID>
<name>OUT_0</name></connection>
<intersection>320.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3931</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,483.5,478.5,483.5</points>
<connection>
<GID>5743</GID>
<name>IN_1</name></connection>
<connection>
<GID>5740</GID>
<name>IN_1</name></connection>
<connection>
<GID>5737</GID>
<name>IN_1</name></connection>
<connection>
<GID>5734</GID>
<name>IN_1</name></connection>
<connection>
<GID>5731</GID>
<name>IN_1</name></connection>
<connection>
<GID>5728</GID>
<name>IN_1</name></connection>
<connection>
<GID>5725</GID>
<name>IN_1</name></connection>
<connection>
<GID>5722</GID>
<name>IN_1</name></connection>
<intersection>242.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,483.5,242.5,486</points>
<connection>
<GID>5671</GID>
<name>OUT_0</name></connection>
<intersection>483.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2388</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>362,-260,364,-260</points>
<connection>
<GID>3331</GID>
<name>OUT</name></connection>
<connection>
<GID>3332</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3932</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,491,466,491</points>
<connection>
<GID>5745</GID>
<name>clock</name></connection>
<connection>
<GID>5742</GID>
<name>clock</name></connection>
<connection>
<GID>5739</GID>
<name>clock</name></connection>
<connection>
<GID>5736</GID>
<name>clock</name></connection>
<connection>
<GID>5733</GID>
<name>clock</name></connection>
<connection>
<GID>5730</GID>
<name>clock</name></connection>
<connection>
<GID>5727</GID>
<name>clock</name></connection>
<connection>
<GID>5724</GID>
<name>clock</name></connection>
<connection>
<GID>5673</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>352,-263,366,-263</points>
<connection>
<GID>3332</GID>
<name>IN_0</name></connection>
<intersection>352 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>352,-263,352,-250.5</points>
<intersection>-263 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>352,-259,356,-259</points>
<connection>
<GID>3331</GID>
<name>IN_0</name></connection>
<intersection>352 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>349.5,-250.5,352,-250.5</points>
<connection>
<GID>3333</GID>
<name>OUT_0</name></connection>
<intersection>352 2</intersection></hsegment></shape></wire>
<wire>
<ID>3933</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,467.5,478,467.5</points>
<connection>
<GID>5719</GID>
<name>IN_1</name></connection>
<connection>
<GID>5716</GID>
<name>IN_1</name></connection>
<connection>
<GID>5713</GID>
<name>IN_1</name></connection>
<connection>
<GID>5710</GID>
<name>IN_1</name></connection>
<connection>
<GID>5707</GID>
<name>IN_1</name></connection>
<connection>
<GID>5704</GID>
<name>IN_1</name></connection>
<connection>
<GID>5701</GID>
<name>IN_1</name></connection>
<connection>
<GID>5698</GID>
<name>IN_1</name></connection>
<intersection>242.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,467.5,242.5,470</points>
<connection>
<GID>5675</GID>
<name>OUT_0</name></connection>
<intersection>467.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2390</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391.5,-260,393.5,-260</points>
<connection>
<GID>3334</GID>
<name>OUT</name></connection>
<connection>
<GID>3335</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3934</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,475,465.5,475</points>
<connection>
<GID>5721</GID>
<name>clock</name></connection>
<connection>
<GID>5718</GID>
<name>clock</name></connection>
<connection>
<GID>5715</GID>
<name>clock</name></connection>
<connection>
<GID>5712</GID>
<name>clock</name></connection>
<connection>
<GID>5709</GID>
<name>clock</name></connection>
<connection>
<GID>5706</GID>
<name>clock</name></connection>
<connection>
<GID>5703</GID>
<name>clock</name></connection>
<connection>
<GID>5700</GID>
<name>clock</name></connection>
<connection>
<GID>5677</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395.5,-263.5,395.5,-263</points>
<connection>
<GID>3335</GID>
<name>IN_0</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381.5,-263.5,395.5,-263.5</points>
<intersection>381.5 2</intersection>
<intersection>395.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381.5,-263.5,381.5,-250.5</points>
<intersection>-263.5 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381.5,-259,385.5,-259</points>
<connection>
<GID>3334</GID>
<name>IN_0</name></connection>
<intersection>381.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379.5,-250.5,381.5,-250.5</points>
<connection>
<GID>3336</GID>
<name>OUT_0</name></connection>
<intersection>381.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3935</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,458,465,458</points>
<connection>
<GID>5697</GID>
<name>clock</name></connection>
<connection>
<GID>5694</GID>
<name>clock</name></connection>
<connection>
<GID>5691</GID>
<name>clock</name></connection>
<connection>
<GID>5688</GID>
<name>clock</name></connection>
<connection>
<GID>5685</GID>
<name>clock</name></connection>
<connection>
<GID>5682</GID>
<name>clock</name></connection>
<connection>
<GID>5681</GID>
<name>OUT</name></connection>
<connection>
<GID>5676</GID>
<name>clock</name></connection>
<connection>
<GID>5668</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2392</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>423,-260,425,-260</points>
<connection>
<GID>3337</GID>
<name>OUT</name></connection>
<connection>
<GID>3338</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3936</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,450.5,477.5,450.5</points>
<connection>
<GID>5695</GID>
<name>IN_1</name></connection>
<connection>
<GID>5692</GID>
<name>IN_1</name></connection>
<connection>
<GID>5689</GID>
<name>IN_1</name></connection>
<connection>
<GID>5686</GID>
<name>IN_1</name></connection>
<connection>
<GID>5683</GID>
<name>IN_1</name></connection>
<connection>
<GID>5678</GID>
<name>IN_1</name></connection>
<connection>
<GID>5672</GID>
<name>IN_1</name></connection>
<connection>
<GID>5666</GID>
<name>IN_1</name></connection>
<intersection>242.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,450.5,242.5,453</points>
<connection>
<GID>5679</GID>
<name>OUT_0</name></connection>
<intersection>450.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2393</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413,-263,427,-263</points>
<connection>
<GID>3338</GID>
<name>IN_0</name></connection>
<intersection>413 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>413,-263,413,-250.5</points>
<intersection>-263 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>413,-259,417,-259</points>
<connection>
<GID>3337</GID>
<name>IN_0</name></connection>
<intersection>413 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410.5,-250.5,413,-250.5</points>
<connection>
<GID>3339</GID>
<name>OUT_0</name></connection>
<intersection>413 2</intersection></hsegment></shape></wire>
<wire>
<ID>3937</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,441.5,465.5,441.5</points>
<connection>
<GID>5659</GID>
<name>OUT</name></connection>
<connection>
<GID>5636</GID>
<name>clock</name></connection>
<connection>
<GID>5633</GID>
<name>clock</name></connection>
<connection>
<GID>5630</GID>
<name>clock</name></connection>
<connection>
<GID>5627</GID>
<name>clock</name></connection>
<connection>
<GID>5624</GID>
<name>clock</name></connection>
<connection>
<GID>5621</GID>
<name>clock</name></connection>
<connection>
<GID>5618</GID>
<name>clock</name></connection>
<connection>
<GID>5615</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2394</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453.5,-260,455.5,-260</points>
<connection>
<GID>3340</GID>
<name>OUT</name></connection>
<connection>
<GID>3341</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3938</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241.5,434,478,434</points>
<connection>
<GID>5634</GID>
<name>IN_1</name></connection>
<connection>
<GID>5631</GID>
<name>IN_1</name></connection>
<connection>
<GID>5628</GID>
<name>IN_1</name></connection>
<connection>
<GID>5625</GID>
<name>IN_1</name></connection>
<connection>
<GID>5622</GID>
<name>IN_1</name></connection>
<connection>
<GID>5619</GID>
<name>IN_1</name></connection>
<connection>
<GID>5616</GID>
<name>IN_1</name></connection>
<connection>
<GID>5613</GID>
<name>IN_1</name></connection>
<intersection>241.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241.5,434,241.5,437</points>
<connection>
<GID>5658</GID>
<name>OUT_0</name></connection>
<intersection>434 1</intersection></vsegment></shape></wire>
<wire>
<ID>2395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,-263.5,457.5,-263</points>
<connection>
<GID>3341</GID>
<name>IN_0</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443.5,-263.5,457.5,-263.5</points>
<intersection>443.5 2</intersection>
<intersection>457.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443.5,-263.5,443.5,-250.5</points>
<intersection>-263.5 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443.5,-259,447.5,-259</points>
<connection>
<GID>3340</GID>
<name>IN_0</name></connection>
<intersection>443.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441.5,-250.5,443.5,-250.5</points>
<connection>
<GID>3342</GID>
<name>OUT_0</name></connection>
<intersection>443.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3939</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,426,465,426</points>
<connection>
<GID>5661</GID>
<name>OUT</name></connection>
<connection>
<GID>5612</GID>
<name>clock</name></connection>
<connection>
<GID>5609</GID>
<name>clock</name></connection>
<connection>
<GID>5606</GID>
<name>clock</name></connection>
<connection>
<GID>5603</GID>
<name>clock</name></connection>
<connection>
<GID>5600</GID>
<name>clock</name></connection>
<connection>
<GID>5597</GID>
<name>clock</name></connection>
<connection>
<GID>5594</GID>
<name>clock</name></connection>
<connection>
<GID>5591</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2396</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>485,-260,487,-260</points>
<connection>
<GID>3343</GID>
<name>OUT</name></connection>
<connection>
<GID>3344</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3940</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241.5,418.5,477.5,418.5</points>
<connection>
<GID>5610</GID>
<name>IN_1</name></connection>
<connection>
<GID>5607</GID>
<name>IN_1</name></connection>
<connection>
<GID>5604</GID>
<name>IN_1</name></connection>
<connection>
<GID>5601</GID>
<name>IN_1</name></connection>
<connection>
<GID>5598</GID>
<name>IN_1</name></connection>
<connection>
<GID>5595</GID>
<name>IN_1</name></connection>
<connection>
<GID>5592</GID>
<name>IN_1</name></connection>
<connection>
<GID>5589</GID>
<name>IN_1</name></connection>
<intersection>241.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241.5,418.5,241.5,421</points>
<connection>
<GID>5660</GID>
<name>OUT_0</name></connection>
<intersection>418.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475,-263,489,-263</points>
<connection>
<GID>3344</GID>
<name>IN_0</name></connection>
<intersection>475 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>475,-263,475,-250.5</points>
<intersection>-263 1</intersection>
<intersection>-259 4</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>475,-259,479,-259</points>
<connection>
<GID>3343</GID>
<name>IN_0</name></connection>
<intersection>475 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472.5,-250.5,475,-250.5</points>
<connection>
<GID>3345</GID>
<name>OUT_0</name></connection>
<intersection>475 2</intersection></hsegment></shape></wire>
<wire>
<ID>3941</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297.5,386.5,299.5,386.5</points>
<connection>
<GID>5545</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5544</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2398</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>269,-244.5,271,-244.5</points>
<connection>
<GID>3346</GID>
<name>OUT</name></connection>
<connection>
<GID>3347</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287.5,383.5,301.5,383.5</points>
<connection>
<GID>5545</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287.5,383.5,287.5,396</points>
<intersection>383.5 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,387.5,291.5,387.5</points>
<connection>
<GID>5544</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285,396,287.5,396</points>
<connection>
<GID>5546</GID>
<name>OUT_0</name></connection>
<intersection>287.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-248,273,-247.5</points>
<connection>
<GID>3347</GID>
<name>IN_0</name></connection>
<intersection>-248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259,-248,273,-248</points>
<intersection>259 2</intersection>
<intersection>273 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>259,-248,259,-235</points>
<intersection>-248 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259,-243.5,263,-243.5</points>
<connection>
<GID>3346</GID>
<name>IN_0</name></connection>
<intersection>259 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>257,-235,259,-235</points>
<connection>
<GID>3348</GID>
<name>OUT_0</name></connection>
<intersection>259 2</intersection></hsegment></shape></wire>
<wire>
<ID>3943</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328,386.5,330,386.5</points>
<connection>
<GID>5548</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5547</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2400</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>300.5,-244.5,302.5,-244.5</points>
<connection>
<GID>3349</GID>
<name>OUT</name></connection>
<connection>
<GID>3350</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,383,332,383.5</points>
<connection>
<GID>5548</GID>
<name>IN_0</name></connection>
<intersection>383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,383,332,383</points>
<intersection>318 2</intersection>
<intersection>332 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318,383,318,396</points>
<intersection>383 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318,387.5,322,387.5</points>
<connection>
<GID>5547</GID>
<name>IN_0</name></connection>
<intersection>318 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316,396,318,396</points>
<connection>
<GID>5549</GID>
<name>OUT_0</name></connection>
<intersection>318 2</intersection></hsegment></shape></wire>
<wire>
<ID>2401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,-247.5,304.5,-247.5</points>
<connection>
<GID>3350</GID>
<name>IN_0</name></connection>
<intersection>290.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>290.5,-247.5,290.5,-235</points>
<intersection>-247.5 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>290.5,-243.5,294.5,-243.5</points>
<connection>
<GID>3349</GID>
<name>IN_0</name></connection>
<intersection>290.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>288,-235,290.5,-235</points>
<connection>
<GID>3351</GID>
<name>OUT_0</name></connection>
<intersection>290.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3945</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359.5,386.5,361.5,386.5</points>
<connection>
<GID>5551</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5550</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2402</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>331,-244.5,333,-244.5</points>
<connection>
<GID>3352</GID>
<name>OUT</name></connection>
<connection>
<GID>3353</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3946</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349.5,383.5,363.5,383.5</points>
<connection>
<GID>5551</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349.5,383.5,349.5,396</points>
<intersection>383.5 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349.5,387.5,353.5,387.5</points>
<connection>
<GID>5550</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347,396,349.5,396</points>
<connection>
<GID>5552</GID>
<name>OUT_0</name></connection>
<intersection>349.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-248,335,-247.5</points>
<connection>
<GID>3353</GID>
<name>IN_0</name></connection>
<intersection>-248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,-248,335,-248</points>
<intersection>321 2</intersection>
<intersection>335 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321,-248,321,-235</points>
<intersection>-248 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321,-243.5,325,-243.5</points>
<connection>
<GID>3352</GID>
<name>IN_0</name></connection>
<intersection>321 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>319,-235,321,-235</points>
<connection>
<GID>3354</GID>
<name>OUT_0</name></connection>
<intersection>321 2</intersection></hsegment></shape></wire>
<wire>
<ID>3947</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389,386.5,391,386.5</points>
<connection>
<GID>5554</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5553</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2404</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>362.5,-244.5,364.5,-244.5</points>
<connection>
<GID>3355</GID>
<name>OUT</name></connection>
<connection>
<GID>3356</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,383,393,383.5</points>
<connection>
<GID>5554</GID>
<name>IN_0</name></connection>
<intersection>383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,383,393,383</points>
<intersection>379 2</intersection>
<intersection>393 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379,383,379,396</points>
<intersection>383 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379,387.5,383,387.5</points>
<connection>
<GID>5553</GID>
<name>IN_0</name></connection>
<intersection>379 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377,396,379,396</points>
<connection>
<GID>5555</GID>
<name>OUT_0</name></connection>
<intersection>379 2</intersection></hsegment></shape></wire>
<wire>
<ID>2405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>352.5,-247.5,366.5,-247.5</points>
<connection>
<GID>3356</GID>
<name>IN_0</name></connection>
<intersection>352.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>352.5,-247.5,352.5,-235</points>
<intersection>-247.5 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>352.5,-243.5,356.5,-243.5</points>
<connection>
<GID>3355</GID>
<name>IN_0</name></connection>
<intersection>352.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>350,-235,352.5,-235</points>
<connection>
<GID>3357</GID>
<name>OUT_0</name></connection>
<intersection>352.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3949</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420.5,386.5,422.5,386.5</points>
<connection>
<GID>5557</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5556</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2406</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>392,-244.5,394,-244.5</points>
<connection>
<GID>3358</GID>
<name>OUT</name></connection>
<connection>
<GID>3359</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3950</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410.5,383.5,424.5,383.5</points>
<connection>
<GID>5557</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410.5,383.5,410.5,396</points>
<intersection>383.5 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410.5,387.5,414.5,387.5</points>
<connection>
<GID>5556</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408,396,410.5,396</points>
<connection>
<GID>5558</GID>
<name>OUT_0</name></connection>
<intersection>410.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396,-248,396,-247.5</points>
<connection>
<GID>3359</GID>
<name>IN_0</name></connection>
<intersection>-248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382,-248,396,-248</points>
<intersection>382 2</intersection>
<intersection>396 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>382,-248,382,-235</points>
<intersection>-248 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>382,-243.5,386,-243.5</points>
<connection>
<GID>3358</GID>
<name>IN_0</name></connection>
<intersection>382 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380,-235,382,-235</points>
<connection>
<GID>3360</GID>
<name>OUT_0</name></connection>
<intersection>382 2</intersection></hsegment></shape></wire>
<wire>
<ID>3951</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451,386.5,453,386.5</points>
<connection>
<GID>5560</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5559</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2408</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>423.5,-244.5,425.5,-244.5</points>
<connection>
<GID>3361</GID>
<name>OUT</name></connection>
<connection>
<GID>3362</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,383,455,383.5</points>
<connection>
<GID>5560</GID>
<name>IN_0</name></connection>
<intersection>383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,383,455,383</points>
<intersection>441 2</intersection>
<intersection>455 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441,383,441,396</points>
<intersection>383 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441,387.5,445,387.5</points>
<connection>
<GID>5559</GID>
<name>IN_0</name></connection>
<intersection>441 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439,396,441,396</points>
<connection>
<GID>5561</GID>
<name>OUT_0</name></connection>
<intersection>441 2</intersection></hsegment></shape></wire>
<wire>
<ID>2409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413.5,-247.5,427.5,-247.5</points>
<connection>
<GID>3362</GID>
<name>IN_0</name></connection>
<intersection>413.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>413.5,-247.5,413.5,-235</points>
<intersection>-247.5 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>413.5,-243.5,417.5,-243.5</points>
<connection>
<GID>3361</GID>
<name>IN_0</name></connection>
<intersection>413.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411,-235,413.5,-235</points>
<connection>
<GID>3363</GID>
<name>OUT_0</name></connection>
<intersection>413.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3953</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482.5,386.5,484.5,386.5</points>
<connection>
<GID>5563</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5562</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2410</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>454,-244.5,456,-244.5</points>
<connection>
<GID>3364</GID>
<name>OUT</name></connection>
<connection>
<GID>3365</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472.5,383.5,486.5,383.5</points>
<connection>
<GID>5563</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472.5,383.5,472.5,396</points>
<intersection>383.5 1</intersection>
<intersection>387.5 4</intersection>
<intersection>396 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472.5,387.5,476.5,387.5</points>
<connection>
<GID>5562</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470,396,472.5,396</points>
<connection>
<GID>5564</GID>
<name>OUT_0</name></connection>
<intersection>472.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,-248,458,-247.5</points>
<connection>
<GID>3365</GID>
<name>IN_0</name></connection>
<intersection>-248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444,-248,458,-248</points>
<intersection>444 2</intersection>
<intersection>458 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>444,-248,444,-235</points>
<intersection>-248 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>444,-243.5,448,-243.5</points>
<connection>
<GID>3364</GID>
<name>IN_0</name></connection>
<intersection>444 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>442,-235,444,-235</points>
<connection>
<GID>3366</GID>
<name>OUT_0</name></connection>
<intersection>444 2</intersection></hsegment></shape></wire>
<wire>
<ID>3955</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266.5,403.5,268.5,403.5</points>
<connection>
<GID>5566</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5565</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2412</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>485.5,-244.5,487.5,-244.5</points>
<connection>
<GID>3367</GID>
<name>OUT</name></connection>
<connection>
<GID>3368</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,400,270.5,400.5</points>
<connection>
<GID>5566</GID>
<name>IN_0</name></connection>
<intersection>400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,400,270.5,400</points>
<intersection>256.5 2</intersection>
<intersection>270.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256.5,400,256.5,413</points>
<intersection>400 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256.5,404.5,260.5,404.5</points>
<connection>
<GID>5565</GID>
<name>IN_0</name></connection>
<intersection>256.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254.5,413,256.5,413</points>
<connection>
<GID>5567</GID>
<name>OUT_0</name></connection>
<intersection>256.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475.5,-247.5,489.5,-247.5</points>
<connection>
<GID>3368</GID>
<name>IN_0</name></connection>
<intersection>475.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>475.5,-247.5,475.5,-235</points>
<intersection>-247.5 1</intersection>
<intersection>-243.5 4</intersection>
<intersection>-235 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>475.5,-243.5,479.5,-243.5</points>
<connection>
<GID>3367</GID>
<name>IN_0</name></connection>
<intersection>475.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>473,-235,475.5,-235</points>
<connection>
<GID>3369</GID>
<name>OUT_0</name></connection>
<intersection>475.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3957</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,403.5,300,403.5</points>
<connection>
<GID>5569</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5568</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-368,247.5,-228.5</points>
<connection>
<GID>3141</GID>
<name>N_in0</name></connection>
<connection>
<GID>3133</GID>
<name>N_in1</name></connection>
<intersection>-348.5 14</intersection>
<intersection>-331.5 12</intersection>
<intersection>-315.5 10</intersection>
<intersection>-300 8</intersection>
<intersection>-283.5 6</intersection>
<intersection>-266.5 4</intersection>
<intersection>-250.5 2</intersection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247.5,-235,251,-235</points>
<connection>
<GID>3348</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-250.5,250.5,-250.5</points>
<connection>
<GID>3324</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>247.5,-266.5,250,-266.5</points>
<connection>
<GID>3300</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>247.5,-283.5,249.5,-283.5</points>
<connection>
<GID>3268</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>247.5,-300,250,-300</points>
<connection>
<GID>3215</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>247.5,-315.5,249.5,-315.5</points>
<connection>
<GID>3191</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>247.5,-331.5,249,-331.5</points>
<connection>
<GID>3167</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>247.5,-348.5,248.5,-348.5</points>
<connection>
<GID>3132</GID>
<name>IN_0</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3958</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,400.5,302,400.5</points>
<connection>
<GID>5569</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288,400.5,288,413</points>
<intersection>400.5 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,404.5,292,404.5</points>
<connection>
<GID>5568</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285.5,413,288,413</points>
<connection>
<GID>5570</GID>
<name>OUT_0</name></connection>
<intersection>288 2</intersection></hsegment></shape></wire>
<wire>
<ID>2415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243,-245.5,479.5,-245.5</points>
<connection>
<GID>3346</GID>
<name>IN_1</name></connection>
<connection>
<GID>3349</GID>
<name>IN_1</name></connection>
<connection>
<GID>3352</GID>
<name>IN_1</name></connection>
<connection>
<GID>3355</GID>
<name>IN_1</name></connection>
<connection>
<GID>3358</GID>
<name>IN_1</name></connection>
<connection>
<GID>3361</GID>
<name>IN_1</name></connection>
<connection>
<GID>3364</GID>
<name>IN_1</name></connection>
<connection>
<GID>3367</GID>
<name>IN_1</name></connection>
<intersection>243 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243,-245.5,243,-242.5</points>
<connection>
<GID>3269</GID>
<name>OUT_0</name></connection>
<intersection>-245.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3959</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328.5,403.5,330.5,403.5</points>
<connection>
<GID>5572</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5571</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237,-238,467,-238</points>
<connection>
<GID>3270</GID>
<name>OUT</name></connection>
<connection>
<GID>3348</GID>
<name>clock</name></connection>
<connection>
<GID>3351</GID>
<name>clock</name></connection>
<connection>
<GID>3354</GID>
<name>clock</name></connection>
<connection>
<GID>3357</GID>
<name>clock</name></connection>
<connection>
<GID>3360</GID>
<name>clock</name></connection>
<connection>
<GID>3363</GID>
<name>clock</name></connection>
<connection>
<GID>3366</GID>
<name>clock</name></connection>
<connection>
<GID>3369</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,400,332.5,400.5</points>
<connection>
<GID>5572</GID>
<name>IN_0</name></connection>
<intersection>400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,400,332.5,400</points>
<intersection>318.5 2</intersection>
<intersection>332.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318.5,400,318.5,413</points>
<intersection>400 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318.5,404.5,322.5,404.5</points>
<connection>
<GID>5571</GID>
<name>IN_0</name></connection>
<intersection>318.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316.5,413,318.5,413</points>
<connection>
<GID>5573</GID>
<name>OUT_0</name></connection>
<intersection>318.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2417</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266.5,-531,271.5,-531</points>
<connection>
<GID>3370</GID>
<name>OUT</name></connection>
<connection>
<GID>3371</GID>
<name>ENABLE_0</name></connection>
<intersection>266.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>266.5,-531,266.5,-530</points>
<intersection>-531 6</intersection>
<intersection>-530 12</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>273.5,-534.5,273.5,-534</points>
<connection>
<GID>3371</GID>
<name>IN_0</name></connection>
<intersection>-534.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>259.5,-534.5,273.5,-534.5</points>
<intersection>259.5 10</intersection>
<intersection>273.5 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>259.5,-534.5,259.5,-521.5</points>
<intersection>-534.5 9</intersection>
<intersection>-530 12</intersection>
<intersection>-521.5 14</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>259.5,-530,266.5,-530</points>
<connection>
<GID>3370</GID>
<name>IN_0</name></connection>
<intersection>259.5 10</intersection>
<intersection>266.5 7</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>257.5,-521.5,259.5,-521.5</points>
<connection>
<GID>3372</GID>
<name>OUT_0</name></connection>
<intersection>259.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>3961</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360,403.5,362,403.5</points>
<connection>
<GID>5575</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5574</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3962</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,400.5,364,400.5</points>
<connection>
<GID>5575</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,400.5,350,413</points>
<intersection>400.5 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350,404.5,354,404.5</points>
<connection>
<GID>5574</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347.5,413,350,413</points>
<connection>
<GID>5576</GID>
<name>OUT_0</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>2419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,-434,482,-434</points>
<connection>
<GID>3562</GID>
<name>IN_1</name></connection>
<connection>
<GID>3565</GID>
<name>IN_1</name></connection>
<connection>
<GID>3568</GID>
<name>IN_1</name></connection>
<connection>
<GID>3571</GID>
<name>IN_1</name></connection>
<connection>
<GID>3574</GID>
<name>IN_1</name></connection>
<connection>
<GID>3577</GID>
<name>IN_1</name></connection>
<connection>
<GID>3580</GID>
<name>IN_1</name></connection>
<connection>
<GID>3583</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,-434,246,-431.5</points>
<connection>
<GID>3511</GID>
<name>OUT_0</name></connection>
<intersection>-434 1</intersection></vsegment></shape></wire>
<wire>
<ID>3963</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389.5,403.5,391.5,403.5</points>
<connection>
<GID>5578</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5577</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-426.5,469.5,-426.5</points>
<connection>
<GID>3513</GID>
<name>OUT</name></connection>
<connection>
<GID>3564</GID>
<name>clock</name></connection>
<connection>
<GID>3567</GID>
<name>clock</name></connection>
<connection>
<GID>3570</GID>
<name>clock</name></connection>
<connection>
<GID>3573</GID>
<name>clock</name></connection>
<connection>
<GID>3576</GID>
<name>clock</name></connection>
<connection>
<GID>3579</GID>
<name>clock</name></connection>
<connection>
<GID>3582</GID>
<name>clock</name></connection>
<connection>
<GID>3585</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,400,393.5,400.5</points>
<connection>
<GID>5578</GID>
<name>IN_0</name></connection>
<intersection>400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,400,393.5,400</points>
<intersection>379.5 2</intersection>
<intersection>393.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379.5,400,379.5,413</points>
<intersection>400 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379.5,404.5,383.5,404.5</points>
<connection>
<GID>5577</GID>
<name>IN_0</name></connection>
<intersection>379.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377.5,413,379.5,413</points>
<connection>
<GID>5579</GID>
<name>OUT_0</name></connection>
<intersection>379.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,-450,481.5,-450</points>
<connection>
<GID>3538</GID>
<name>IN_1</name></connection>
<connection>
<GID>3541</GID>
<name>IN_1</name></connection>
<connection>
<GID>3544</GID>
<name>IN_1</name></connection>
<connection>
<GID>3547</GID>
<name>IN_1</name></connection>
<connection>
<GID>3550</GID>
<name>IN_1</name></connection>
<connection>
<GID>3553</GID>
<name>IN_1</name></connection>
<connection>
<GID>3556</GID>
<name>IN_1</name></connection>
<connection>
<GID>3559</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,-450,246,-447.5</points>
<connection>
<GID>3515</GID>
<name>OUT_0</name></connection>
<intersection>-450 1</intersection></vsegment></shape></wire>
<wire>
<ID>3965</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421,403.5,423,403.5</points>
<connection>
<GID>5581</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5580</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-442.5,469,-442.5</points>
<connection>
<GID>3517</GID>
<name>OUT</name></connection>
<connection>
<GID>3540</GID>
<name>clock</name></connection>
<connection>
<GID>3543</GID>
<name>clock</name></connection>
<connection>
<GID>3546</GID>
<name>clock</name></connection>
<connection>
<GID>3549</GID>
<name>clock</name></connection>
<connection>
<GID>3552</GID>
<name>clock</name></connection>
<connection>
<GID>3555</GID>
<name>clock</name></connection>
<connection>
<GID>3558</GID>
<name>clock</name></connection>
<connection>
<GID>3561</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411,400.5,425,400.5</points>
<connection>
<GID>5581</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411,400.5,411,413</points>
<intersection>400.5 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411,404.5,415,404.5</points>
<connection>
<GID>5580</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408.5,413,411,413</points>
<connection>
<GID>5582</GID>
<name>OUT_0</name></connection>
<intersection>411 2</intersection></hsegment></shape></wire>
<wire>
<ID>2423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-459.5,468.5,-459.5</points>
<connection>
<GID>3537</GID>
<name>clock</name></connection>
<connection>
<GID>3534</GID>
<name>clock</name></connection>
<connection>
<GID>3531</GID>
<name>clock</name></connection>
<connection>
<GID>3528</GID>
<name>clock</name></connection>
<connection>
<GID>3525</GID>
<name>clock</name></connection>
<connection>
<GID>3522</GID>
<name>clock</name></connection>
<connection>
<GID>3521</GID>
<name>OUT</name></connection>
<connection>
<GID>3516</GID>
<name>clock</name></connection>
<connection>
<GID>3508</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3967</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451.5,403.5,453.5,403.5</points>
<connection>
<GID>5584</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5583</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,-467,481,-467</points>
<connection>
<GID>3506</GID>
<name>IN_1</name></connection>
<connection>
<GID>3512</GID>
<name>IN_1</name></connection>
<connection>
<GID>3518</GID>
<name>IN_1</name></connection>
<connection>
<GID>3523</GID>
<name>IN_1</name></connection>
<connection>
<GID>3526</GID>
<name>IN_1</name></connection>
<connection>
<GID>3529</GID>
<name>IN_1</name></connection>
<connection>
<GID>3532</GID>
<name>IN_1</name></connection>
<connection>
<GID>3535</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,-467,246,-464.5</points>
<connection>
<GID>3519</GID>
<name>OUT_0</name></connection>
<intersection>-467 1</intersection></vsegment></shape></wire>
<wire>
<ID>3968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,400,455.5,400.5</points>
<connection>
<GID>5584</GID>
<name>IN_0</name></connection>
<intersection>400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,400,455.5,400</points>
<intersection>441.5 2</intersection>
<intersection>455.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441.5,400,441.5,413</points>
<intersection>400 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441.5,404.5,445.5,404.5</points>
<connection>
<GID>5583</GID>
<name>IN_0</name></connection>
<intersection>441.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439.5,413,441.5,413</points>
<connection>
<GID>5585</GID>
<name>OUT_0</name></connection>
<intersection>441.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-476,469,-476</points>
<connection>
<GID>3499</GID>
<name>OUT</name></connection>
<connection>
<GID>3476</GID>
<name>clock</name></connection>
<connection>
<GID>3473</GID>
<name>clock</name></connection>
<connection>
<GID>3470</GID>
<name>clock</name></connection>
<connection>
<GID>3467</GID>
<name>clock</name></connection>
<connection>
<GID>3464</GID>
<name>clock</name></connection>
<connection>
<GID>3461</GID>
<name>clock</name></connection>
<connection>
<GID>3458</GID>
<name>clock</name></connection>
<connection>
<GID>3455</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3969</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483,403.5,485,403.5</points>
<connection>
<GID>5587</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5586</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-483.5,481.5,-483.5</points>
<connection>
<GID>3453</GID>
<name>IN_1</name></connection>
<connection>
<GID>3456</GID>
<name>IN_1</name></connection>
<connection>
<GID>3459</GID>
<name>IN_1</name></connection>
<connection>
<GID>3462</GID>
<name>IN_1</name></connection>
<connection>
<GID>3465</GID>
<name>IN_1</name></connection>
<connection>
<GID>3468</GID>
<name>IN_1</name></connection>
<connection>
<GID>3471</GID>
<name>IN_1</name></connection>
<connection>
<GID>3474</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-483.5,245,-480.5</points>
<connection>
<GID>3498</GID>
<name>OUT_0</name></connection>
<intersection>-483.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3970</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473,400.5,487,400.5</points>
<connection>
<GID>5587</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473,400.5,473,413</points>
<intersection>400.5 1</intersection>
<intersection>404.5 4</intersection>
<intersection>413 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473,404.5,477,404.5</points>
<connection>
<GID>5586</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470.5,413,473,413</points>
<connection>
<GID>5588</GID>
<name>OUT_0</name></connection>
<intersection>473 2</intersection></hsegment></shape></wire>
<wire>
<ID>2427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-491.5,468.5,-491.5</points>
<connection>
<GID>3501</GID>
<name>OUT</name></connection>
<connection>
<GID>3452</GID>
<name>clock</name></connection>
<connection>
<GID>3449</GID>
<name>clock</name></connection>
<connection>
<GID>3446</GID>
<name>clock</name></connection>
<connection>
<GID>3443</GID>
<name>clock</name></connection>
<connection>
<GID>3440</GID>
<name>clock</name></connection>
<connection>
<GID>3437</GID>
<name>clock</name></connection>
<connection>
<GID>3434</GID>
<name>clock</name></connection>
<connection>
<GID>3431</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>3971</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267,419.5,269,419.5</points>
<connection>
<GID>5590</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5589</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-499,481,-499</points>
<connection>
<GID>3429</GID>
<name>IN_1</name></connection>
<connection>
<GID>3432</GID>
<name>IN_1</name></connection>
<connection>
<GID>3435</GID>
<name>IN_1</name></connection>
<connection>
<GID>3438</GID>
<name>IN_1</name></connection>
<connection>
<GID>3441</GID>
<name>IN_1</name></connection>
<connection>
<GID>3444</GID>
<name>IN_1</name></connection>
<connection>
<GID>3447</GID>
<name>IN_1</name></connection>
<connection>
<GID>3450</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-499,245,-496.5</points>
<connection>
<GID>3500</GID>
<name>OUT_0</name></connection>
<intersection>-499 1</intersection></vsegment></shape></wire>
<wire>
<ID>3972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,416,271,416.5</points>
<connection>
<GID>5590</GID>
<name>IN_0</name></connection>
<intersection>416 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,416,271,416</points>
<intersection>257 2</intersection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257,416,257,429</points>
<intersection>416 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,420.5,261,420.5</points>
<connection>
<GID>5589</GID>
<name>IN_0</name></connection>
<intersection>257 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255,429,257,429</points>
<connection>
<GID>5591</GID>
<name>OUT_0</name></connection>
<intersection>257 2</intersection></hsegment></shape></wire>
<wire>
<ID>2429</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301,-531,303,-531</points>
<connection>
<GID>3384</GID>
<name>OUT</name></connection>
<connection>
<GID>3385</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3973</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,419.5,300.5,419.5</points>
<connection>
<GID>5593</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5592</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291,-534,305,-534</points>
<connection>
<GID>3385</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291,-534,291,-521.5</points>
<intersection>-534 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291,-530,295,-530</points>
<connection>
<GID>3384</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>288.5,-521.5,291,-521.5</points>
<connection>
<GID>3386</GID>
<name>OUT_0</name></connection>
<intersection>291 2</intersection></hsegment></shape></wire>
<wire>
<ID>3974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288.5,416.5,302.5,416.5</points>
<connection>
<GID>5593</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288.5,416.5,288.5,429</points>
<intersection>416.5 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,420.5,292.5,420.5</points>
<connection>
<GID>5592</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,429,288.5,429</points>
<connection>
<GID>5594</GID>
<name>OUT_0</name></connection>
<intersection>288.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2431</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>331.5,-531,333.5,-531</points>
<connection>
<GID>3387</GID>
<name>OUT</name></connection>
<connection>
<GID>3388</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3975</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329,419.5,331,419.5</points>
<connection>
<GID>5596</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5595</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-534.5,335.5,-534</points>
<connection>
<GID>3388</GID>
<name>IN_0</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-534.5,335.5,-534.5</points>
<intersection>321.5 2</intersection>
<intersection>335.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321.5,-534.5,321.5,-521.5</points>
<intersection>-534.5 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321.5,-530,325.5,-530</points>
<connection>
<GID>3387</GID>
<name>IN_0</name></connection>
<intersection>321.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>319.5,-521.5,321.5,-521.5</points>
<connection>
<GID>3389</GID>
<name>OUT_0</name></connection>
<intersection>321.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,416,333,416.5</points>
<connection>
<GID>5596</GID>
<name>IN_0</name></connection>
<intersection>416 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,416,333,416</points>
<intersection>319 2</intersection>
<intersection>333 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319,416,319,429</points>
<intersection>416 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,420.5,323,420.5</points>
<connection>
<GID>5595</GID>
<name>IN_0</name></connection>
<intersection>319 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317,429,319,429</points>
<connection>
<GID>5597</GID>
<name>OUT_0</name></connection>
<intersection>319 2</intersection></hsegment></shape></wire>
<wire>
<ID>2433</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363,-531,365,-531</points>
<connection>
<GID>3390</GID>
<name>OUT</name></connection>
<connection>
<GID>3391</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3977</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360.5,419.5,362.5,419.5</points>
<connection>
<GID>5599</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5598</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353,-534,367,-534</points>
<connection>
<GID>3391</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353,-534,353,-521.5</points>
<intersection>-534 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353,-530,357,-530</points>
<connection>
<GID>3390</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>350.5,-521.5,353,-521.5</points>
<connection>
<GID>3392</GID>
<name>OUT_0</name></connection>
<intersection>353 2</intersection></hsegment></shape></wire>
<wire>
<ID>3978</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350.5,416.5,364.5,416.5</points>
<connection>
<GID>5599</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,416.5,350.5,429</points>
<intersection>416.5 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350.5,420.5,354.5,420.5</points>
<connection>
<GID>5598</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348,429,350.5,429</points>
<connection>
<GID>5600</GID>
<name>OUT_0</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2435</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>392.5,-531,394.5,-531</points>
<connection>
<GID>3393</GID>
<name>OUT</name></connection>
<connection>
<GID>3394</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3979</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390,419.5,392,419.5</points>
<connection>
<GID>5602</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5601</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-534.5,396.5,-534</points>
<connection>
<GID>3394</GID>
<name>IN_0</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382.5,-534.5,396.5,-534.5</points>
<intersection>382.5 2</intersection>
<intersection>396.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>382.5,-534.5,382.5,-521.5</points>
<intersection>-534.5 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>382.5,-530,386.5,-530</points>
<connection>
<GID>3393</GID>
<name>IN_0</name></connection>
<intersection>382.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380.5,-521.5,382.5,-521.5</points>
<connection>
<GID>3395</GID>
<name>OUT_0</name></connection>
<intersection>382.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,416,394,416.5</points>
<connection>
<GID>5602</GID>
<name>IN_0</name></connection>
<intersection>416 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,416,394,416</points>
<intersection>380 2</intersection>
<intersection>394 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380,416,380,429</points>
<intersection>416 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,420.5,384,420.5</points>
<connection>
<GID>5601</GID>
<name>IN_0</name></connection>
<intersection>380 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378,429,380,429</points>
<connection>
<GID>5603</GID>
<name>OUT_0</name></connection>
<intersection>380 2</intersection></hsegment></shape></wire>
<wire>
<ID>2437</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424,-531,426,-531</points>
<connection>
<GID>3396</GID>
<name>OUT</name></connection>
<connection>
<GID>3397</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3981</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421.5,419.5,423.5,419.5</points>
<connection>
<GID>5605</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5604</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414,-534,428,-534</points>
<connection>
<GID>3397</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414,-534,414,-521.5</points>
<intersection>-534 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414,-530,418,-530</points>
<connection>
<GID>3396</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411.5,-521.5,414,-521.5</points>
<connection>
<GID>3398</GID>
<name>OUT_0</name></connection>
<intersection>414 2</intersection></hsegment></shape></wire>
<wire>
<ID>3982</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411.5,416.5,425.5,416.5</points>
<connection>
<GID>5605</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411.5,416.5,411.5,429</points>
<intersection>416.5 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411.5,420.5,415.5,420.5</points>
<connection>
<GID>5604</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409,429,411.5,429</points>
<connection>
<GID>5606</GID>
<name>OUT_0</name></connection>
<intersection>411.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2439</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>454.5,-531,456.5,-531</points>
<connection>
<GID>3399</GID>
<name>OUT</name></connection>
<connection>
<GID>3400</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3983</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452,419.5,454,419.5</points>
<connection>
<GID>5608</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5607</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-534.5,458.5,-534</points>
<connection>
<GID>3400</GID>
<name>IN_0</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,-534.5,458.5,-534.5</points>
<intersection>444.5 2</intersection>
<intersection>458.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>444.5,-534.5,444.5,-521.5</points>
<intersection>-534.5 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>444.5,-530,448.5,-530</points>
<connection>
<GID>3399</GID>
<name>IN_0</name></connection>
<intersection>444.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>442.5,-521.5,444.5,-521.5</points>
<connection>
<GID>3401</GID>
<name>OUT_0</name></connection>
<intersection>444.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,416,456,416.5</points>
<connection>
<GID>5608</GID>
<name>IN_0</name></connection>
<intersection>416 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,416,456,416</points>
<intersection>442 2</intersection>
<intersection>456 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442,416,442,429</points>
<intersection>416 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442,420.5,446,420.5</points>
<connection>
<GID>5607</GID>
<name>IN_0</name></connection>
<intersection>442 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,429,442,429</points>
<connection>
<GID>5609</GID>
<name>OUT_0</name></connection>
<intersection>442 2</intersection></hsegment></shape></wire>
<wire>
<ID>2441</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486,-531,488,-531</points>
<connection>
<GID>3402</GID>
<name>OUT</name></connection>
<connection>
<GID>3403</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3985</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483.5,419.5,485.5,419.5</points>
<connection>
<GID>5611</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5610</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2442</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476,-534,490,-534</points>
<connection>
<GID>3403</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476,-534,476,-521.5</points>
<intersection>-534 1</intersection>
<intersection>-530 4</intersection>
<intersection>-521.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476,-530,480,-530</points>
<connection>
<GID>3402</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>473.5,-521.5,476,-521.5</points>
<connection>
<GID>3404</GID>
<name>OUT_0</name></connection>
<intersection>476 2</intersection></hsegment></shape></wire>
<wire>
<ID>3986</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473.5,416.5,487.5,416.5</points>
<connection>
<GID>5611</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473.5,416.5,473.5,429</points>
<intersection>416.5 1</intersection>
<intersection>420.5 4</intersection>
<intersection>429 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473.5,420.5,477.5,420.5</points>
<connection>
<GID>5610</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471,429,473.5,429</points>
<connection>
<GID>5612</GID>
<name>OUT_0</name></connection>
<intersection>473.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2443</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270,-514,272,-514</points>
<connection>
<GID>3405</GID>
<name>OUT</name></connection>
<connection>
<GID>3406</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3987</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267.5,435,269.5,435</points>
<connection>
<GID>5614</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5613</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-517.5,274,-517</points>
<connection>
<GID>3406</GID>
<name>IN_0</name></connection>
<intersection>-517.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-517.5,274,-517.5</points>
<intersection>260 2</intersection>
<intersection>274 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260,-517.5,260,-504.5</points>
<intersection>-517.5 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260,-513,264,-513</points>
<connection>
<GID>3405</GID>
<name>IN_0</name></connection>
<intersection>260 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258,-504.5,260,-504.5</points>
<connection>
<GID>3407</GID>
<name>OUT_0</name></connection>
<intersection>260 2</intersection></hsegment></shape></wire>
<wire>
<ID>3988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,431.5,271.5,432</points>
<connection>
<GID>5614</GID>
<name>IN_0</name></connection>
<intersection>431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,431.5,271.5,431.5</points>
<intersection>257.5 2</intersection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257.5,431.5,257.5,444.5</points>
<intersection>431.5 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257.5,436,261.5,436</points>
<connection>
<GID>5613</GID>
<name>IN_0</name></connection>
<intersection>257.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255.5,444.5,257.5,444.5</points>
<connection>
<GID>5615</GID>
<name>OUT_0</name></connection>
<intersection>257.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2445</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,-514,303.5,-514</points>
<connection>
<GID>3408</GID>
<name>OUT</name></connection>
<connection>
<GID>3409</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3989</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299,435,301,435</points>
<connection>
<GID>5617</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5616</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,-517,305.5,-517</points>
<connection>
<GID>3409</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291.5,-517,291.5,-504.5</points>
<intersection>-517 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291.5,-513,295.5,-513</points>
<connection>
<GID>3408</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289,-504.5,291.5,-504.5</points>
<connection>
<GID>3410</GID>
<name>OUT_0</name></connection>
<intersection>291.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3990</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,432,303,432</points>
<connection>
<GID>5617</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289,432,289,444.5</points>
<intersection>432 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289,436,293,436</points>
<connection>
<GID>5616</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286.5,444.5,289,444.5</points>
<connection>
<GID>5618</GID>
<name>OUT_0</name></connection>
<intersection>289 2</intersection></hsegment></shape></wire>
<wire>
<ID>2447</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332,-514,334,-514</points>
<connection>
<GID>3411</GID>
<name>OUT</name></connection>
<connection>
<GID>3412</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3991</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329.5,435,331.5,435</points>
<connection>
<GID>5620</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5619</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,-517.5,336,-517</points>
<connection>
<GID>3412</GID>
<name>IN_0</name></connection>
<intersection>-517.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-517.5,336,-517.5</points>
<intersection>322 2</intersection>
<intersection>336 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322,-517.5,322,-504.5</points>
<intersection>-517.5 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322,-513,326,-513</points>
<connection>
<GID>3411</GID>
<name>IN_0</name></connection>
<intersection>322 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320,-504.5,322,-504.5</points>
<connection>
<GID>3413</GID>
<name>OUT_0</name></connection>
<intersection>322 2</intersection></hsegment></shape></wire>
<wire>
<ID>3992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,431.5,333.5,432</points>
<connection>
<GID>5620</GID>
<name>IN_0</name></connection>
<intersection>431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,431.5,333.5,431.5</points>
<intersection>319.5 2</intersection>
<intersection>333.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319.5,431.5,319.5,444.5</points>
<intersection>431.5 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319.5,436,323.5,436</points>
<connection>
<GID>5619</GID>
<name>IN_0</name></connection>
<intersection>319.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317.5,444.5,319.5,444.5</points>
<connection>
<GID>5621</GID>
<name>OUT_0</name></connection>
<intersection>319.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2449</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363.5,-514,365.5,-514</points>
<connection>
<GID>3414</GID>
<name>OUT</name></connection>
<connection>
<GID>3415</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3993</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361,435,363,435</points>
<connection>
<GID>5623</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5622</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353.5,-517,367.5,-517</points>
<connection>
<GID>3415</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353.5,-517,353.5,-504.5</points>
<intersection>-517 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353.5,-513,357.5,-513</points>
<connection>
<GID>3414</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351,-504.5,353.5,-504.5</points>
<connection>
<GID>3416</GID>
<name>OUT_0</name></connection>
<intersection>353.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3994</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351,432,365,432</points>
<connection>
<GID>5623</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351,432,351,444.5</points>
<intersection>432 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351,436,355,436</points>
<connection>
<GID>5622</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348.5,444.5,351,444.5</points>
<connection>
<GID>5624</GID>
<name>OUT_0</name></connection>
<intersection>351 2</intersection></hsegment></shape></wire>
<wire>
<ID>2451</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393,-514,395,-514</points>
<connection>
<GID>3417</GID>
<name>OUT</name></connection>
<connection>
<GID>3418</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3995</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390.5,435,392.5,435</points>
<connection>
<GID>5626</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5625</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,-517.5,397,-517</points>
<connection>
<GID>3418</GID>
<name>IN_0</name></connection>
<intersection>-517.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383,-517.5,397,-517.5</points>
<intersection>383 2</intersection>
<intersection>397 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,-517.5,383,-504.5</points>
<intersection>-517.5 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383,-513,387,-513</points>
<connection>
<GID>3417</GID>
<name>IN_0</name></connection>
<intersection>383 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381,-504.5,383,-504.5</points>
<connection>
<GID>3419</GID>
<name>OUT_0</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>3996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,431.5,394.5,432</points>
<connection>
<GID>5626</GID>
<name>IN_0</name></connection>
<intersection>431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,431.5,394.5,431.5</points>
<intersection>380.5 2</intersection>
<intersection>394.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380.5,431.5,380.5,444.5</points>
<intersection>431.5 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380.5,436,384.5,436</points>
<connection>
<GID>5625</GID>
<name>IN_0</name></connection>
<intersection>380.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378.5,444.5,380.5,444.5</points>
<connection>
<GID>5627</GID>
<name>OUT_0</name></connection>
<intersection>380.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2453</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424.5,-514,426.5,-514</points>
<connection>
<GID>3420</GID>
<name>OUT</name></connection>
<connection>
<GID>3421</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3997</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422,435,424,435</points>
<connection>
<GID>5629</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5628</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414.5,-517,428.5,-517</points>
<connection>
<GID>3421</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414.5,-517,414.5,-504.5</points>
<intersection>-517 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414.5,-513,418.5,-513</points>
<connection>
<GID>3420</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412,-504.5,414.5,-504.5</points>
<connection>
<GID>3422</GID>
<name>OUT_0</name></connection>
<intersection>414.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3998</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,432,426,432</points>
<connection>
<GID>5629</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412,432,412,444.5</points>
<intersection>432 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412,436,416,436</points>
<connection>
<GID>5628</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409.5,444.5,412,444.5</points>
<connection>
<GID>5630</GID>
<name>OUT_0</name></connection>
<intersection>412 2</intersection></hsegment></shape></wire>
<wire>
<ID>2455</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455,-514,457,-514</points>
<connection>
<GID>3423</GID>
<name>OUT</name></connection>
<connection>
<GID>3424</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3999</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452.5,435,454.5,435</points>
<connection>
<GID>5632</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5631</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-517.5,459,-517</points>
<connection>
<GID>3424</GID>
<name>IN_0</name></connection>
<intersection>-517.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,-517.5,459,-517.5</points>
<intersection>445 2</intersection>
<intersection>459 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445,-517.5,445,-504.5</points>
<intersection>-517.5 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445,-513,449,-513</points>
<connection>
<GID>3423</GID>
<name>IN_0</name></connection>
<intersection>445 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443,-504.5,445,-504.5</points>
<connection>
<GID>3425</GID>
<name>OUT_0</name></connection>
<intersection>445 2</intersection></hsegment></shape></wire>
<wire>
<ID>4000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,431.5,456.5,432</points>
<connection>
<GID>5632</GID>
<name>IN_0</name></connection>
<intersection>431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,431.5,456.5,431.5</points>
<intersection>442.5 2</intersection>
<intersection>456.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442.5,431.5,442.5,444.5</points>
<intersection>431.5 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442.5,436,446.5,436</points>
<connection>
<GID>5631</GID>
<name>IN_0</name></connection>
<intersection>442.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,444.5,442.5,444.5</points>
<connection>
<GID>5633</GID>
<name>OUT_0</name></connection>
<intersection>442.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2457</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486.5,-514,488.5,-514</points>
<connection>
<GID>3426</GID>
<name>OUT</name></connection>
<connection>
<GID>3427</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4001</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484,435,486,435</points>
<connection>
<GID>5635</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5634</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476.5,-517,490.5,-517</points>
<connection>
<GID>3427</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476.5,-517,476.5,-504.5</points>
<intersection>-517 1</intersection>
<intersection>-513 4</intersection>
<intersection>-504.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476.5,-513,480.5,-513</points>
<connection>
<GID>3426</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474,-504.5,476.5,-504.5</points>
<connection>
<GID>3428</GID>
<name>OUT_0</name></connection>
<intersection>476.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4002</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474,432,488,432</points>
<connection>
<GID>5635</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474,432,474,444.5</points>
<intersection>432 1</intersection>
<intersection>436 4</intersection>
<intersection>444.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474,436,478,436</points>
<connection>
<GID>5634</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471.5,444.5,474,444.5</points>
<connection>
<GID>5636</GID>
<name>OUT_0</name></connection>
<intersection>474 2</intersection></hsegment></shape></wire>
<wire>
<ID>2459</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270.5,-498,272.5,-498</points>
<connection>
<GID>3429</GID>
<name>OUT</name></connection>
<connection>
<GID>3430</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4003</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,410,464.5,410</points>
<connection>
<GID>5663</GID>
<name>OUT</name></connection>
<connection>
<GID>5588</GID>
<name>clock</name></connection>
<connection>
<GID>5585</GID>
<name>clock</name></connection>
<connection>
<GID>5582</GID>
<name>clock</name></connection>
<connection>
<GID>5579</GID>
<name>clock</name></connection>
<connection>
<GID>5576</GID>
<name>clock</name></connection>
<connection>
<GID>5573</GID>
<name>clock</name></connection>
<connection>
<GID>5570</GID>
<name>clock</name></connection>
<connection>
<GID>5567</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-501.5,274.5,-501</points>
<connection>
<GID>3430</GID>
<name>IN_0</name></connection>
<intersection>-501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-501.5,274.5,-501.5</points>
<intersection>260.5 2</intersection>
<intersection>274.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260.5,-501.5,260.5,-488.5</points>
<intersection>-501.5 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,-497,264.5,-497</points>
<connection>
<GID>3429</GID>
<name>IN_0</name></connection>
<intersection>260.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258.5,-488.5,260.5,-488.5</points>
<connection>
<GID>3431</GID>
<name>OUT_0</name></connection>
<intersection>260.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4004</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241.5,402.5,477,402.5</points>
<connection>
<GID>5586</GID>
<name>IN_1</name></connection>
<connection>
<GID>5583</GID>
<name>IN_1</name></connection>
<connection>
<GID>5580</GID>
<name>IN_1</name></connection>
<connection>
<GID>5577</GID>
<name>IN_1</name></connection>
<connection>
<GID>5574</GID>
<name>IN_1</name></connection>
<connection>
<GID>5571</GID>
<name>IN_1</name></connection>
<connection>
<GID>5568</GID>
<name>IN_1</name></connection>
<connection>
<GID>5565</GID>
<name>IN_1</name></connection>
<intersection>241.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241.5,402.5,241.5,405</points>
<connection>
<GID>5662</GID>
<name>OUT_0</name></connection>
<intersection>402.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2461</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302,-498,304,-498</points>
<connection>
<GID>3432</GID>
<name>OUT</name></connection>
<connection>
<GID>3433</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4005</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,393,464,393</points>
<connection>
<GID>5665</GID>
<name>OUT</name></connection>
<connection>
<GID>5564</GID>
<name>clock</name></connection>
<connection>
<GID>5561</GID>
<name>clock</name></connection>
<connection>
<GID>5558</GID>
<name>clock</name></connection>
<connection>
<GID>5555</GID>
<name>clock</name></connection>
<connection>
<GID>5552</GID>
<name>clock</name></connection>
<connection>
<GID>5549</GID>
<name>clock</name></connection>
<connection>
<GID>5546</GID>
<name>clock</name></connection>
<connection>
<GID>5532</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-501,306,-501</points>
<connection>
<GID>3433</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292,-501,292,-488.5</points>
<intersection>-501 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292,-497,296,-497</points>
<connection>
<GID>3432</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289.5,-488.5,292,-488.5</points>
<connection>
<GID>3434</GID>
<name>OUT_0</name></connection>
<intersection>292 2</intersection></hsegment></shape></wire>
<wire>
<ID>4006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,385.5,242.5,388</points>
<intersection>385.5 2</intersection>
<intersection>388 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>242.5,385.5,476.5,385.5</points>
<connection>
<GID>5562</GID>
<name>IN_1</name></connection>
<connection>
<GID>5559</GID>
<name>IN_1</name></connection>
<connection>
<GID>5556</GID>
<name>IN_1</name></connection>
<connection>
<GID>5553</GID>
<name>IN_1</name></connection>
<connection>
<GID>5550</GID>
<name>IN_1</name></connection>
<connection>
<GID>5547</GID>
<name>IN_1</name></connection>
<connection>
<GID>5544</GID>
<name>IN_1</name></connection>
<connection>
<GID>5530</GID>
<name>IN_1</name></connection>
<intersection>242.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>241.5,388,242.5,388</points>
<connection>
<GID>5664</GID>
<name>OUT_0</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2463</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332.5,-498,334.5,-498</points>
<connection>
<GID>3435</GID>
<name>OUT</name></connection>
<connection>
<GID>3436</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4007</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,376,278,509.5</points>
<connection>
<GID>5534</GID>
<name>N_in1</name></connection>
<intersection>396 1</intersection>
<intersection>413 3</intersection>
<intersection>429 4</intersection>
<intersection>444.5 5</intersection>
<intersection>461 6</intersection>
<intersection>478 7</intersection>
<intersection>494 8</intersection>
<intersection>509.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,396,279,396</points>
<connection>
<GID>5546</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278,509.5,281.5,509.5</points>
<connection>
<GID>5751</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>278,413,279.5,413</points>
<connection>
<GID>5570</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>278,429,280,429</points>
<connection>
<GID>5594</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>278,444.5,280.5,444.5</points>
<connection>
<GID>5618</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>278,461,280,461</points>
<connection>
<GID>5676</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>278,478,280.5,478</points>
<connection>
<GID>5703</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>278,494,281,494</points>
<connection>
<GID>5727</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>2464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,-501.5,336.5,-501</points>
<connection>
<GID>3436</GID>
<name>IN_0</name></connection>
<intersection>-501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,-501.5,336.5,-501.5</points>
<intersection>322.5 2</intersection>
<intersection>336.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322.5,-501.5,322.5,-488.5</points>
<intersection>-501.5 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322.5,-497,326.5,-497</points>
<connection>
<GID>3435</GID>
<name>IN_0</name></connection>
<intersection>322.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320.5,-488.5,322.5,-488.5</points>
<connection>
<GID>3437</GID>
<name>OUT_0</name></connection>
<intersection>322.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,376,310,509.5</points>
<connection>
<GID>5535</GID>
<name>N_in1</name></connection>
<connection>
<GID>5549</GID>
<name>IN_0</name></connection>
<intersection>413 9</intersection>
<intersection>429 10</intersection>
<intersection>444.5 7</intersection>
<intersection>461 11</intersection>
<intersection>478 5</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,509.5,312.5,509.5</points>
<connection>
<GID>5754</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,494,312,494</points>
<connection>
<GID>5730</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>310,478,311.5,478</points>
<connection>
<GID>5706</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>310,444.5,311.5,444.5</points>
<connection>
<GID>5621</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>310,413,310.5,413</points>
<connection>
<GID>5573</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>310,429,311,429</points>
<connection>
<GID>5597</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>310,461,311,461</points>
<connection>
<GID>5682</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>2465</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364,-498,366,-498</points>
<connection>
<GID>3438</GID>
<name>OUT</name></connection>
<connection>
<GID>3439</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4009</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341,377,341,509.5</points>
<connection>
<GID>5552</GID>
<name>IN_0</name></connection>
<connection>
<GID>5536</GID>
<name>N_in1</name></connection>
<intersection>413 38</intersection>
<intersection>429 21</intersection>
<intersection>444.5 7</intersection>
<intersection>461 20</intersection>
<intersection>478 5</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>341,509.5,343.5,509.5</points>
<connection>
<GID>5757</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341,494,343,494</points>
<connection>
<GID>5733</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>341,478,342.5,478</points>
<connection>
<GID>5709</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>341,444.5,342.5,444.5</points>
<connection>
<GID>5624</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>341,461,342,461</points>
<connection>
<GID>5685</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>341,429,342,429</points>
<connection>
<GID>5600</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>341,413,341.5,413</points>
<connection>
<GID>5576</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection></hsegment></shape></wire>
<wire>
<ID>2466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354,-501,368,-501</points>
<connection>
<GID>3439</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354,-501,354,-488.5</points>
<intersection>-501 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354,-497,358,-497</points>
<connection>
<GID>3438</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351.5,-488.5,354,-488.5</points>
<connection>
<GID>3440</GID>
<name>OUT_0</name></connection>
<intersection>354 2</intersection></hsegment></shape></wire>
<wire>
<ID>4010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,413,372,509.5</points>
<connection>
<GID>5688</GID>
<name>IN_0</name></connection>
<connection>
<GID>5603</GID>
<name>IN_0</name></connection>
<intersection>413 9</intersection>
<intersection>444.5 7</intersection>
<intersection>478 5</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372,509.5,373.5,509.5</points>
<connection>
<GID>5760</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,494,373,494</points>
<connection>
<GID>5736</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>372,478,372.5,478</points>
<connection>
<GID>5712</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>372,444.5,372.5,444.5</points>
<connection>
<GID>5627</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>371,413,372,413</points>
<connection>
<GID>5579</GID>
<name>IN_0</name></connection>
<intersection>371 10</intersection>
<intersection>372 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>371,378,371,413</points>
<connection>
<GID>5555</GID>
<name>IN_0</name></connection>
<connection>
<GID>5537</GID>
<name>N_in1</name></connection>
<intersection>413 9</intersection></vsegment></shape></wire>
<wire>
<ID>2467</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393.5,-498,395.5,-498</points>
<connection>
<GID>3441</GID>
<name>OUT</name></connection>
<connection>
<GID>3442</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402,378.5,402,509.5</points>
<connection>
<GID>5558</GID>
<name>IN_0</name></connection>
<connection>
<GID>5538</GID>
<name>N_in1</name></connection>
<intersection>413 13</intersection>
<intersection>429 11</intersection>
<intersection>444.5 9</intersection>
<intersection>461 7</intersection>
<intersection>478 5</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,509.5,404.5,509.5</points>
<connection>
<GID>5763</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>402,494,404,494</points>
<connection>
<GID>5739</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>402,478,403.5,478</points>
<connection>
<GID>5715</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>402,461,403,461</points>
<connection>
<GID>5691</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>402,444.5,403.5,444.5</points>
<connection>
<GID>5630</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>402,429,403,429</points>
<connection>
<GID>5606</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>402,413,402.5,413</points>
<connection>
<GID>5582</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment></shape></wire>
<wire>
<ID>2468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,-501.5,397.5,-501</points>
<connection>
<GID>3442</GID>
<name>IN_0</name></connection>
<intersection>-501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,-501.5,397.5,-501.5</points>
<intersection>383.5 2</intersection>
<intersection>397.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,-501.5,383.5,-488.5</points>
<intersection>-501.5 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383.5,-497,387.5,-497</points>
<connection>
<GID>3441</GID>
<name>IN_0</name></connection>
<intersection>383.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381.5,-488.5,383.5,-488.5</points>
<connection>
<GID>3443</GID>
<name>OUT_0</name></connection>
<intersection>383.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433,379.5,433,509.5</points>
<connection>
<GID>5561</GID>
<name>IN_0</name></connection>
<connection>
<GID>5540</GID>
<name>N_in1</name></connection>
<intersection>413 13</intersection>
<intersection>429 11</intersection>
<intersection>444.5 9</intersection>
<intersection>461 7</intersection>
<intersection>478 5</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433,509.5,435.5,509.5</points>
<connection>
<GID>5766</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433,494,435,494</points>
<connection>
<GID>5742</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>433,478,434.5,478</points>
<connection>
<GID>5718</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>433,461,434,461</points>
<connection>
<GID>5694</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>433,444.5,434.5,444.5</points>
<connection>
<GID>5633</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>433,429,434,429</points>
<connection>
<GID>5609</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>433,413,433.5,413</points>
<connection>
<GID>5585</GID>
<name>IN_0</name></connection>
<intersection>433 0</intersection></hsegment></shape></wire>
<wire>
<ID>2469</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425,-498,427,-498</points>
<connection>
<GID>3444</GID>
<name>OUT</name></connection>
<connection>
<GID>3445</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464,377.5,464,509.5</points>
<connection>
<GID>5564</GID>
<name>IN_0</name></connection>
<connection>
<GID>5539</GID>
<name>N_in1</name></connection>
<intersection>413 13</intersection>
<intersection>429 10</intersection>
<intersection>444.5 8</intersection>
<intersection>461 6</intersection>
<intersection>478 4</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>464,509.5,466.5,509.5</points>
<connection>
<GID>5769</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,494,466,494</points>
<connection>
<GID>5745</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>464,478,465.5,478</points>
<connection>
<GID>5721</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>464,461,465,461</points>
<connection>
<GID>5697</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>464,444.5,465.5,444.5</points>
<connection>
<GID>5636</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>464,429,465,429</points>
<connection>
<GID>5612</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>464,413,464.5,413</points>
<connection>
<GID>5588</GID>
<name>IN_0</name></connection>
<intersection>464 0</intersection></hsegment></shape></wire>
<wire>
<ID>2470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415,-501,429,-501</points>
<connection>
<GID>3445</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415,-501,415,-488.5</points>
<intersection>-501 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415,-497,419,-497</points>
<connection>
<GID>3444</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412.5,-488.5,415,-488.5</points>
<connection>
<GID>3446</GID>
<name>OUT_0</name></connection>
<intersection>415 2</intersection></hsegment></shape></wire>
<wire>
<ID>4014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,368,276,523</points>
<connection>
<GID>5642</GID>
<name>N_in0</name></connection>
<connection>
<GID>5643</GID>
<name>N_in1</name></connection>
<intersection>388 13</intersection>
<intersection>405 12</intersection>
<intersection>421 11</intersection>
<intersection>436.5 10</intersection>
<intersection>453 9</intersection>
<intersection>470 8</intersection>
<intersection>487.5 7</intersection>
<intersection>502.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>272.5,502.5,276,502.5</points>
<connection>
<GID>5747</GID>
<name>OUT_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>272,487.5,276,487.5</points>
<intersection>272 22</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>271.5,470,276,470</points>
<intersection>271.5 21</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>271,453,276,453</points>
<intersection>271 20</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>271.5,436.5,276,436.5</points>
<intersection>271.5 17</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>271,421,276,421</points>
<intersection>271 16</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>270.5,405,276,405</points>
<intersection>270.5 15</intersection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>270,388,276,388</points>
<intersection>270 14</intersection>
<intersection>276 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>270,388,270,389</points>
<connection>
<GID>5531</GID>
<name>OUT_0</name></connection>
<intersection>388 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>270.5,405,270.5,406</points>
<connection>
<GID>5566</GID>
<name>OUT_0</name></connection>
<intersection>405 12</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>271,421,271,422</points>
<connection>
<GID>5590</GID>
<name>OUT_0</name></connection>
<intersection>421 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>271.5,436.5,271.5,437.5</points>
<connection>
<GID>5614</GID>
<name>OUT_0</name></connection>
<intersection>436.5 10</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>271,453,271,454</points>
<connection>
<GID>5667</GID>
<name>OUT_0</name></connection>
<intersection>453 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>271.5,470,271.5,471</points>
<connection>
<GID>5699</GID>
<name>OUT_0</name></connection>
<intersection>470 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>272,487,272,487.5</points>
<connection>
<GID>5723</GID>
<name>OUT_0</name></connection>
<intersection>487.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>2471</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455.5,-498,457.5,-498</points>
<connection>
<GID>3447</GID>
<name>OUT</name></connection>
<connection>
<GID>3448</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,368.5,305.5,523</points>
<connection>
<GID>5771</GID>
<name>N_in1</name></connection>
<intersection>389 13</intersection>
<intersection>406 12</intersection>
<intersection>422 11</intersection>
<intersection>437.5 10</intersection>
<intersection>454 9</intersection>
<intersection>471 8</intersection>
<intersection>487 7</intersection>
<intersection>502.5 6</intersection>
<intersection>523 23</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>304,502.5,305.5,502.5</points>
<connection>
<GID>5750</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>303.5,487,305.5,487</points>
<connection>
<GID>5726</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>303,471,305.5,471</points>
<connection>
<GID>5702</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>302.5,454,305.5,454</points>
<connection>
<GID>5674</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>303,437.5,305.5,437.5</points>
<connection>
<GID>5617</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>302.5,422,305.5,422</points>
<connection>
<GID>5593</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>302,406,305.5,406</points>
<connection>
<GID>5569</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>301.5,389,305.5,389</points>
<connection>
<GID>5545</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>305.5,523,307,523</points>
<connection>
<GID>5656</GID>
<name>N_in0</name></connection>
<intersection>305.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-501.5,459.5,-501</points>
<connection>
<GID>3448</GID>
<name>IN_0</name></connection>
<intersection>-501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,-501.5,459.5,-501.5</points>
<intersection>445.5 2</intersection>
<intersection>459.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445.5,-501.5,445.5,-488.5</points>
<intersection>-501.5 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445.5,-497,449.5,-497</points>
<connection>
<GID>3447</GID>
<name>IN_0</name></connection>
<intersection>445.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443.5,-488.5,445.5,-488.5</points>
<connection>
<GID>3449</GID>
<name>OUT_0</name></connection>
<intersection>445.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339,369,339,523</points>
<connection>
<GID>5655</GID>
<name>N_in0</name></connection>
<connection>
<GID>5644</GID>
<name>N_in1</name></connection>
<intersection>389 13</intersection>
<intersection>406 12</intersection>
<intersection>422 11</intersection>
<intersection>437.5 10</intersection>
<intersection>454 9</intersection>
<intersection>471 8</intersection>
<intersection>487 7</intersection>
<intersection>502.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>334.5,502.5,339,502.5</points>
<connection>
<GID>5753</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>334,487,339,487</points>
<connection>
<GID>5729</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>333.5,471,339,471</points>
<connection>
<GID>5705</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>333,454,339,454</points>
<connection>
<GID>5680</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>333.5,437.5,339,437.5</points>
<connection>
<GID>5620</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>333,422,339,422</points>
<connection>
<GID>5596</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>332.5,406,339,406</points>
<connection>
<GID>5572</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>332,389,339,389</points>
<connection>
<GID>5548</GID>
<name>OUT_0</name></connection>
<intersection>339 0</intersection></hsegment></shape></wire>
<wire>
<ID>2473</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487,-498,489,-498</points>
<connection>
<GID>3450</GID>
<name>OUT</name></connection>
<connection>
<GID>3451</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369.5,369.5,369.5,523</points>
<connection>
<GID>5654</GID>
<name>N_in0</name></connection>
<connection>
<GID>5645</GID>
<name>N_in1</name></connection>
<intersection>389 18</intersection>
<intersection>406 17</intersection>
<intersection>422 16</intersection>
<intersection>437.5 15</intersection>
<intersection>454 14</intersection>
<intersection>471 13</intersection>
<intersection>487 12</intersection>
<intersection>502.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>366,502.5,369.5,502.5</points>
<connection>
<GID>5756</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>365.5,487,369.5,487</points>
<connection>
<GID>5732</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>365,471,369.5,471</points>
<connection>
<GID>5708</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>364.5,454,369.5,454</points>
<connection>
<GID>5684</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>365,437.5,369.5,437.5</points>
<connection>
<GID>5623</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>364.5,422,369.5,422</points>
<connection>
<GID>5599</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>364,406,369.5,406</points>
<connection>
<GID>5575</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>363.5,389,369.5,389</points>
<connection>
<GID>5551</GID>
<name>OUT_0</name></connection>
<intersection>369.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,-501,491,-501</points>
<connection>
<GID>3451</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477,-501,477,-488.5</points>
<intersection>-501 1</intersection>
<intersection>-497 4</intersection>
<intersection>-488.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477,-497,481,-497</points>
<connection>
<GID>3450</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474.5,-488.5,477,-488.5</points>
<connection>
<GID>3452</GID>
<name>OUT_0</name></connection>
<intersection>477 2</intersection></hsegment></shape></wire>
<wire>
<ID>4018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,369.5,400,523</points>
<connection>
<GID>5653</GID>
<name>N_in0</name></connection>
<connection>
<GID>5646</GID>
<name>N_in1</name></connection>
<intersection>389 9</intersection>
<intersection>406 10</intersection>
<intersection>422 11</intersection>
<intersection>437.5 12</intersection>
<intersection>454 13</intersection>
<intersection>471 14</intersection>
<intersection>487 15</intersection>
<intersection>502.5 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>393,389,400,389</points>
<connection>
<GID>5554</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>393.5,406,400,406</points>
<connection>
<GID>5578</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>394,422,400,422</points>
<connection>
<GID>5602</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>394.5,437.5,400,437.5</points>
<connection>
<GID>5626</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>394,454,400,454</points>
<connection>
<GID>5687</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>394.5,471,400,471</points>
<connection>
<GID>5711</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>395,487,400,487</points>
<connection>
<GID>5735</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>395.5,502.5,400,502.5</points>
<connection>
<GID>5759</GID>
<name>OUT_0</name></connection>
<intersection>400 0</intersection></hsegment></shape></wire>
<wire>
<ID>2475</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271,-482.5,273,-482.5</points>
<connection>
<GID>3453</GID>
<name>OUT</name></connection>
<connection>
<GID>3454</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431,369.5,431,523</points>
<connection>
<GID>5652</GID>
<name>N_in0</name></connection>
<connection>
<GID>5647</GID>
<name>N_in1</name></connection>
<intersection>389 6</intersection>
<intersection>406 7</intersection>
<intersection>422 8</intersection>
<intersection>437.5 9</intersection>
<intersection>454 10</intersection>
<intersection>471 11</intersection>
<intersection>487 12</intersection>
<intersection>502.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>424.5,389,431,389</points>
<connection>
<GID>5557</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>425,406,431,406</points>
<connection>
<GID>5581</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>425.5,422,431,422</points>
<connection>
<GID>5605</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>426,437.5,431,437.5</points>
<connection>
<GID>5629</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>425.5,454,431,454</points>
<connection>
<GID>5690</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>426,471,431,471</points>
<connection>
<GID>5714</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>426.5,487,431,487</points>
<connection>
<GID>5738</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>427,502.5,431,502.5</points>
<connection>
<GID>5762</GID>
<name>OUT_0</name></connection>
<intersection>431 0</intersection></hsegment></shape></wire>
<wire>
<ID>2476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-486,275,-485.5</points>
<connection>
<GID>3454</GID>
<name>IN_0</name></connection>
<intersection>-486 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-486,275,-486</points>
<intersection>261 2</intersection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261,-486,261,-473</points>
<intersection>-486 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,-481.5,265,-481.5</points>
<connection>
<GID>3453</GID>
<name>IN_0</name></connection>
<intersection>261 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259,-473,261,-473</points>
<connection>
<GID>3455</GID>
<name>OUT_0</name></connection>
<intersection>261 2</intersection></hsegment></shape></wire>
<wire>
<ID>4020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462,369,462,524</points>
<connection>
<GID>5651</GID>
<name>N_in0</name></connection>
<connection>
<GID>5648</GID>
<name>N_in1</name></connection>
<intersection>389 6</intersection>
<intersection>406 7</intersection>
<intersection>422 8</intersection>
<intersection>437.5 9</intersection>
<intersection>454 10</intersection>
<intersection>471 11</intersection>
<intersection>487 12</intersection>
<intersection>502.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>455,389,462,389</points>
<connection>
<GID>5560</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>455.5,406,462,406</points>
<connection>
<GID>5584</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>456,422,462,422</points>
<connection>
<GID>5608</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>456.5,437.5,462,437.5</points>
<connection>
<GID>5632</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>456,454,462,454</points>
<connection>
<GID>5693</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>456.5,471,462,471</points>
<connection>
<GID>5717</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>457,487,462,487</points>
<connection>
<GID>5741</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>457.5,502.5,462,502.5</points>
<connection>
<GID>5765</GID>
<name>OUT_0</name></connection>
<intersection>462 0</intersection></hsegment></shape></wire>
<wire>
<ID>2477</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302.5,-482.5,304.5,-482.5</points>
<connection>
<GID>3456</GID>
<name>OUT</name></connection>
<connection>
<GID>3457</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,369.5,492.5,524.5</points>
<connection>
<GID>5650</GID>
<name>N_in0</name></connection>
<connection>
<GID>5649</GID>
<name>N_in1</name></connection>
<intersection>389 3</intersection>
<intersection>406 4</intersection>
<intersection>422 5</intersection>
<intersection>437.5 6</intersection>
<intersection>454 7</intersection>
<intersection>471 8</intersection>
<intersection>487 9</intersection>
<intersection>502.5 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>486.5,389,492.5,389</points>
<connection>
<GID>5563</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>487,406,492.5,406</points>
<connection>
<GID>5587</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>487.5,422,492.5,422</points>
<connection>
<GID>5611</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>488,437.5,492.5,437.5</points>
<connection>
<GID>5635</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>487.5,454,492.5,454</points>
<connection>
<GID>5696</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>488,471,492.5,471</points>
<connection>
<GID>5720</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>488.5,487,492.5,487</points>
<connection>
<GID>5744</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>489,502.5,492.5,502.5</points>
<connection>
<GID>5768</GID>
<name>OUT_0</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-485.5,306.5,-485.5</points>
<connection>
<GID>3457</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292.5,-485.5,292.5,-473</points>
<intersection>-485.5 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-481.5,296.5,-481.5</points>
<connection>
<GID>3456</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290,-473,292.5,-473</points>
<connection>
<GID>3458</GID>
<name>OUT_0</name></connection>
<intersection>292.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,455,201,504</points>
<intersection>455 2</intersection>
<intersection>504 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,504,240,504</points>
<connection>
<GID>5669</GID>
<name>ENABLE_0</name></connection>
<intersection>201 0</intersection>
<intersection>226 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,455,201,455</points>
<connection>
<GID>5657</GID>
<name>OUT_7</name></connection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226,504,226,507.5</points>
<intersection>504 1</intersection>
<intersection>507.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226,507.5,230.5,507.5</points>
<connection>
<GID>5670</GID>
<name>IN_0</name></connection>
<intersection>226 4</intersection></hsegment></shape></wire>
<wire>
<ID>2479</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333,-482.5,335,-482.5</points>
<connection>
<GID>3459</GID>
<name>OUT</name></connection>
<connection>
<GID>3460</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,454,203,488.5</points>
<intersection>454 2</intersection>
<intersection>488.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,488.5,240,488.5</points>
<intersection>203 0</intersection>
<intersection>226 4</intersection>
<intersection>240 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,454,203,454</points>
<connection>
<GID>5657</GID>
<name>OUT_6</name></connection>
<intersection>203 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240,488,240,488.5</points>
<connection>
<GID>5671</GID>
<name>ENABLE_0</name></connection>
<intersection>488.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>226,488.5,226,492</points>
<intersection>488.5 1</intersection>
<intersection>492 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226,492,230,492</points>
<connection>
<GID>5673</GID>
<name>IN_0</name></connection>
<intersection>226 4</intersection></hsegment></shape></wire>
<wire>
<ID>2480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-486,337,-485.5</points>
<connection>
<GID>3460</GID>
<name>IN_0</name></connection>
<intersection>-486 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,-486,337,-486</points>
<intersection>323 2</intersection>
<intersection>337 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323,-486,323,-473</points>
<intersection>-486 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323,-481.5,327,-481.5</points>
<connection>
<GID>3459</GID>
<name>IN_0</name></connection>
<intersection>323 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321,-473,323,-473</points>
<connection>
<GID>3461</GID>
<name>OUT_0</name></connection>
<intersection>323 2</intersection></hsegment></shape></wire>
<wire>
<ID>4024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,453,205,476</points>
<intersection>453 2</intersection>
<intersection>476 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205,476,230,476</points>
<connection>
<GID>5677</GID>
<name>IN_0</name></connection>
<intersection>205 0</intersection>
<intersection>226 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,453,205,453</points>
<connection>
<GID>5657</GID>
<name>OUT_5</name></connection>
<intersection>205 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>226,472,226,476</points>
<intersection>472 4</intersection>
<intersection>476 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>226,472,240,472</points>
<connection>
<GID>5675</GID>
<name>ENABLE_0</name></connection>
<intersection>226 3</intersection></hsegment></shape></wire>
<wire>
<ID>2481</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364.5,-482.5,366.5,-482.5</points>
<connection>
<GID>3462</GID>
<name>OUT</name></connection>
<connection>
<GID>3463</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4025</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,452,207,459</points>
<intersection>452 2</intersection>
<intersection>459 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,459,230,459</points>
<connection>
<GID>5681</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection>
<intersection>226 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,452,207,452</points>
<connection>
<GID>5657</GID>
<name>OUT_4</name></connection>
<intersection>207 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>226,455,226,459</points>
<intersection>455 4</intersection>
<intersection>459 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>226,455,240,455</points>
<connection>
<GID>5679</GID>
<name>ENABLE_0</name></connection>
<intersection>226 3</intersection></hsegment></shape></wire>
<wire>
<ID>2482</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-485.5,368.5,-485.5</points>
<connection>
<GID>3463</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354.5,-485.5,354.5,-473</points>
<intersection>-485.5 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354.5,-481.5,358.5,-481.5</points>
<connection>
<GID>3462</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352,-473,354.5,-473</points>
<connection>
<GID>3464</GID>
<name>OUT_0</name></connection>
<intersection>354.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4026</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,439,207,451</points>
<intersection>439 1</intersection>
<intersection>451 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,439,239,439</points>
<connection>
<GID>5658</GID>
<name>ENABLE_0</name></connection>
<intersection>207 0</intersection>
<intersection>226 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,451,207,451</points>
<connection>
<GID>5657</GID>
<name>OUT_3</name></connection>
<intersection>207 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226,439,226,442.5</points>
<intersection>439 1</intersection>
<intersection>442.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226,442.5,230,442.5</points>
<connection>
<GID>5659</GID>
<name>IN_0</name></connection>
<intersection>226 4</intersection></hsegment></shape></wire>
<wire>
<ID>2483</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394,-482.5,396,-482.5</points>
<connection>
<GID>3465</GID>
<name>OUT</name></connection>
<connection>
<GID>3466</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4027</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,423,205,450</points>
<intersection>423 1</intersection>
<intersection>450 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205,423,239,423</points>
<connection>
<GID>5660</GID>
<name>ENABLE_0</name></connection>
<intersection>205 0</intersection>
<intersection>226 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,450,205,450</points>
<connection>
<GID>5657</GID>
<name>OUT_2</name></connection>
<intersection>205 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226,423,226,427</points>
<intersection>423 1</intersection>
<intersection>427 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226,427,230,427</points>
<connection>
<GID>5661</GID>
<name>IN_0</name></connection>
<intersection>226 4</intersection></hsegment></shape></wire>
<wire>
<ID>2484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,-486,398,-485.5</points>
<connection>
<GID>3466</GID>
<name>IN_0</name></connection>
<intersection>-486 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-486,398,-486</points>
<intersection>384 2</intersection>
<intersection>398 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384,-486,384,-473</points>
<intersection>-486 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384,-481.5,388,-481.5</points>
<connection>
<GID>3465</GID>
<name>IN_0</name></connection>
<intersection>384 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382,-473,384,-473</points>
<connection>
<GID>3467</GID>
<name>OUT_0</name></connection>
<intersection>384 2</intersection></hsegment></shape></wire>
<wire>
<ID>4028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,407.5,203,449</points>
<intersection>407.5 1</intersection>
<intersection>449 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,407.5,239,407.5</points>
<intersection>203 0</intersection>
<intersection>226 4</intersection>
<intersection>239 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,449,203,449</points>
<connection>
<GID>5657</GID>
<name>OUT_1</name></connection>
<intersection>203 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239,407,239,407.5</points>
<connection>
<GID>5662</GID>
<name>ENABLE_0</name></connection>
<intersection>407.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>226,407.5,226,411</points>
<intersection>407.5 1</intersection>
<intersection>411 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226,411,230,411</points>
<connection>
<GID>5663</GID>
<name>IN_0</name></connection>
<intersection>226 4</intersection></hsegment></shape></wire>
<wire>
<ID>2485</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425.5,-482.5,427.5,-482.5</points>
<connection>
<GID>3468</GID>
<name>OUT</name></connection>
<connection>
<GID>3469</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4029</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,390,201,448</points>
<intersection>390 1</intersection>
<intersection>448 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,390,239,390</points>
<connection>
<GID>5664</GID>
<name>ENABLE_0</name></connection>
<intersection>201 0</intersection>
<intersection>226 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,448,201,448</points>
<connection>
<GID>5657</GID>
<name>OUT_0</name></connection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>226,390,226,394</points>
<intersection>390 1</intersection>
<intersection>394 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>226,394,230,394</points>
<connection>
<GID>5665</GID>
<name>IN_0</name></connection>
<intersection>226 4</intersection></hsegment></shape></wire>
<wire>
<ID>2486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415.5,-485.5,429.5,-485.5</points>
<connection>
<GID>3469</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415.5,-485.5,415.5,-473</points>
<intersection>-485.5 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415.5,-481.5,419.5,-481.5</points>
<connection>
<GID>3468</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413,-473,415.5,-473</points>
<connection>
<GID>3470</GID>
<name>OUT_0</name></connection>
<intersection>415.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4030</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267,451.5,269,451.5</points>
<connection>
<GID>5667</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5666</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2487</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456,-482.5,458,-482.5</points>
<connection>
<GID>3471</GID>
<name>OUT</name></connection>
<connection>
<GID>3472</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,448,271,448.5</points>
<connection>
<GID>5667</GID>
<name>IN_0</name></connection>
<intersection>448 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,448,271,448</points>
<intersection>257 2</intersection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257,448,257,461</points>
<intersection>448 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,452.5,261,452.5</points>
<connection>
<GID>5666</GID>
<name>IN_0</name></connection>
<intersection>257 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255,461,257,461</points>
<connection>
<GID>5668</GID>
<name>OUT_0</name></connection>
<intersection>257 2</intersection></hsegment></shape></wire>
<wire>
<ID>2488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460,-486,460,-485.5</points>
<connection>
<GID>3472</GID>
<name>IN_0</name></connection>
<intersection>-486 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446,-486,460,-486</points>
<intersection>446 2</intersection>
<intersection>460 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446,-486,446,-473</points>
<intersection>-486 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446,-481.5,450,-481.5</points>
<connection>
<GID>3471</GID>
<name>IN_0</name></connection>
<intersection>446 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444,-473,446,-473</points>
<connection>
<GID>3473</GID>
<name>OUT_0</name></connection>
<intersection>446 2</intersection></hsegment></shape></wire>
<wire>
<ID>4032</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,451.5,300.5,451.5</points>
<connection>
<GID>5674</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5672</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2489</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487.5,-482.5,489.5,-482.5</points>
<connection>
<GID>3474</GID>
<name>OUT</name></connection>
<connection>
<GID>3475</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288.5,448.5,302.5,448.5</points>
<connection>
<GID>5674</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288.5,448.5,288.5,461</points>
<intersection>448.5 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,452.5,292.5,452.5</points>
<connection>
<GID>5672</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,461,288.5,461</points>
<connection>
<GID>5676</GID>
<name>OUT_0</name></connection>
<intersection>288.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2490</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-485.5,491.5,-485.5</points>
<connection>
<GID>3475</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477.5,-485.5,477.5,-473</points>
<intersection>-485.5 1</intersection>
<intersection>-481.5 4</intersection>
<intersection>-473 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477.5,-481.5,481.5,-481.5</points>
<connection>
<GID>3474</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475,-473,477.5,-473</points>
<connection>
<GID>3476</GID>
<name>OUT_0</name></connection>
<intersection>477.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4034</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329,451.5,331,451.5</points>
<connection>
<GID>5680</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5678</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-507.5,468,-507.5</points>
<connection>
<GID>3503</GID>
<name>OUT</name></connection>
<connection>
<GID>3428</GID>
<name>clock</name></connection>
<connection>
<GID>3425</GID>
<name>clock</name></connection>
<connection>
<GID>3422</GID>
<name>clock</name></connection>
<connection>
<GID>3419</GID>
<name>clock</name></connection>
<connection>
<GID>3416</GID>
<name>clock</name></connection>
<connection>
<GID>3413</GID>
<name>clock</name></connection>
<connection>
<GID>3410</GID>
<name>clock</name></connection>
<connection>
<GID>3407</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,448,333,448.5</points>
<connection>
<GID>5680</GID>
<name>IN_0</name></connection>
<intersection>448 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,448,333,448</points>
<intersection>319 2</intersection>
<intersection>333 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319,448,319,461</points>
<intersection>448 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,452.5,323,452.5</points>
<connection>
<GID>5678</GID>
<name>IN_0</name></connection>
<intersection>319 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317,461,319,461</points>
<connection>
<GID>5682</GID>
<name>OUT_0</name></connection>
<intersection>319 2</intersection></hsegment></shape></wire>
<wire>
<ID>2492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-515,480.5,-515</points>
<connection>
<GID>3405</GID>
<name>IN_1</name></connection>
<connection>
<GID>3408</GID>
<name>IN_1</name></connection>
<connection>
<GID>3411</GID>
<name>IN_1</name></connection>
<connection>
<GID>3414</GID>
<name>IN_1</name></connection>
<connection>
<GID>3417</GID>
<name>IN_1</name></connection>
<connection>
<GID>3420</GID>
<name>IN_1</name></connection>
<connection>
<GID>3423</GID>
<name>IN_1</name></connection>
<connection>
<GID>3426</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,-515,245,-512.5</points>
<connection>
<GID>3502</GID>
<name>OUT_0</name></connection>
<intersection>-515 1</intersection></vsegment></shape></wire>
<wire>
<ID>4036</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360.5,451.5,362.5,451.5</points>
<connection>
<GID>5684</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5683</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,-524.5,467.5,-524.5</points>
<connection>
<GID>3505</GID>
<name>OUT</name></connection>
<connection>
<GID>3404</GID>
<name>clock</name></connection>
<connection>
<GID>3401</GID>
<name>clock</name></connection>
<connection>
<GID>3398</GID>
<name>clock</name></connection>
<connection>
<GID>3395</GID>
<name>clock</name></connection>
<connection>
<GID>3392</GID>
<name>clock</name></connection>
<connection>
<GID>3389</GID>
<name>clock</name></connection>
<connection>
<GID>3386</GID>
<name>clock</name></connection>
<connection>
<GID>3372</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350.5,448.5,364.5,448.5</points>
<connection>
<GID>5684</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,448.5,350.5,461</points>
<intersection>448.5 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350.5,452.5,354.5,452.5</points>
<connection>
<GID>5683</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348,461,350.5,461</points>
<connection>
<GID>5685</GID>
<name>OUT_0</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-532,246,-529.5</points>
<intersection>-532 2</intersection>
<intersection>-529.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>246,-532,480,-532</points>
<connection>
<GID>3370</GID>
<name>IN_1</name></connection>
<connection>
<GID>3384</GID>
<name>IN_1</name></connection>
<connection>
<GID>3387</GID>
<name>IN_1</name></connection>
<connection>
<GID>3390</GID>
<name>IN_1</name></connection>
<connection>
<GID>3393</GID>
<name>IN_1</name></connection>
<connection>
<GID>3396</GID>
<name>IN_1</name></connection>
<connection>
<GID>3399</GID>
<name>IN_1</name></connection>
<connection>
<GID>3402</GID>
<name>IN_1</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>245,-529.5,246,-529.5</points>
<connection>
<GID>3504</GID>
<name>OUT_0</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>4038</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390,451.5,392,451.5</points>
<connection>
<GID>5687</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5686</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-541.5,281.5,-401.5</points>
<connection>
<GID>3374</GID>
<name>N_in1</name></connection>
<connection>
<GID>3382</GID>
<name>N_in0</name></connection>
<intersection>-521.5 1</intersection>
<intersection>-504.5 3</intersection>
<intersection>-488.5 4</intersection>
<intersection>-473 5</intersection>
<intersection>-456.5 6</intersection>
<intersection>-439.5 7</intersection>
<intersection>-423.5 8</intersection>
<intersection>-408 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-521.5,282.5,-521.5</points>
<connection>
<GID>3386</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-408,285,-408</points>
<connection>
<GID>3591</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281.5,-504.5,283,-504.5</points>
<connection>
<GID>3410</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>281.5,-488.5,283.5,-488.5</points>
<connection>
<GID>3434</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>281.5,-473,284,-473</points>
<connection>
<GID>3458</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>281.5,-456.5,283.5,-456.5</points>
<connection>
<GID>3516</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>281.5,-439.5,284,-439.5</points>
<connection>
<GID>3543</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>281.5,-423.5,284.5,-423.5</points>
<connection>
<GID>3567</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,448,394,448.5</points>
<connection>
<GID>5687</GID>
<name>IN_0</name></connection>
<intersection>448 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,448,394,448</points>
<intersection>380 2</intersection>
<intersection>394 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380,448,380,461</points>
<intersection>448 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,452.5,384,452.5</points>
<connection>
<GID>5686</GID>
<name>IN_0</name></connection>
<intersection>380 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378,461,380,461</points>
<connection>
<GID>5688</GID>
<name>OUT_0</name></connection>
<intersection>380 2</intersection></hsegment></shape></wire>
<wire>
<ID>2496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-541.5,313.5,-401.5</points>
<connection>
<GID>3389</GID>
<name>IN_0</name></connection>
<connection>
<GID>3375</GID>
<name>N_in1</name></connection>
<connection>
<GID>3383</GID>
<name>N_in0</name></connection>
<intersection>-504.5 9</intersection>
<intersection>-488.5 10</intersection>
<intersection>-473 7</intersection>
<intersection>-456.5 11</intersection>
<intersection>-439.5 5</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,-408,316,-408</points>
<connection>
<GID>3594</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313.5,-423.5,315.5,-423.5</points>
<connection>
<GID>3570</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>313.5,-439.5,315,-439.5</points>
<connection>
<GID>3546</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>313.5,-473,315,-473</points>
<connection>
<GID>3461</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>313.5,-504.5,314,-504.5</points>
<connection>
<GID>3413</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>313.5,-488.5,314.5,-488.5</points>
<connection>
<GID>3437</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>313.5,-456.5,314.5,-456.5</points>
<connection>
<GID>3522</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4040</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421.5,451.5,423.5,451.5</points>
<connection>
<GID>5690</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5689</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,-540.5,344.5,-401.5</points>
<connection>
<GID>3392</GID>
<name>IN_0</name></connection>
<connection>
<GID>3376</GID>
<name>N_in1</name></connection>
<connection>
<GID>3477</GID>
<name>N_in0</name></connection>
<intersection>-504.5 38</intersection>
<intersection>-488.5 21</intersection>
<intersection>-473 7</intersection>
<intersection>-456.5 20</intersection>
<intersection>-439.5 5</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,-408,347,-408</points>
<connection>
<GID>3597</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>344.5,-423.5,346.5,-423.5</points>
<connection>
<GID>3573</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>344.5,-439.5,346,-439.5</points>
<connection>
<GID>3549</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>344.5,-473,346,-473</points>
<connection>
<GID>3464</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>344.5,-456.5,345.5,-456.5</points>
<connection>
<GID>3525</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>344.5,-488.5,345.5,-488.5</points>
<connection>
<GID>3440</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>344.5,-504.5,345,-504.5</points>
<connection>
<GID>3416</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411.5,448.5,425.5,448.5</points>
<connection>
<GID>5690</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411.5,448.5,411.5,461</points>
<intersection>448.5 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411.5,452.5,415.5,452.5</points>
<connection>
<GID>5689</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409,461,411.5,461</points>
<connection>
<GID>5691</GID>
<name>OUT_0</name></connection>
<intersection>411.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-504.5,375.5,-402</points>
<connection>
<GID>3528</GID>
<name>IN_0</name></connection>
<connection>
<GID>3443</GID>
<name>IN_0</name></connection>
<connection>
<GID>3478</GID>
<name>N_in0</name></connection>
<intersection>-504.5 9</intersection>
<intersection>-473 7</intersection>
<intersection>-439.5 5</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-408,377,-408</points>
<connection>
<GID>3600</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-423.5,376.5,-423.5</points>
<connection>
<GID>3576</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>375.5,-439.5,376,-439.5</points>
<connection>
<GID>3552</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>375.5,-473,376,-473</points>
<connection>
<GID>3467</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>374.5,-504.5,375.5,-504.5</points>
<connection>
<GID>3419</GID>
<name>IN_0</name></connection>
<intersection>374.5 10</intersection>
<intersection>375.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>374.5,-539.5,374.5,-504.5</points>
<connection>
<GID>3395</GID>
<name>IN_0</name></connection>
<connection>
<GID>3377</GID>
<name>N_in1</name></connection>
<intersection>-504.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>4042</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452,451.5,454,451.5</points>
<connection>
<GID>5693</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5692</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405.5,-539,405.5,-401.5</points>
<connection>
<GID>3398</GID>
<name>IN_0</name></connection>
<connection>
<GID>3378</GID>
<name>N_in1</name></connection>
<connection>
<GID>3479</GID>
<name>N_in0</name></connection>
<intersection>-504.5 13</intersection>
<intersection>-488.5 11</intersection>
<intersection>-473 9</intersection>
<intersection>-456.5 7</intersection>
<intersection>-439.5 5</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>405.5,-408,408,-408</points>
<connection>
<GID>3603</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>405.5,-423.5,407.5,-423.5</points>
<connection>
<GID>3579</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>405.5,-439.5,407,-439.5</points>
<connection>
<GID>3555</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>405.5,-456.5,406.5,-456.5</points>
<connection>
<GID>3531</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>405.5,-473,407,-473</points>
<connection>
<GID>3470</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>405.5,-488.5,406.5,-488.5</points>
<connection>
<GID>3446</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>405.5,-504.5,406,-504.5</points>
<connection>
<GID>3422</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,448,456,448.5</points>
<connection>
<GID>5693</GID>
<name>IN_0</name></connection>
<intersection>448 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,448,456,448</points>
<intersection>442 2</intersection>
<intersection>456 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442,448,442,461</points>
<intersection>448 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442,452.5,446,452.5</points>
<connection>
<GID>5692</GID>
<name>IN_0</name></connection>
<intersection>442 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,461,442,461</points>
<connection>
<GID>5694</GID>
<name>OUT_0</name></connection>
<intersection>442 2</intersection></hsegment></shape></wire>
<wire>
<ID>2500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,-538,436.5,-401.5</points>
<connection>
<GID>3401</GID>
<name>IN_0</name></connection>
<connection>
<GID>3380</GID>
<name>N_in1</name></connection>
<connection>
<GID>3480</GID>
<name>N_in0</name></connection>
<intersection>-504.5 13</intersection>
<intersection>-488.5 11</intersection>
<intersection>-473 9</intersection>
<intersection>-456.5 7</intersection>
<intersection>-439.5 5</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,-408,439,-408</points>
<connection>
<GID>3606</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436.5,-423.5,438.5,-423.5</points>
<connection>
<GID>3582</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>436.5,-439.5,438,-439.5</points>
<connection>
<GID>3558</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>436.5,-456.5,437.5,-456.5</points>
<connection>
<GID>3534</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>436.5,-473,438,-473</points>
<connection>
<GID>3473</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>436.5,-488.5,437.5,-488.5</points>
<connection>
<GID>3449</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>436.5,-504.5,437,-504.5</points>
<connection>
<GID>3425</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4044</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483.5,451.5,485.5,451.5</points>
<connection>
<GID>5696</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5695</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467.5,-540,467.5,-402</points>
<connection>
<GID>3404</GID>
<name>IN_0</name></connection>
<connection>
<GID>3379</GID>
<name>N_in1</name></connection>
<connection>
<GID>3481</GID>
<name>N_in0</name></connection>
<intersection>-504.5 13</intersection>
<intersection>-488.5 10</intersection>
<intersection>-473 8</intersection>
<intersection>-456.5 6</intersection>
<intersection>-439.5 4</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467.5,-408,470,-408</points>
<connection>
<GID>3609</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>467.5,-423.5,469.5,-423.5</points>
<connection>
<GID>3585</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>467.5,-439.5,469,-439.5</points>
<connection>
<GID>3561</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>467.5,-456.5,468.5,-456.5</points>
<connection>
<GID>3537</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>467.5,-473,469,-473</points>
<connection>
<GID>3476</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>467.5,-488.5,468.5,-488.5</points>
<connection>
<GID>3452</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>467.5,-504.5,468,-504.5</points>
<connection>
<GID>3428</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473.5,448.5,487.5,448.5</points>
<connection>
<GID>5696</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473.5,448.5,473.5,461</points>
<intersection>448.5 1</intersection>
<intersection>452.5 4</intersection>
<intersection>461 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473.5,452.5,477.5,452.5</points>
<connection>
<GID>5695</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471,461,473.5,461</points>
<connection>
<GID>5697</GID>
<name>OUT_0</name></connection>
<intersection>473.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-549.5,279.5,-394.5</points>
<connection>
<GID>3483</GID>
<name>N_in1</name></connection>
<connection>
<GID>3482</GID>
<name>N_in0</name></connection>
<intersection>-526.5 13</intersection>
<intersection>-509.5 12</intersection>
<intersection>-493.5 11</intersection>
<intersection>-478 10</intersection>
<intersection>-461.5 9</intersection>
<intersection>-444.5 8</intersection>
<intersection>-428.5 7</intersection>
<intersection>-413 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>276,-413,279.5,-413</points>
<intersection>276 23</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>275.5,-428.5,279.5,-428.5</points>
<intersection>275.5 22</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>275,-444.5,279.5,-444.5</points>
<intersection>275 21</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>274.5,-461.5,279.5,-461.5</points>
<intersection>274.5 20</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>275,-478,279.5,-478</points>
<intersection>275 17</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>274.5,-493.5,279.5,-493.5</points>
<intersection>274.5 16</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>274,-509.5,279.5,-509.5</points>
<intersection>274 15</intersection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>273.5,-526.5,279.5,-526.5</points>
<intersection>273.5 14</intersection>
<intersection>279.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>273.5,-528.5,273.5,-526.5</points>
<connection>
<GID>3371</GID>
<name>OUT_0</name></connection>
<intersection>-526.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>274,-511.5,274,-509.5</points>
<connection>
<GID>3406</GID>
<name>OUT_0</name></connection>
<intersection>-509.5 12</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>274.5,-495.5,274.5,-493.5</points>
<connection>
<GID>3430</GID>
<name>OUT_0</name></connection>
<intersection>-493.5 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>275,-480,275,-478</points>
<connection>
<GID>3454</GID>
<name>OUT_0</name></connection>
<intersection>-478 10</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>274.5,-463.5,274.5,-461.5</points>
<connection>
<GID>3507</GID>
<name>OUT_0</name></connection>
<intersection>-461.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>275,-446.5,275,-444.5</points>
<connection>
<GID>3539</GID>
<name>OUT_0</name></connection>
<intersection>-444.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>275.5,-430.5,275.5,-428.5</points>
<connection>
<GID>3563</GID>
<name>OUT_0</name></connection>
<intersection>-428.5 7</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>276,-415,276,-413</points>
<connection>
<GID>3587</GID>
<name>OUT_0</name></connection>
<intersection>-413 6</intersection></vsegment></shape></wire>
<wire>
<ID>4046</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267.5,468.5,269.5,468.5</points>
<connection>
<GID>5699</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5698</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-528.5,310.5,-394.5</points>
<connection>
<GID>3496</GID>
<name>N_in0</name></connection>
<intersection>-528.5 13</intersection>
<intersection>-511.5 12</intersection>
<intersection>-495.5 11</intersection>
<intersection>-480 10</intersection>
<intersection>-463.5 9</intersection>
<intersection>-446.5 8</intersection>
<intersection>-430.5 7</intersection>
<intersection>-415 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>307.5,-415,310.5,-415</points>
<connection>
<GID>3590</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>307,-430.5,310.5,-430.5</points>
<connection>
<GID>3566</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>306.5,-446.5,310.5,-446.5</points>
<connection>
<GID>3542</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>306,-463.5,310.5,-463.5</points>
<connection>
<GID>3514</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>306.5,-480,310.5,-480</points>
<connection>
<GID>3457</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>306,-495.5,310.5,-495.5</points>
<connection>
<GID>3433</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>305.5,-511.5,310.5,-511.5</points>
<connection>
<GID>3409</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>305,-528.5,310.5,-528.5</points>
<connection>
<GID>3385</GID>
<name>OUT_0</name></connection>
<intersection>308.5 22</intersection>
<intersection>310.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>308.5,-553,308.5,-528.5</points>
<intersection>-553 23</intersection>
<intersection>-528.5 13</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>306,-553,308.5,-553</points>
<connection>
<GID>5783</GID>
<name>N_in1</name></connection>
<intersection>308.5 22</intersection></hsegment></shape></wire>
<wire>
<ID>4047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,465,271.5,465.5</points>
<connection>
<GID>5699</GID>
<name>IN_0</name></connection>
<intersection>465 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,465,271.5,465</points>
<intersection>257.5 2</intersection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257.5,465,257.5,478</points>
<intersection>465 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257.5,469.5,261.5,469.5</points>
<connection>
<GID>5698</GID>
<name>IN_0</name></connection>
<intersection>257.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255.5,478,257.5,478</points>
<connection>
<GID>5700</GID>
<name>OUT_0</name></connection>
<intersection>257.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342.5,-548.5,342.5,-394.5</points>
<connection>
<GID>3484</GID>
<name>N_in1</name></connection>
<connection>
<GID>3495</GID>
<name>N_in0</name></connection>
<intersection>-528.5 13</intersection>
<intersection>-511.5 12</intersection>
<intersection>-495.5 11</intersection>
<intersection>-480 10</intersection>
<intersection>-463.5 9</intersection>
<intersection>-446.5 8</intersection>
<intersection>-430.5 7</intersection>
<intersection>-415 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>338,-415,342.5,-415</points>
<connection>
<GID>3593</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>337.5,-430.5,342.5,-430.5</points>
<connection>
<GID>3569</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>337,-446.5,342.5,-446.5</points>
<connection>
<GID>3545</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>336.5,-463.5,342.5,-463.5</points>
<connection>
<GID>3520</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>337,-480,342.5,-480</points>
<connection>
<GID>3460</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>336.5,-495.5,342.5,-495.5</points>
<connection>
<GID>3436</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>336,-511.5,342.5,-511.5</points>
<connection>
<GID>3412</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>335.5,-528.5,342.5,-528.5</points>
<connection>
<GID>3388</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4048</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299,468.5,301,468.5</points>
<connection>
<GID>5702</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5701</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,-548,373,-394.5</points>
<connection>
<GID>3485</GID>
<name>N_in1</name></connection>
<connection>
<GID>3494</GID>
<name>N_in0</name></connection>
<intersection>-528.5 18</intersection>
<intersection>-511.5 17</intersection>
<intersection>-495.5 16</intersection>
<intersection>-480 15</intersection>
<intersection>-463.5 14</intersection>
<intersection>-446.5 13</intersection>
<intersection>-430.5 12</intersection>
<intersection>-415 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>369.5,-415,373,-415</points>
<connection>
<GID>3596</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>369,-430.5,373,-430.5</points>
<connection>
<GID>3572</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>368.5,-446.5,373,-446.5</points>
<connection>
<GID>3548</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>368,-463.5,373,-463.5</points>
<connection>
<GID>3524</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>368.5,-480,373,-480</points>
<connection>
<GID>3463</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>368,-495.5,373,-495.5</points>
<connection>
<GID>3439</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>367.5,-511.5,373,-511.5</points>
<connection>
<GID>3415</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>367,-528.5,373,-528.5</points>
<connection>
<GID>3391</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment></shape></wire>
<wire>
<ID>4049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,465.5,303,465.5</points>
<connection>
<GID>5702</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289,465.5,289,478</points>
<intersection>465.5 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289,469.5,293,469.5</points>
<connection>
<GID>5701</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286.5,478,289,478</points>
<connection>
<GID>5703</GID>
<name>OUT_0</name></connection>
<intersection>289 2</intersection></hsegment></shape></wire>
<wire>
<ID>2506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,-548,403.5,-394.5</points>
<connection>
<GID>3486</GID>
<name>N_in1</name></connection>
<connection>
<GID>3493</GID>
<name>N_in0</name></connection>
<intersection>-528.5 9</intersection>
<intersection>-511.5 10</intersection>
<intersection>-495.5 11</intersection>
<intersection>-480 12</intersection>
<intersection>-463.5 13</intersection>
<intersection>-446.5 14</intersection>
<intersection>-430.5 15</intersection>
<intersection>-415 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>396.5,-528.5,403.5,-528.5</points>
<connection>
<GID>3394</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>397,-511.5,403.5,-511.5</points>
<connection>
<GID>3418</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>397.5,-495.5,403.5,-495.5</points>
<connection>
<GID>3442</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>398,-480,403.5,-480</points>
<connection>
<GID>3466</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>397.5,-463.5,403.5,-463.5</points>
<connection>
<GID>3527</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>398,-446.5,403.5,-446.5</points>
<connection>
<GID>3551</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>398.5,-430.5,403.5,-430.5</points>
<connection>
<GID>3575</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>399,-415,403.5,-415</points>
<connection>
<GID>3599</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4050</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329.5,468.5,331.5,468.5</points>
<connection>
<GID>5705</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5704</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-548,434.5,-394.5</points>
<connection>
<GID>3487</GID>
<name>N_in1</name></connection>
<connection>
<GID>3492</GID>
<name>N_in0</name></connection>
<intersection>-528.5 6</intersection>
<intersection>-511.5 7</intersection>
<intersection>-495.5 8</intersection>
<intersection>-480 9</intersection>
<intersection>-463.5 10</intersection>
<intersection>-446.5 11</intersection>
<intersection>-430.5 12</intersection>
<intersection>-415 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>428,-528.5,434.5,-528.5</points>
<connection>
<GID>3397</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>428.5,-511.5,434.5,-511.5</points>
<connection>
<GID>3421</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>429,-495.5,434.5,-495.5</points>
<connection>
<GID>3445</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>429.5,-480,434.5,-480</points>
<connection>
<GID>3469</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>429,-463.5,434.5,-463.5</points>
<connection>
<GID>3530</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>429.5,-446.5,434.5,-446.5</points>
<connection>
<GID>3554</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>430,-430.5,434.5,-430.5</points>
<connection>
<GID>3578</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>430.5,-415,434.5,-415</points>
<connection>
<GID>3602</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,465,333.5,465.5</points>
<connection>
<GID>5705</GID>
<name>IN_0</name></connection>
<intersection>465 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,465,333.5,465</points>
<intersection>319.5 2</intersection>
<intersection>333.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319.5,465,319.5,478</points>
<intersection>465 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319.5,469.5,323.5,469.5</points>
<connection>
<GID>5704</GID>
<name>IN_0</name></connection>
<intersection>319.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317.5,478,319.5,478</points>
<connection>
<GID>5706</GID>
<name>OUT_0</name></connection>
<intersection>319.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465.5,-548.5,465.5,-393.5</points>
<connection>
<GID>3488</GID>
<name>N_in1</name></connection>
<connection>
<GID>3491</GID>
<name>N_in0</name></connection>
<intersection>-528.5 6</intersection>
<intersection>-511.5 7</intersection>
<intersection>-495.5 8</intersection>
<intersection>-480 9</intersection>
<intersection>-463.5 10</intersection>
<intersection>-446.5 11</intersection>
<intersection>-430.5 12</intersection>
<intersection>-415 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>458.5,-528.5,465.5,-528.5</points>
<connection>
<GID>3400</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>459,-511.5,465.5,-511.5</points>
<connection>
<GID>3424</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>459.5,-495.5,465.5,-495.5</points>
<connection>
<GID>3448</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>460,-480,465.5,-480</points>
<connection>
<GID>3472</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>459.5,-463.5,465.5,-463.5</points>
<connection>
<GID>3533</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>460,-446.5,465.5,-446.5</points>
<connection>
<GID>3557</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>460.5,-430.5,465.5,-430.5</points>
<connection>
<GID>3581</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>461,-415,465.5,-415</points>
<connection>
<GID>3605</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4052</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361,468.5,363,468.5</points>
<connection>
<GID>5708</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5707</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496,-548,496,-393</points>
<connection>
<GID>3489</GID>
<name>N_in1</name></connection>
<connection>
<GID>3490</GID>
<name>N_in0</name></connection>
<intersection>-528.5 3</intersection>
<intersection>-511.5 4</intersection>
<intersection>-495.5 5</intersection>
<intersection>-480 6</intersection>
<intersection>-463.5 7</intersection>
<intersection>-446.5 8</intersection>
<intersection>-430.5 9</intersection>
<intersection>-415 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>490,-528.5,496,-528.5</points>
<connection>
<GID>3403</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>490.5,-511.5,496,-511.5</points>
<connection>
<GID>3427</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>491,-495.5,496,-495.5</points>
<connection>
<GID>3451</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>491.5,-480,496,-480</points>
<connection>
<GID>3475</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>491,-463.5,496,-463.5</points>
<connection>
<GID>3536</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>491.5,-446.5,496,-446.5</points>
<connection>
<GID>3560</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>492,-430.5,496,-430.5</points>
<connection>
<GID>3584</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>492.5,-415,496,-415</points>
<connection>
<GID>3608</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment></shape></wire>
<wire>
<ID>4053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351,465.5,365,465.5</points>
<connection>
<GID>5708</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351,465.5,351,478</points>
<intersection>465.5 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351,469.5,355,469.5</points>
<connection>
<GID>5707</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348.5,478,351,478</points>
<connection>
<GID>5709</GID>
<name>OUT_0</name></connection>
<intersection>351 2</intersection></hsegment></shape></wire>
<wire>
<ID>2510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-462.5,204.5,-413.5</points>
<intersection>-462.5 2</intersection>
<intersection>-413.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-413.5,243.5,-413.5</points>
<connection>
<GID>3509</GID>
<name>ENABLE_0</name></connection>
<intersection>204.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-462.5,204.5,-462.5</points>
<connection>
<GID>3497</GID>
<name>OUT_7</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-413.5,229.5,-410</points>
<intersection>-413.5 1</intersection>
<intersection>-410 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-410,234,-410</points>
<connection>
<GID>3510</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4054</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390.5,468.5,392.5,468.5</points>
<connection>
<GID>5711</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5710</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-463.5,206.5,-429</points>
<intersection>-463.5 2</intersection>
<intersection>-429 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,-429,243.5,-429</points>
<intersection>206.5 0</intersection>
<intersection>229.5 4</intersection>
<intersection>243.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-463.5,206.5,-463.5</points>
<connection>
<GID>3497</GID>
<name>OUT_6</name></connection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243.5,-429.5,243.5,-429</points>
<connection>
<GID>3511</GID>
<name>ENABLE_0</name></connection>
<intersection>-429 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-429,229.5,-425.5</points>
<intersection>-429 1</intersection>
<intersection>-425.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-425.5,233.5,-425.5</points>
<connection>
<GID>3513</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,465,394.5,465.5</points>
<connection>
<GID>5711</GID>
<name>IN_0</name></connection>
<intersection>465 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,465,394.5,465</points>
<intersection>380.5 2</intersection>
<intersection>394.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380.5,465,380.5,478</points>
<intersection>465 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380.5,469.5,384.5,469.5</points>
<connection>
<GID>5710</GID>
<name>IN_0</name></connection>
<intersection>380.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378.5,478,380.5,478</points>
<connection>
<GID>5712</GID>
<name>OUT_0</name></connection>
<intersection>380.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-464.5,208.5,-441.5</points>
<intersection>-464.5 2</intersection>
<intersection>-441.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-441.5,233.5,-441.5</points>
<connection>
<GID>3517</GID>
<name>IN_0</name></connection>
<intersection>208.5 0</intersection>
<intersection>229.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-464.5,208.5,-464.5</points>
<connection>
<GID>3497</GID>
<name>OUT_5</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229.5,-445.5,229.5,-441.5</points>
<intersection>-445.5 4</intersection>
<intersection>-441.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229.5,-445.5,243.5,-445.5</points>
<connection>
<GID>3515</GID>
<name>ENABLE_0</name></connection>
<intersection>229.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>4056</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422,468.5,424,468.5</points>
<connection>
<GID>5714</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5713</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,-465.5,210.5,-458.5</points>
<intersection>-465.5 2</intersection>
<intersection>-458.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,-458.5,233.5,-458.5</points>
<connection>
<GID>3521</GID>
<name>IN_0</name></connection>
<intersection>210.5 0</intersection>
<intersection>229.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-465.5,210.5,-465.5</points>
<connection>
<GID>3497</GID>
<name>OUT_4</name></connection>
<intersection>210.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229.5,-462.5,229.5,-458.5</points>
<intersection>-462.5 4</intersection>
<intersection>-458.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229.5,-462.5,243.5,-462.5</points>
<connection>
<GID>3519</GID>
<name>ENABLE_0</name></connection>
<intersection>229.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>4057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,465.5,426,465.5</points>
<connection>
<GID>5714</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412,465.5,412,478</points>
<intersection>465.5 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412,469.5,416,469.5</points>
<connection>
<GID>5713</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409.5,478,412,478</points>
<connection>
<GID>5715</GID>
<name>OUT_0</name></connection>
<intersection>412 2</intersection></hsegment></shape></wire>
<wire>
<ID>2514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,-478.5,210.5,-466.5</points>
<intersection>-478.5 1</intersection>
<intersection>-466.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,-478.5,242.5,-478.5</points>
<connection>
<GID>3498</GID>
<name>ENABLE_0</name></connection>
<intersection>210.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-466.5,210.5,-466.5</points>
<connection>
<GID>3497</GID>
<name>OUT_3</name></connection>
<intersection>210.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-478.5,229.5,-475</points>
<intersection>-478.5 1</intersection>
<intersection>-475 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-475,233.5,-475</points>
<connection>
<GID>3499</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4058</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452.5,468.5,454.5,468.5</points>
<connection>
<GID>5717</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5716</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-494.5,208.5,-467.5</points>
<intersection>-494.5 1</intersection>
<intersection>-467.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-494.5,242.5,-494.5</points>
<connection>
<GID>3500</GID>
<name>ENABLE_0</name></connection>
<intersection>208.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-467.5,208.5,-467.5</points>
<connection>
<GID>3497</GID>
<name>OUT_2</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-494.5,229.5,-490.5</points>
<intersection>-494.5 1</intersection>
<intersection>-490.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-490.5,233.5,-490.5</points>
<connection>
<GID>3501</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,465,456.5,465.5</points>
<connection>
<GID>5717</GID>
<name>IN_0</name></connection>
<intersection>465 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,465,456.5,465</points>
<intersection>442.5 2</intersection>
<intersection>456.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442.5,465,442.5,478</points>
<intersection>465 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442.5,469.5,446.5,469.5</points>
<connection>
<GID>5716</GID>
<name>IN_0</name></connection>
<intersection>442.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,478,442.5,478</points>
<connection>
<GID>5718</GID>
<name>OUT_0</name></connection>
<intersection>442.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-510,206.5,-468.5</points>
<intersection>-510 1</intersection>
<intersection>-468.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,-510,242.5,-510</points>
<intersection>206.5 0</intersection>
<intersection>229.5 4</intersection>
<intersection>242.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-468.5,206.5,-468.5</points>
<connection>
<GID>3497</GID>
<name>OUT_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,-510.5,242.5,-510</points>
<connection>
<GID>3502</GID>
<name>ENABLE_0</name></connection>
<intersection>-510 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-510,229.5,-506.5</points>
<intersection>-510 1</intersection>
<intersection>-506.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-506.5,233.5,-506.5</points>
<connection>
<GID>3503</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4060</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484,468.5,486,468.5</points>
<connection>
<GID>5720</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5719</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-527.5,204.5,-469.5</points>
<intersection>-527.5 1</intersection>
<intersection>-469.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-527.5,242.5,-527.5</points>
<connection>
<GID>3504</GID>
<name>ENABLE_0</name></connection>
<intersection>204.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-469.5,204.5,-469.5</points>
<connection>
<GID>3497</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,-527.5,229.5,-523.5</points>
<intersection>-527.5 1</intersection>
<intersection>-523.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-523.5,233.5,-523.5</points>
<connection>
<GID>3505</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>4061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474,465.5,488,465.5</points>
<connection>
<GID>5720</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474,465.5,474,478</points>
<intersection>465.5 1</intersection>
<intersection>469.5 4</intersection>
<intersection>478 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474,469.5,478,469.5</points>
<connection>
<GID>5719</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471.5,478,474,478</points>
<connection>
<GID>5721</GID>
<name>OUT_0</name></connection>
<intersection>474 2</intersection></hsegment></shape></wire>
<wire>
<ID>2518</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270.5,-466,272.5,-466</points>
<connection>
<GID>3506</GID>
<name>OUT</name></connection>
<connection>
<GID>3507</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4062</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268,484.5,270,484.5</points>
<connection>
<GID>5723</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5722</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-469.5,274.5,-469</points>
<connection>
<GID>3507</GID>
<name>IN_0</name></connection>
<intersection>-469.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,-469.5,274.5,-469.5</points>
<intersection>260.5 2</intersection>
<intersection>274.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260.5,-469.5,260.5,-456.5</points>
<intersection>-469.5 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,-465,264.5,-465</points>
<connection>
<GID>3506</GID>
<name>IN_0</name></connection>
<intersection>260.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258.5,-456.5,260.5,-456.5</points>
<connection>
<GID>3508</GID>
<name>OUT_0</name></connection>
<intersection>260.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4063</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,481,272,481.5</points>
<connection>
<GID>5723</GID>
<name>IN_0</name></connection>
<intersection>481 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,481,272,481</points>
<intersection>258 2</intersection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,481,258,494</points>
<intersection>481 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258,485.5,262,485.5</points>
<connection>
<GID>5722</GID>
<name>IN_0</name></connection>
<intersection>258 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256,494,258,494</points>
<connection>
<GID>5724</GID>
<name>OUT_0</name></connection>
<intersection>258 2</intersection></hsegment></shape></wire>
<wire>
<ID>2520</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302,-466,304,-466</points>
<connection>
<GID>3512</GID>
<name>OUT</name></connection>
<connection>
<GID>3514</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4064</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299.5,484.5,301.5,484.5</points>
<connection>
<GID>5726</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5725</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,-469,306,-469</points>
<connection>
<GID>3514</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292,-469,292,-456.5</points>
<intersection>-469 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292,-465,296,-465</points>
<connection>
<GID>3512</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289.5,-456.5,292,-456.5</points>
<connection>
<GID>3516</GID>
<name>OUT_0</name></connection>
<intersection>292 2</intersection></hsegment></shape></wire>
<wire>
<ID>4065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,481.5,303.5,481.5</points>
<connection>
<GID>5726</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289.5,481.5,289.5,494</points>
<intersection>481.5 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289.5,485.5,293.5,485.5</points>
<connection>
<GID>5725</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287,494,289.5,494</points>
<connection>
<GID>5727</GID>
<name>OUT_0</name></connection>
<intersection>289.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2522</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332.5,-466,334.5,-466</points>
<connection>
<GID>3518</GID>
<name>OUT</name></connection>
<connection>
<GID>3520</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4066</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330,484.5,332,484.5</points>
<connection>
<GID>5729</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5728</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,-469.5,336.5,-469</points>
<connection>
<GID>3520</GID>
<name>IN_0</name></connection>
<intersection>-469.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,-469.5,336.5,-469.5</points>
<intersection>322.5 2</intersection>
<intersection>336.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322.5,-469.5,322.5,-456.5</points>
<intersection>-469.5 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322.5,-465,326.5,-465</points>
<connection>
<GID>3518</GID>
<name>IN_0</name></connection>
<intersection>322.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320.5,-456.5,322.5,-456.5</points>
<connection>
<GID>3522</GID>
<name>OUT_0</name></connection>
<intersection>322.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4067</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,481,334,481.5</points>
<connection>
<GID>5729</GID>
<name>IN_0</name></connection>
<intersection>481 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,481,334,481</points>
<intersection>320 2</intersection>
<intersection>334 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320,481,320,494</points>
<intersection>481 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320,485.5,324,485.5</points>
<connection>
<GID>5728</GID>
<name>IN_0</name></connection>
<intersection>320 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318,494,320,494</points>
<connection>
<GID>5730</GID>
<name>OUT_0</name></connection>
<intersection>320 2</intersection></hsegment></shape></wire>
<wire>
<ID>2524</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364,-466,366,-466</points>
<connection>
<GID>3523</GID>
<name>OUT</name></connection>
<connection>
<GID>3524</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4068</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361.5,484.5,363.5,484.5</points>
<connection>
<GID>5732</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5731</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354,-469,368,-469</points>
<connection>
<GID>3524</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354,-469,354,-456.5</points>
<intersection>-469 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354,-465,358,-465</points>
<connection>
<GID>3523</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351.5,-456.5,354,-456.5</points>
<connection>
<GID>3525</GID>
<name>OUT_0</name></connection>
<intersection>354 2</intersection></hsegment></shape></wire>
<wire>
<ID>4069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351.5,481.5,365.5,481.5</points>
<connection>
<GID>5732</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351.5,481.5,351.5,494</points>
<intersection>481.5 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351.5,485.5,355.5,485.5</points>
<connection>
<GID>5731</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>349,494,351.5,494</points>
<connection>
<GID>5733</GID>
<name>OUT_0</name></connection>
<intersection>351.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2526</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393.5,-466,395.5,-466</points>
<connection>
<GID>3526</GID>
<name>OUT</name></connection>
<connection>
<GID>3527</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4070</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391,484.5,393,484.5</points>
<connection>
<GID>5735</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5734</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,-469.5,397.5,-469</points>
<connection>
<GID>3527</GID>
<name>IN_0</name></connection>
<intersection>-469.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,-469.5,397.5,-469.5</points>
<intersection>383.5 2</intersection>
<intersection>397.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,-469.5,383.5,-456.5</points>
<intersection>-469.5 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383.5,-465,387.5,-465</points>
<connection>
<GID>3526</GID>
<name>IN_0</name></connection>
<intersection>383.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381.5,-456.5,383.5,-456.5</points>
<connection>
<GID>3528</GID>
<name>OUT_0</name></connection>
<intersection>383.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395,481,395,481.5</points>
<connection>
<GID>5735</GID>
<name>IN_0</name></connection>
<intersection>481 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,481,395,481</points>
<intersection>381 2</intersection>
<intersection>395 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381,481,381,494</points>
<intersection>481 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381,485.5,385,485.5</points>
<connection>
<GID>5734</GID>
<name>IN_0</name></connection>
<intersection>381 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379,494,381,494</points>
<connection>
<GID>5736</GID>
<name>OUT_0</name></connection>
<intersection>381 2</intersection></hsegment></shape></wire>
<wire>
<ID>2528</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425,-466,427,-466</points>
<connection>
<GID>3529</GID>
<name>OUT</name></connection>
<connection>
<GID>3530</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4072</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422.5,484.5,424.5,484.5</points>
<connection>
<GID>5738</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5737</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415,-469,429,-469</points>
<connection>
<GID>3530</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415,-469,415,-456.5</points>
<intersection>-469 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415,-465,419,-465</points>
<connection>
<GID>3529</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412.5,-456.5,415,-456.5</points>
<connection>
<GID>3531</GID>
<name>OUT_0</name></connection>
<intersection>415 2</intersection></hsegment></shape></wire>
<wire>
<ID>4073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,481.5,426.5,481.5</points>
<connection>
<GID>5738</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412.5,481.5,412.5,494</points>
<intersection>481.5 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412.5,485.5,416.5,485.5</points>
<connection>
<GID>5737</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410,494,412.5,494</points>
<connection>
<GID>5739</GID>
<name>OUT_0</name></connection>
<intersection>412.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2530</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455.5,-466,457.5,-466</points>
<connection>
<GID>3532</GID>
<name>OUT</name></connection>
<connection>
<GID>3533</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4074</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453,484.5,455,484.5</points>
<connection>
<GID>5741</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5740</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-469.5,459.5,-469</points>
<connection>
<GID>3533</GID>
<name>IN_0</name></connection>
<intersection>-469.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,-469.5,459.5,-469.5</points>
<intersection>445.5 2</intersection>
<intersection>459.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445.5,-469.5,445.5,-456.5</points>
<intersection>-469.5 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445.5,-465,449.5,-465</points>
<connection>
<GID>3532</GID>
<name>IN_0</name></connection>
<intersection>445.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443.5,-456.5,445.5,-456.5</points>
<connection>
<GID>3534</GID>
<name>OUT_0</name></connection>
<intersection>445.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,481,457,481.5</points>
<connection>
<GID>5741</GID>
<name>IN_0</name></connection>
<intersection>481 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443,481,457,481</points>
<intersection>443 2</intersection>
<intersection>457 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443,481,443,494</points>
<intersection>481 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443,485.5,447,485.5</points>
<connection>
<GID>5740</GID>
<name>IN_0</name></connection>
<intersection>443 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441,494,443,494</points>
<connection>
<GID>5742</GID>
<name>OUT_0</name></connection>
<intersection>443 2</intersection></hsegment></shape></wire>
<wire>
<ID>2532</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487,-466,489,-466</points>
<connection>
<GID>3535</GID>
<name>OUT</name></connection>
<connection>
<GID>3536</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4076</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484.5,484.5,486.5,484.5</points>
<connection>
<GID>5744</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5743</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,-469,491,-469</points>
<connection>
<GID>3536</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477,-469,477,-456.5</points>
<intersection>-469 1</intersection>
<intersection>-465 4</intersection>
<intersection>-456.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477,-465,481,-465</points>
<connection>
<GID>3535</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474.5,-456.5,477,-456.5</points>
<connection>
<GID>3537</GID>
<name>OUT_0</name></connection>
<intersection>477 2</intersection></hsegment></shape></wire>
<wire>
<ID>4077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474.5,481.5,488.5,481.5</points>
<connection>
<GID>5744</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474.5,481.5,474.5,494</points>
<intersection>481.5 1</intersection>
<intersection>485.5 4</intersection>
<intersection>494 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474.5,485.5,478.5,485.5</points>
<connection>
<GID>5743</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472,494,474.5,494</points>
<connection>
<GID>5745</GID>
<name>OUT_0</name></connection>
<intersection>474.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2534</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271,-449,273,-449</points>
<connection>
<GID>3538</GID>
<name>OUT</name></connection>
<connection>
<GID>3539</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4078</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268.5,500,270.5,500</points>
<connection>
<GID>5747</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5746</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-452.5,275,-452</points>
<connection>
<GID>3539</GID>
<name>IN_0</name></connection>
<intersection>-452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-452.5,275,-452.5</points>
<intersection>261 2</intersection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261,-452.5,261,-439.5</points>
<intersection>-452.5 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,-448,265,-448</points>
<connection>
<GID>3538</GID>
<name>IN_0</name></connection>
<intersection>261 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259,-439.5,261,-439.5</points>
<connection>
<GID>3540</GID>
<name>OUT_0</name></connection>
<intersection>261 2</intersection></hsegment></shape></wire>
<wire>
<ID>4079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,496.5,272.5,497</points>
<connection>
<GID>5747</GID>
<name>IN_0</name></connection>
<intersection>496.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258.5,496.5,272.5,496.5</points>
<intersection>258.5 2</intersection>
<intersection>272.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258.5,496.5,258.5,509.5</points>
<intersection>496.5 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258.5,501,262.5,501</points>
<connection>
<GID>5746</GID>
<name>IN_0</name></connection>
<intersection>258.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256.5,509.5,258.5,509.5</points>
<connection>
<GID>5748</GID>
<name>OUT_0</name></connection>
<intersection>258.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2536</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302.5,-449,304.5,-449</points>
<connection>
<GID>3541</GID>
<name>OUT</name></connection>
<connection>
<GID>3542</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4080</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>300,500,302,500</points>
<connection>
<GID>5750</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5749</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-452,306.5,-452</points>
<connection>
<GID>3542</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292.5,-452,292.5,-439.5</points>
<intersection>-452 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292.5,-448,296.5,-448</points>
<connection>
<GID>3541</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290,-439.5,292.5,-439.5</points>
<connection>
<GID>3543</GID>
<name>OUT_0</name></connection>
<intersection>292.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4081</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,497,304,497</points>
<connection>
<GID>5750</GID>
<name>IN_0</name></connection>
<intersection>290 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>290,497,290,509.5</points>
<intersection>497 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>290,501,294,501</points>
<connection>
<GID>5749</GID>
<name>IN_0</name></connection>
<intersection>290 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287.5,509.5,290,509.5</points>
<connection>
<GID>5751</GID>
<name>OUT_0</name></connection>
<intersection>290 2</intersection></hsegment></shape></wire>
<wire>
<ID>2538</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333,-449,335,-449</points>
<connection>
<GID>3544</GID>
<name>OUT</name></connection>
<connection>
<GID>3545</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4082</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330.5,500,332.5,500</points>
<connection>
<GID>5753</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5752</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-452.5,337,-452</points>
<connection>
<GID>3545</GID>
<name>IN_0</name></connection>
<intersection>-452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,-452.5,337,-452.5</points>
<intersection>323 2</intersection>
<intersection>337 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323,-452.5,323,-439.5</points>
<intersection>-452.5 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323,-448,327,-448</points>
<connection>
<GID>3544</GID>
<name>IN_0</name></connection>
<intersection>323 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321,-439.5,323,-439.5</points>
<connection>
<GID>3546</GID>
<name>OUT_0</name></connection>
<intersection>323 2</intersection></hsegment></shape></wire>
<wire>
<ID>4083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334.5,496.5,334.5,497</points>
<connection>
<GID>5753</GID>
<name>IN_0</name></connection>
<intersection>496.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,496.5,334.5,496.5</points>
<intersection>320.5 2</intersection>
<intersection>334.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320.5,496.5,320.5,509.5</points>
<intersection>496.5 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320.5,501,324.5,501</points>
<connection>
<GID>5752</GID>
<name>IN_0</name></connection>
<intersection>320.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318.5,509.5,320.5,509.5</points>
<connection>
<GID>5754</GID>
<name>OUT_0</name></connection>
<intersection>320.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2540</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364.5,-449,366.5,-449</points>
<connection>
<GID>3547</GID>
<name>OUT</name></connection>
<connection>
<GID>3548</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4084</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>362,500,364,500</points>
<connection>
<GID>5756</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5755</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2541</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-452,368.5,-452</points>
<connection>
<GID>3548</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354.5,-452,354.5,-439.5</points>
<intersection>-452 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354.5,-448,358.5,-448</points>
<connection>
<GID>3547</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352,-439.5,354.5,-439.5</points>
<connection>
<GID>3549</GID>
<name>OUT_0</name></connection>
<intersection>354.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2542</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394,-449,396,-449</points>
<connection>
<GID>3550</GID>
<name>OUT</name></connection>
<connection>
<GID>3551</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4086</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391.5,500,393.5,500</points>
<connection>
<GID>5759</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5758</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,-452.5,398,-452</points>
<connection>
<GID>3551</GID>
<name>IN_0</name></connection>
<intersection>-452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-452.5,398,-452.5</points>
<intersection>384 2</intersection>
<intersection>398 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384,-452.5,384,-439.5</points>
<intersection>-452.5 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384,-448,388,-448</points>
<connection>
<GID>3550</GID>
<name>IN_0</name></connection>
<intersection>384 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382,-439.5,384,-439.5</points>
<connection>
<GID>3552</GID>
<name>OUT_0</name></connection>
<intersection>384 2</intersection></hsegment></shape></wire>
<wire>
<ID>4087</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395.5,496.5,395.5,497</points>
<connection>
<GID>5759</GID>
<name>IN_0</name></connection>
<intersection>496.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381.5,496.5,395.5,496.5</points>
<intersection>381.5 2</intersection>
<intersection>395.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381.5,496.5,381.5,509.5</points>
<intersection>496.5 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381.5,501,385.5,501</points>
<connection>
<GID>5758</GID>
<name>IN_0</name></connection>
<intersection>381.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379.5,509.5,381.5,509.5</points>
<connection>
<GID>5760</GID>
<name>OUT_0</name></connection>
<intersection>381.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2544</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425.5,-449,427.5,-449</points>
<connection>
<GID>3553</GID>
<name>OUT</name></connection>
<connection>
<GID>3554</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4088</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>423,500,425,500</points>
<connection>
<GID>5762</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5761</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2545</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415.5,-452,429.5,-452</points>
<connection>
<GID>3554</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415.5,-452,415.5,-439.5</points>
<intersection>-452 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415.5,-448,419.5,-448</points>
<connection>
<GID>3553</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413,-439.5,415.5,-439.5</points>
<connection>
<GID>3555</GID>
<name>OUT_0</name></connection>
<intersection>415.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413,497,427,497</points>
<connection>
<GID>5762</GID>
<name>IN_0</name></connection>
<intersection>413 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>413,497,413,509.5</points>
<intersection>497 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>413,501,417,501</points>
<connection>
<GID>5761</GID>
<name>IN_0</name></connection>
<intersection>413 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410.5,509.5,413,509.5</points>
<connection>
<GID>5763</GID>
<name>OUT_0</name></connection>
<intersection>413 2</intersection></hsegment></shape></wire>
<wire>
<ID>2546</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456,-449,458,-449</points>
<connection>
<GID>3556</GID>
<name>OUT</name></connection>
<connection>
<GID>3557</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4090</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453.5,500,455.5,500</points>
<connection>
<GID>5765</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5764</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460,-452.5,460,-452</points>
<connection>
<GID>3557</GID>
<name>IN_0</name></connection>
<intersection>-452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446,-452.5,460,-452.5</points>
<intersection>446 2</intersection>
<intersection>460 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446,-452.5,446,-439.5</points>
<intersection>-452.5 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446,-448,450,-448</points>
<connection>
<GID>3556</GID>
<name>IN_0</name></connection>
<intersection>446 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444,-439.5,446,-439.5</points>
<connection>
<GID>3558</GID>
<name>OUT_0</name></connection>
<intersection>446 2</intersection></hsegment></shape></wire>
<wire>
<ID>4091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,496.5,457.5,497</points>
<connection>
<GID>5765</GID>
<name>IN_0</name></connection>
<intersection>496.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443.5,496.5,457.5,496.5</points>
<intersection>443.5 2</intersection>
<intersection>457.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443.5,496.5,443.5,509.5</points>
<intersection>496.5 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443.5,501,447.5,501</points>
<connection>
<GID>5764</GID>
<name>IN_0</name></connection>
<intersection>443.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441.5,509.5,443.5,509.5</points>
<connection>
<GID>5766</GID>
<name>OUT_0</name></connection>
<intersection>443.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2548</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487.5,-449,489.5,-449</points>
<connection>
<GID>3559</GID>
<name>OUT</name></connection>
<connection>
<GID>3560</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4092</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>485,500,487,500</points>
<connection>
<GID>5768</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>5767</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-452,491.5,-452</points>
<connection>
<GID>3560</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477.5,-452,477.5,-439.5</points>
<intersection>-452 1</intersection>
<intersection>-448 4</intersection>
<intersection>-439.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477.5,-448,481.5,-448</points>
<connection>
<GID>3559</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475,-439.5,477.5,-439.5</points>
<connection>
<GID>3561</GID>
<name>OUT_0</name></connection>
<intersection>477.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4093</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475,497,489,497</points>
<connection>
<GID>5768</GID>
<name>IN_0</name></connection>
<intersection>475 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>475,497,475,509.5</points>
<intersection>497 1</intersection>
<intersection>501 4</intersection>
<intersection>509.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>475,501,479,501</points>
<connection>
<GID>5767</GID>
<name>IN_0</name></connection>
<intersection>475 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472.5,509.5,475,509.5</points>
<connection>
<GID>5769</GID>
<name>OUT_0</name></connection>
<intersection>475 2</intersection></hsegment></shape></wire>
<wire>
<ID>2550</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271.5,-433,273.5,-433</points>
<connection>
<GID>3562</GID>
<name>OUT</name></connection>
<connection>
<GID>3563</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,376.5,247,509.5</points>
<connection>
<GID>5533</GID>
<name>N_in1</name></connection>
<intersection>396 14</intersection>
<intersection>413 12</intersection>
<intersection>429 10</intersection>
<intersection>444.5 8</intersection>
<intersection>461 6</intersection>
<intersection>478 4</intersection>
<intersection>494 2</intersection>
<intersection>509.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,509.5,250.5,509.5</points>
<connection>
<GID>5748</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>247,494,250,494</points>
<connection>
<GID>5724</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>247,478,249.5,478</points>
<connection>
<GID>5700</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>247,461,249,461</points>
<connection>
<GID>5668</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>247,444.5,249.5,444.5</points>
<connection>
<GID>5615</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>247,429,249,429</points>
<connection>
<GID>5591</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>247,413,248.5,413</points>
<connection>
<GID>5567</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>247,396,248,396</points>
<connection>
<GID>5532</GID>
<name>IN_0</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>2551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-436.5,275.5,-436</points>
<connection>
<GID>3563</GID>
<name>IN_0</name></connection>
<intersection>-436.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-436.5,275.5,-436.5</points>
<intersection>261.5 2</intersection>
<intersection>275.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261.5,-436.5,261.5,-423.5</points>
<intersection>-436.5 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261.5,-432,265.5,-432</points>
<connection>
<GID>3562</GID>
<name>IN_0</name></connection>
<intersection>261.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259.5,-423.5,261.5,-423.5</points>
<connection>
<GID>3564</GID>
<name>OUT_0</name></connection>
<intersection>261.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4095</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242.5,499,479,499</points>
<connection>
<GID>5767</GID>
<name>IN_1</name></connection>
<connection>
<GID>5764</GID>
<name>IN_1</name></connection>
<connection>
<GID>5761</GID>
<name>IN_1</name></connection>
<connection>
<GID>5758</GID>
<name>IN_1</name></connection>
<connection>
<GID>5755</GID>
<name>IN_1</name></connection>
<connection>
<GID>5752</GID>
<name>IN_1</name></connection>
<connection>
<GID>5749</GID>
<name>IN_1</name></connection>
<connection>
<GID>5746</GID>
<name>IN_1</name></connection>
<intersection>242.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,499,242.5,502</points>
<connection>
<GID>5669</GID>
<name>OUT_0</name></connection>
<intersection>499 1</intersection></vsegment></shape></wire>
<wire>
<ID>2552</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>303,-433,305,-433</points>
<connection>
<GID>3565</GID>
<name>OUT</name></connection>
<connection>
<GID>3566</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4096</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,506.5,466.5,506.5</points>
<connection>
<GID>5769</GID>
<name>clock</name></connection>
<connection>
<GID>5766</GID>
<name>clock</name></connection>
<connection>
<GID>5763</GID>
<name>clock</name></connection>
<connection>
<GID>5760</GID>
<name>clock</name></connection>
<connection>
<GID>5757</GID>
<name>clock</name></connection>
<connection>
<GID>5754</GID>
<name>clock</name></connection>
<connection>
<GID>5751</GID>
<name>clock</name></connection>
<connection>
<GID>5748</GID>
<name>clock</name></connection>
<connection>
<GID>5670</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2553</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293,-436,307,-436</points>
<connection>
<GID>3566</GID>
<name>IN_0</name></connection>
<intersection>293 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>293,-436,293,-423.5</points>
<intersection>-436 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>293,-432,297,-432</points>
<connection>
<GID>3565</GID>
<name>IN_0</name></connection>
<intersection>293 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290.5,-423.5,293,-423.5</points>
<connection>
<GID>3567</GID>
<name>OUT_0</name></connection>
<intersection>293 2</intersection></hsegment></shape></wire>
<wire>
<ID>4097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,334.5,245.5,354.5</points>
<connection>
<GID>4821</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>247,354.5,247,374.5</points>
<connection>
<GID>5533</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>245.5,354.5,247,354.5</points>
<intersection>245.5 0</intersection>
<intersection>247 1</intersection></hsegment></shape></wire>
<wire>
<ID>2554</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333.5,-433,335.5,-433</points>
<connection>
<GID>3568</GID>
<name>OUT</name></connection>
<connection>
<GID>3569</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,341.5,274.5,353.5</points>
<connection>
<GID>4922</GID>
<name>N_in1</name></connection>
<intersection>353.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>276,353.5,276,366</points>
<connection>
<GID>5643</GID>
<name>N_in0</name></connection>
<intersection>353.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>274.5,353.5,276,353.5</points>
<intersection>274.5 0</intersection>
<intersection>276 1</intersection></hsegment></shape></wire>
<wire>
<ID>2555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,-436.5,337.5,-436</points>
<connection>
<GID>3569</GID>
<name>IN_0</name></connection>
<intersection>-436.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,-436.5,337.5,-436.5</points>
<intersection>323.5 2</intersection>
<intersection>337.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323.5,-436.5,323.5,-423.5</points>
<intersection>-436.5 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323.5,-432,327.5,-432</points>
<connection>
<GID>3568</GID>
<name>IN_0</name></connection>
<intersection>323.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321.5,-423.5,323.5,-423.5</points>
<connection>
<GID>3570</GID>
<name>OUT_0</name></connection>
<intersection>323.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,334.5,276.5,354</points>
<connection>
<GID>4822</GID>
<name>N_in1</name></connection>
<intersection>354 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>278,354,278,374</points>
<connection>
<GID>5534</GID>
<name>N_in0</name></connection>
<intersection>354 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>276.5,354,278,354</points>
<intersection>276.5 0</intersection>
<intersection>278 1</intersection></hsegment></shape></wire>
<wire>
<ID>2556</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>365,-433,367,-433</points>
<connection>
<GID>3571</GID>
<name>OUT</name></connection>
<connection>
<GID>3572</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,-436,369,-436</points>
<connection>
<GID>3572</GID>
<name>IN_0</name></connection>
<intersection>355 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>355,-436,355,-423.5</points>
<intersection>-436 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>355,-432,359,-432</points>
<connection>
<GID>3571</GID>
<name>IN_0</name></connection>
<intersection>355 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352.5,-423.5,355,-423.5</points>
<connection>
<GID>3573</GID>
<name>OUT_0</name></connection>
<intersection>355 2</intersection></hsegment></shape></wire>
<wire>
<ID>4101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,341.5,305.5,366.5</points>
<connection>
<GID>4936</GID>
<name>N_in1</name></connection>
<connection>
<GID>5771</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>2558</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394.5,-433,396.5,-433</points>
<connection>
<GID>3574</GID>
<name>OUT</name></connection>
<connection>
<GID>3575</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,334.5,308.5,354</points>
<connection>
<GID>4823</GID>
<name>N_in1</name></connection>
<intersection>354 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>310,354,310,374</points>
<connection>
<GID>5535</GID>
<name>N_in0</name></connection>
<intersection>354 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308.5,354,310,354</points>
<intersection>308.5 0</intersection>
<intersection>310 1</intersection></hsegment></shape></wire>
<wire>
<ID>2559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398.5,-436.5,398.5,-436</points>
<connection>
<GID>3575</GID>
<name>IN_0</name></connection>
<intersection>-436.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-436.5,398.5,-436.5</points>
<intersection>384.5 2</intersection>
<intersection>398.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384.5,-436.5,384.5,-423.5</points>
<intersection>-436.5 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384.5,-432,388.5,-432</points>
<connection>
<GID>3574</GID>
<name>IN_0</name></connection>
<intersection>384.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382.5,-423.5,384.5,-423.5</points>
<connection>
<GID>3576</GID>
<name>OUT_0</name></connection>
<intersection>384.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,341.5,337.5,354</points>
<connection>
<GID>4935</GID>
<name>N_in1</name></connection>
<intersection>354 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>339,354,339,367</points>
<connection>
<GID>5644</GID>
<name>N_in0</name></connection>
<intersection>354 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,354,339,354</points>
<intersection>337.5 0</intersection>
<intersection>339 1</intersection></hsegment></shape></wire>
<wire>
<ID>2560</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>426,-433,428,-433</points>
<connection>
<GID>3577</GID>
<name>OUT</name></connection>
<connection>
<GID>3578</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,334.5,339.5,354.5</points>
<connection>
<GID>4917</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>341,354.5,341,375</points>
<connection>
<GID>5536</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>339.5,354.5,341,354.5</points>
<intersection>339.5 0</intersection>
<intersection>341 1</intersection></hsegment></shape></wire>
<wire>
<ID>2561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>416,-436,430,-436</points>
<connection>
<GID>3578</GID>
<name>IN_0</name></connection>
<intersection>416 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>416,-436,416,-423.5</points>
<intersection>-436 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>416,-432,420,-432</points>
<connection>
<GID>3577</GID>
<name>IN_0</name></connection>
<intersection>416 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413.5,-423.5,416,-423.5</points>
<connection>
<GID>3579</GID>
<name>OUT_0</name></connection>
<intersection>416 2</intersection></hsegment></shape></wire>
<wire>
<ID>4105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,341.5,368,354.5</points>
<connection>
<GID>4934</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>369.5,354.5,369.5,367.5</points>
<connection>
<GID>5645</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368,354.5,369.5,354.5</points>
<intersection>368 0</intersection>
<intersection>369.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2562</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456.5,-433,458.5,-433</points>
<connection>
<GID>3580</GID>
<name>OUT</name></connection>
<connection>
<GID>3581</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370.5,334,370.5,355</points>
<connection>
<GID>4918</GID>
<name>N_in1</name></connection>
<intersection>355 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>371,355,371,376</points>
<connection>
<GID>5537</GID>
<name>N_in0</name></connection>
<intersection>355 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>370.5,355,371,355</points>
<intersection>370.5 0</intersection>
<intersection>371 1</intersection></hsegment></shape></wire>
<wire>
<ID>2563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460.5,-436.5,460.5,-436</points>
<connection>
<GID>3581</GID>
<name>IN_0</name></connection>
<intersection>-436.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446.5,-436.5,460.5,-436.5</points>
<intersection>446.5 2</intersection>
<intersection>460.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446.5,-436.5,446.5,-423.5</points>
<intersection>-436.5 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446.5,-432,450.5,-432</points>
<connection>
<GID>3580</GID>
<name>IN_0</name></connection>
<intersection>446.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444.5,-423.5,446.5,-423.5</points>
<connection>
<GID>3582</GID>
<name>OUT_0</name></connection>
<intersection>446.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398.5,341.5,398.5,354.5</points>
<connection>
<GID>4933</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>400,354.5,400,367.5</points>
<connection>
<GID>5646</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>398.5,354.5,400,354.5</points>
<intersection>398.5 0</intersection>
<intersection>400 1</intersection></hsegment></shape></wire>
<wire>
<ID>2564</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>488,-433,490,-433</points>
<connection>
<GID>3583</GID>
<name>OUT</name></connection>
<connection>
<GID>3584</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,334.5,400.5,355.5</points>
<connection>
<GID>4919</GID>
<name>N_in1</name></connection>
<intersection>355.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>402,355.5,402,376.5</points>
<connection>
<GID>5538</GID>
<name>N_in0</name></connection>
<intersection>355.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>400.5,355.5,402,355.5</points>
<intersection>400.5 0</intersection>
<intersection>402 1</intersection></hsegment></shape></wire>
<wire>
<ID>2565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>478,-436,492,-436</points>
<connection>
<GID>3584</GID>
<name>IN_0</name></connection>
<intersection>478 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>478,-436,478,-423.5</points>
<intersection>-436 1</intersection>
<intersection>-432 4</intersection>
<intersection>-423.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>478,-432,482,-432</points>
<connection>
<GID>3583</GID>
<name>IN_0</name></connection>
<intersection>478 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475.5,-423.5,478,-423.5</points>
<connection>
<GID>3585</GID>
<name>OUT_0</name></connection>
<intersection>478 2</intersection></hsegment></shape></wire>
<wire>
<ID>4109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,341.5,429.5,354.5</points>
<connection>
<GID>4932</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>431,354.5,431,367.5</points>
<connection>
<GID>5647</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>429.5,354.5,431,354.5</points>
<intersection>429.5 0</intersection>
<intersection>431 1</intersection></hsegment></shape></wire>
<wire>
<ID>2566</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>272,-417.5,274,-417.5</points>
<connection>
<GID>3586</GID>
<name>OUT</name></connection>
<connection>
<GID>3587</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,334.5,431.5,356</points>
<connection>
<GID>4920</GID>
<name>N_in1</name></connection>
<intersection>356 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>433,356,433,377.5</points>
<connection>
<GID>5540</GID>
<name>N_in0</name></connection>
<intersection>356 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>431.5,356,433,356</points>
<intersection>431.5 0</intersection>
<intersection>433 1</intersection></hsegment></shape></wire>
<wire>
<ID>2567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-421,276,-420.5</points>
<connection>
<GID>3587</GID>
<name>IN_0</name></connection>
<intersection>-421 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-421,276,-421</points>
<intersection>262 2</intersection>
<intersection>276 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>262,-421,262,-408</points>
<intersection>-421 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>262,-416.5,266,-416.5</points>
<connection>
<GID>3586</GID>
<name>IN_0</name></connection>
<intersection>262 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>260,-408,262,-408</points>
<connection>
<GID>3588</GID>
<name>OUT_0</name></connection>
<intersection>262 2</intersection></hsegment></shape></wire>
<wire>
<ID>4111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460.5,342.5,460.5,354.5</points>
<connection>
<GID>4931</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>462,354.5,462,367</points>
<connection>
<GID>5648</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>460.5,354.5,462,354.5</points>
<intersection>460.5 0</intersection>
<intersection>462 1</intersection></hsegment></shape></wire>
<wire>
<ID>2568</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>303.5,-417.5,305.5,-417.5</points>
<connection>
<GID>3589</GID>
<name>OUT</name></connection>
<connection>
<GID>3590</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,334,462.5,354.5</points>
<connection>
<GID>4921</GID>
<name>N_in1</name></connection>
<intersection>354.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>464,354.5,464,375.5</points>
<connection>
<GID>5539</GID>
<name>N_in0</name></connection>
<intersection>354.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462.5,354.5,464,354.5</points>
<intersection>462.5 0</intersection>
<intersection>464 1</intersection></hsegment></shape></wire>
<wire>
<ID>2569</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293.5,-420.5,307.5,-420.5</points>
<connection>
<GID>3590</GID>
<name>IN_0</name></connection>
<intersection>293.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>293.5,-420.5,293.5,-408</points>
<intersection>-420.5 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>293.5,-416.5,297.5,-416.5</points>
<connection>
<GID>3589</GID>
<name>IN_0</name></connection>
<intersection>293.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>291,-408,293.5,-408</points>
<connection>
<GID>3591</GID>
<name>OUT_0</name></connection>
<intersection>293.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,343,491,355</points>
<connection>
<GID>4930</GID>
<name>N_in1</name></connection>
<intersection>355 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>492.5,355,492.5,367.5</points>
<connection>
<GID>5649</GID>
<name>N_in0</name></connection>
<intersection>355 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>491,355,492.5,355</points>
<intersection>491 0</intersection>
<intersection>492.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2570</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>334,-417.5,336,-417.5</points>
<connection>
<GID>3592</GID>
<name>OUT</name></connection>
<connection>
<GID>3593</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,173,491,184</points>
<connection>
<GID>4929</GID>
<name>N_in0</name></connection>
<intersection>173 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>496,162,496,173</points>
<connection>
<GID>4210</GID>
<name>N_in1</name></connection>
<intersection>173 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>491,173,496,173</points>
<intersection>491 0</intersection>
<intersection>496 1</intersection></hsegment></shape></wire>
<wire>
<ID>2571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338,-421,338,-420.5</points>
<connection>
<GID>3593</GID>
<name>IN_0</name></connection>
<intersection>-421 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324,-421,338,-421</points>
<intersection>324 2</intersection>
<intersection>338 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>324,-421,324,-408</points>
<intersection>-421 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>324,-416.5,328,-416.5</points>
<connection>
<GID>3592</GID>
<name>IN_0</name></connection>
<intersection>324 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>322,-408,324,-408</points>
<connection>
<GID>3594</GID>
<name>OUT_0</name></connection>
<intersection>324 2</intersection></hsegment></shape></wire>
<wire>
<ID>4115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,174.5,462.5,192</points>
<connection>
<GID>4819</GID>
<name>N_in0</name></connection>
<intersection>174.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>467.5,153,467.5,174.5</points>
<connection>
<GID>4201</GID>
<name>N_in1</name></connection>
<intersection>174.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462.5,174.5,467.5,174.5</points>
<intersection>462.5 0</intersection>
<intersection>467.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2572</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>365.5,-417.5,367.5,-417.5</points>
<connection>
<GID>3595</GID>
<name>OUT</name></connection>
<connection>
<GID>3596</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460.5,172.5,460.5,183.5</points>
<connection>
<GID>4928</GID>
<name>N_in0</name></connection>
<intersection>172.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>465.5,161.5,465.5,172.5</points>
<connection>
<GID>4211</GID>
<name>N_in1</name></connection>
<intersection>172.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>460.5,172.5,465.5,172.5</points>
<intersection>460.5 0</intersection>
<intersection>465.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355.5,-420.5,369.5,-420.5</points>
<connection>
<GID>3596</GID>
<name>IN_0</name></connection>
<intersection>355.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>355.5,-420.5,355.5,-408</points>
<intersection>-420.5 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>355.5,-416.5,359.5,-416.5</points>
<connection>
<GID>3595</GID>
<name>IN_0</name></connection>
<intersection>355.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>353,-408,355.5,-408</points>
<connection>
<GID>3597</GID>
<name>OUT_0</name></connection>
<intersection>355.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,153.5,436.5,173.5</points>
<connection>
<GID>4200</GID>
<name>N_in1</name></connection>
<intersection>173.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>431.5,173.5,431.5,194</points>
<connection>
<GID>4820</GID>
<name>N_in0</name></connection>
<intersection>173.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>431.5,173.5,436.5,173.5</points>
<intersection>431.5 1</intersection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2574</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>395,-417.5,397,-417.5</points>
<connection>
<GID>3598</GID>
<name>OUT</name></connection>
<connection>
<GID>3599</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,172,429.5,184</points>
<connection>
<GID>4927</GID>
<name>N_in0</name></connection>
<intersection>172 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>434.5,160.5,434.5,172</points>
<connection>
<GID>4212</GID>
<name>N_in1</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>429.5,172,434.5,172</points>
<intersection>429.5 0</intersection>
<intersection>434.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,-421,399,-420.5</points>
<connection>
<GID>3599</GID>
<name>IN_0</name></connection>
<intersection>-421 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>385,-421,399,-421</points>
<intersection>385 2</intersection>
<intersection>399 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>385,-421,385,-408</points>
<intersection>-421 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>385,-416.5,389,-416.5</points>
<connection>
<GID>3598</GID>
<name>IN_0</name></connection>
<intersection>385 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>383,-408,385,-408</points>
<connection>
<GID>3600</GID>
<name>OUT_0</name></connection>
<intersection>385 2</intersection></hsegment></shape></wire>
<wire>
<ID>4119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,160.5,403.5,172</points>
<connection>
<GID>4213</GID>
<name>N_in1</name></connection>
<intersection>172 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>398.5,172,398.5,184</points>
<connection>
<GID>4926</GID>
<name>N_in0</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>398.5,172,403.5,172</points>
<intersection>398.5 1</intersection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2576</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>426.5,-417.5,428.5,-417.5</points>
<connection>
<GID>3601</GID>
<name>OUT</name></connection>
<connection>
<GID>3602</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405.5,153.5,405.5,173</points>
<connection>
<GID>4199</GID>
<name>N_in1</name></connection>
<intersection>173 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>400.5,173,400.5,193</points>
<connection>
<GID>4818</GID>
<name>N_in0</name></connection>
<intersection>173 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>400.5,173,405.5,173</points>
<intersection>400.5 1</intersection>
<intersection>405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>416.5,-420.5,430.5,-420.5</points>
<connection>
<GID>3602</GID>
<name>IN_0</name></connection>
<intersection>416.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>416.5,-420.5,416.5,-408</points>
<intersection>-420.5 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>416.5,-416.5,420.5,-416.5</points>
<connection>
<GID>3601</GID>
<name>IN_0</name></connection>
<intersection>416.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>414,-408,416.5,-408</points>
<connection>
<GID>3603</GID>
<name>OUT_0</name></connection>
<intersection>416.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,160.5,373,172</points>
<connection>
<GID>4214</GID>
<name>N_in1</name></connection>
<intersection>172 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>368,172,368,184</points>
<connection>
<GID>4925</GID>
<name>N_in0</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368,172,373,172</points>
<intersection>368 1</intersection>
<intersection>373 0</intersection></hsegment></shape></wire>
<wire>
<ID>2578</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>457,-417.5,459,-417.5</points>
<connection>
<GID>3604</GID>
<name>OUT</name></connection>
<connection>
<GID>3605</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,153,375.5,172.5</points>
<connection>
<GID>4198</GID>
<name>N_in1</name></connection>
<intersection>172.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>369.5,172.5,369.5,192.5</points>
<connection>
<GID>4817</GID>
<name>N_in0</name></connection>
<intersection>172.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>369.5,172.5,375.5,172.5</points>
<intersection>369.5 1</intersection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461,-421,461,-420.5</points>
<connection>
<GID>3605</GID>
<name>IN_0</name></connection>
<intersection>-421 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>447,-421,461,-421</points>
<intersection>447 2</intersection>
<intersection>461 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>447,-421,447,-408</points>
<intersection>-421 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>447,-416.5,451,-416.5</points>
<connection>
<GID>3604</GID>
<name>IN_0</name></connection>
<intersection>447 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>445,-408,447,-408</points>
<connection>
<GID>3606</GID>
<name>OUT_0</name></connection>
<intersection>447 2</intersection></hsegment></shape></wire>
<wire>
<ID>4123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342.5,160.5,342.5,172</points>
<connection>
<GID>4215</GID>
<name>N_in1</name></connection>
<intersection>172 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>337.5,172,337.5,183.5</points>
<connection>
<GID>4924</GID>
<name>N_in0</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>337.5,172,342.5,172</points>
<intersection>337.5 1</intersection>
<intersection>342.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2580</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>488.5,-417.5,490.5,-417.5</points>
<connection>
<GID>3607</GID>
<name>OUT</name></connection>
<connection>
<GID>3608</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,153.5,344.5,172.5</points>
<connection>
<GID>4197</GID>
<name>N_in1</name></connection>
<intersection>172.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>339.5,172.5,339.5,191.5</points>
<connection>
<GID>4816</GID>
<name>N_in0</name></connection>
<intersection>172.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>339.5,172.5,344.5,172.5</points>
<intersection>339.5 1</intersection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>478.5,-420.5,492.5,-420.5</points>
<connection>
<GID>3608</GID>
<name>IN_0</name></connection>
<intersection>478.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>478.5,-420.5,478.5,-408</points>
<intersection>-420.5 1</intersection>
<intersection>-416.5 4</intersection>
<intersection>-408 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>478.5,-416.5,482.5,-416.5</points>
<connection>
<GID>3607</GID>
<name>IN_0</name></connection>
<intersection>478.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>476,-408,478.5,-408</points>
<connection>
<GID>3609</GID>
<name>OUT_0</name></connection>
<intersection>478.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>4125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,153.5,313.5,177</points>
<connection>
<GID>4103</GID>
<name>N_in1</name></connection>
<intersection>177 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>308.5,177,308.5,190.5</points>
<connection>
<GID>4815</GID>
<name>N_in0</name></connection>
<intersection>177 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308.5,177,313.5,177</points>
<intersection>308.5 1</intersection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2582</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-541,250.5,-401.5</points>
<connection>
<GID>3373</GID>
<name>N_in1</name></connection>
<connection>
<GID>3381</GID>
<name>N_in0</name></connection>
<intersection>-521.5 14</intersection>
<intersection>-504.5 12</intersection>
<intersection>-488.5 10</intersection>
<intersection>-473 8</intersection>
<intersection>-456.5 6</intersection>
<intersection>-439.5 4</intersection>
<intersection>-423.5 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-408,254,-408</points>
<connection>
<GID>3588</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>250.5,-423.5,253.5,-423.5</points>
<connection>
<GID>3564</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>250.5,-439.5,253,-439.5</points>
<connection>
<GID>3540</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>250.5,-456.5,252.5,-456.5</points>
<connection>
<GID>3508</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>250.5,-473,253,-473</points>
<connection>
<GID>3455</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>250.5,-488.5,252.5,-488.5</points>
<connection>
<GID>3431</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>250.5,-504.5,252,-504.5</points>
<connection>
<GID>3407</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>250.5,-521.5,251.5,-521.5</points>
<connection>
<GID>3372</GID>
<name>IN_0</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,160.5,279.5,171.5</points>
<connection>
<GID>4202</GID>
<name>N_in1</name></connection>
<intersection>171.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>274.5,171.5,274.5,182.5</points>
<connection>
<GID>4923</GID>
<name>N_in0</name></connection>
<intersection>171.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>274.5,171.5,279.5,171.5</points>
<intersection>274.5 1</intersection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,-418.5,482.5,-418.5</points>
<connection>
<GID>3586</GID>
<name>IN_1</name></connection>
<connection>
<GID>3589</GID>
<name>IN_1</name></connection>
<connection>
<GID>3592</GID>
<name>IN_1</name></connection>
<connection>
<GID>3595</GID>
<name>IN_1</name></connection>
<connection>
<GID>3598</GID>
<name>IN_1</name></connection>
<connection>
<GID>3601</GID>
<name>IN_1</name></connection>
<connection>
<GID>3604</GID>
<name>IN_1</name></connection>
<connection>
<GID>3607</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,-418.5,246,-415.5</points>
<connection>
<GID>3509</GID>
<name>OUT_0</name></connection>
<intersection>-418.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,153.5,281.5,172</points>
<connection>
<GID>4102</GID>
<name>N_in1</name></connection>
<intersection>172 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>276.5,172,276.5,190.5</points>
<connection>
<GID>4814</GID>
<name>N_in0</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>276.5,172,281.5,172</points>
<intersection>276.5 1</intersection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>240,-411,470,-411</points>
<connection>
<GID>3510</GID>
<name>OUT</name></connection>
<connection>
<GID>3588</GID>
<name>clock</name></connection>
<connection>
<GID>3591</GID>
<name>clock</name></connection>
<connection>
<GID>3594</GID>
<name>clock</name></connection>
<connection>
<GID>3597</GID>
<name>clock</name></connection>
<connection>
<GID>3600</GID>
<name>clock</name></connection>
<connection>
<GID>3603</GID>
<name>clock</name></connection>
<connection>
<GID>3606</GID>
<name>clock</name></connection>
<connection>
<GID>3609</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>4128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,153.5,250.5,172</points>
<connection>
<GID>4101</GID>
<name>N_in1</name></connection>
<intersection>172 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>245.5,172,245.5,191</points>
<connection>
<GID>4813</GID>
<name>N_in0</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>245.5,172,250.5,172</points>
<intersection>245.5 1</intersection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,160.5,310.5,175.5</points>
<connection>
<GID>4216</GID>
<name>N_in1</name></connection>
<intersection>175.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>303.5,175.5,303.5,190.5</points>
<connection>
<GID>5773</GID>
<name>N_in0</name></connection>
<intersection>175.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>303.5,175.5,310.5,175.5</points>
<intersection>303.5 1</intersection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-50.5,249.5,-20</points>
<connection>
<GID>2181</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>250.5,-20,250.5,10</points>
<connection>
<GID>4093</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-20,250.5,-20</points>
<intersection>249.5 0</intersection>
<intersection>250.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-43.5,278.5,-21</points>
<connection>
<GID>2282</GID>
<name>N_in1</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>279.5,-21,279.5,1.5</points>
<connection>
<GID>4203</GID>
<name>N_in0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>278.5,-21,279.5,-21</points>
<intersection>278.5 0</intersection>
<intersection>279.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-50.5,280.5,-20.5</points>
<connection>
<GID>2182</GID>
<name>N_in1</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>281.5,-20.5,281.5,9.5</points>
<connection>
<GID>4094</GID>
<name>N_in0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>280.5,-20.5,281.5,-20.5</points>
<intersection>280.5 0</intersection>
<intersection>281.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-43.5,309.5,-20</points>
<connection>
<GID>2296</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>309,-20,309,3</points>
<connection>
<GID>5775</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>309,-20,309.5,-20</points>
<intersection>309 1</intersection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-50.5,312.5,-20.5</points>
<connection>
<GID>2183</GID>
<name>N_in1</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>313.5,-20.5,313.5,9.5</points>
<connection>
<GID>4095</GID>
<name>N_in0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>312.5,-20.5,313.5,-20.5</points>
<intersection>312.5 0</intersection>
<intersection>313.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-43.5,341.5,-20.5</points>
<connection>
<GID>2295</GID>
<name>N_in1</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>342.5,-20.5,342.5,2.5</points>
<connection>
<GID>4204</GID>
<name>N_in0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-20.5,342.5,-20.5</points>
<intersection>341.5 0</intersection>
<intersection>342.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343.5,-50.5,343.5,-20</points>
<connection>
<GID>2277</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>344.5,-20,344.5,10.5</points>
<connection>
<GID>4096</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>343.5,-20,344.5,-20</points>
<intersection>343.5 0</intersection>
<intersection>344.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-43.5,372,-20</points>
<connection>
<GID>2294</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>373,-20,373,3</points>
<connection>
<GID>4205</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>372,-20,373,-20</points>
<intersection>372 0</intersection>
<intersection>373 1</intersection></hsegment></shape></wire>
<wire>
<ID>4138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374.5,-51,374.5,11.5</points>
<connection>
<GID>2278</GID>
<name>N_in1</name></connection>
<connection>
<GID>4097</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-43.5,402.5,-20</points>
<connection>
<GID>2293</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>403.5,-20,403.5,3</points>
<connection>
<GID>4206</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>402.5,-20,403.5,-20</points>
<intersection>402.5 0</intersection>
<intersection>403.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404.5,-50.5,404.5,-19</points>
<connection>
<GID>2279</GID>
<name>N_in1</name></connection>
<intersection>-19 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>405.5,-19,405.5,12</points>
<connection>
<GID>4098</GID>
<name>N_in0</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>404.5,-19,405.5,-19</points>
<intersection>404.5 0</intersection>
<intersection>405.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,-43.5,433.5,-20</points>
<connection>
<GID>2292</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>434.5,-20,434.5,3</points>
<connection>
<GID>4207</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-20,434.5,-20</points>
<intersection>433.5 0</intersection>
<intersection>434.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,-50.5,435.5,-18.5</points>
<connection>
<GID>2280</GID>
<name>N_in1</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>436.5,-18.5,436.5,13</points>
<connection>
<GID>4100</GID>
<name>N_in0</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>435.5,-18.5,436.5,-18.5</points>
<intersection>435.5 0</intersection>
<intersection>436.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,-42.5,464.5,-20</points>
<connection>
<GID>2291</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>465.5,-20,465.5,2.5</points>
<connection>
<GID>4208</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>464.5,-20,465.5,-20</points>
<intersection>464.5 0</intersection>
<intersection>465.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466.5,-51,466.5,-20</points>
<connection>
<GID>2281</GID>
<name>N_in1</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>467.5,-20,467.5,11</points>
<connection>
<GID>4099</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>466.5,-20,467.5,-20</points>
<intersection>466.5 0</intersection>
<intersection>467.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495,-42,495,-19.5</points>
<connection>
<GID>2290</GID>
<name>N_in1</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>496,-19.5,496,3</points>
<connection>
<GID>4209</GID>
<name>N_in0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>495,-19.5,496,-19.5</points>
<intersection>495 0</intersection>
<intersection>496 1</intersection></hsegment></shape></wire>
<wire>
<ID>4146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495,-209.5,495,-201</points>
<connection>
<GID>2289</GID>
<name>N_in0</name></connection>
<intersection>-209.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>493,-218,493,-209.5</points>
<connection>
<GID>3250</GID>
<name>N_in1</name></connection>
<intersection>-209.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>493,-209.5,495,-209.5</points>
<intersection>493 1</intersection>
<intersection>495 0</intersection></hsegment></shape></wire>
<wire>
<ID>4147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466.5,-227,466.5,-193</points>
<connection>
<GID>2179</GID>
<name>N_in0</name></connection>
<intersection>-227 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>464.5,-227,466.5,-227</points>
<connection>
<GID>3241</GID>
<name>N_in1</name></connection>
<intersection>466.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>464.5,-210,464.5,-201.5</points>
<connection>
<GID>2288</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>462.5,-218.5,462.5,-210</points>
<connection>
<GID>3251</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462.5,-210,464.5,-210</points>
<intersection>462.5 1</intersection>
<intersection>464.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-226.5,434.5,-208.5</points>
<intersection>-226.5 3</intersection>
<intersection>-208.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>435.5,-208.5,435.5,-191</points>
<connection>
<GID>2180</GID>
<name>N_in0</name></connection>
<intersection>-208.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434.5,-208.5,435.5,-208.5</points>
<intersection>434.5 0</intersection>
<intersection>435.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>433.5,-226.5,434.5,-226.5</points>
<connection>
<GID>3240</GID>
<name>N_in1</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,-219.5,431.5,-210</points>
<connection>
<GID>3252</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>433.5,-210,433.5,-201</points>
<connection>
<GID>2287</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-210,433.5,-210</points>
<intersection>431.5 0</intersection>
<intersection>433.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,-226.5,403.5,-209</points>
<intersection>-226.5 3</intersection>
<intersection>-209 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>404.5,-209,404.5,-192</points>
<connection>
<GID>2178</GID>
<name>N_in0</name></connection>
<intersection>-209 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>403.5,-209,404.5,-209</points>
<intersection>403.5 0</intersection>
<intersection>404.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>402.5,-226.5,403.5,-226.5</points>
<connection>
<GID>3239</GID>
<name>N_in1</name></connection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,-219.5,400.5,-210</points>
<connection>
<GID>3253</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>402.5,-210,402.5,-201</points>
<connection>
<GID>2286</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>400.5,-210,402.5,-210</points>
<intersection>400.5 0</intersection>
<intersection>402.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,-219.5,370,-210</points>
<connection>
<GID>3254</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>372,-210,372,-201</points>
<connection>
<GID>2285</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>370,-210,372,-210</points>
<intersection>370 0</intersection>
<intersection>372 1</intersection></hsegment></shape></wire>
<wire>
<ID>4154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372.5,-227,372.5,-209.5</points>
<connection>
<GID>3238</GID>
<name>N_in1</name></connection>
<intersection>-209.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>373.5,-209.5,373.5,-192.5</points>
<connection>
<GID>2177</GID>
<name>N_in0</name></connection>
<intersection>-209.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-209.5,373.5,-209.5</points>
<intersection>372.5 0</intersection>
<intersection>373.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,-219.5,339.5,-210.5</points>
<connection>
<GID>3255</GID>
<name>N_in1</name></connection>
<intersection>-210.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>341.5,-210.5,341.5,-201.5</points>
<connection>
<GID>2284</GID>
<name>N_in0</name></connection>
<intersection>-210.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-210.5,341.5,-210.5</points>
<intersection>339.5 0</intersection>
<intersection>341.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-226.5,341.5,-210</points>
<connection>
<GID>3237</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>343.5,-210,343.5,-193.5</points>
<connection>
<GID>2176</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-210,343.5,-210</points>
<intersection>341.5 0</intersection>
<intersection>343.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-219.5,307.5,-210</points>
<connection>
<GID>3256</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>306,-210,306,-200.5</points>
<connection>
<GID>5777</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>306,-210,307.5,-210</points>
<intersection>306 1</intersection>
<intersection>307.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-226.5,310.5,-210.5</points>
<connection>
<GID>3143</GID>
<name>N_in1</name></connection>
<intersection>-210.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>312.5,-210.5,312.5,-194.5</points>
<connection>
<GID>2175</GID>
<name>N_in0</name></connection>
<intersection>-210.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>310.5,-210.5,312.5,-210.5</points>
<intersection>310.5 0</intersection>
<intersection>312.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,-219.5,276.5,-211</points>
<connection>
<GID>3242</GID>
<name>N_in1</name></connection>
<intersection>-211 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>278.5,-211,278.5,-202.5</points>
<connection>
<GID>2283</GID>
<name>N_in0</name></connection>
<intersection>-211 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>276.5,-211,278.5,-211</points>
<intersection>276.5 0</intersection>
<intersection>278.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-226.5,279.5,-210.5</points>
<intersection>-226.5 3</intersection>
<intersection>-210.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>280.5,-210.5,280.5,-194.5</points>
<connection>
<GID>2174</GID>
<name>N_in0</name></connection>
<intersection>-210.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>279.5,-210.5,280.5,-210.5</points>
<intersection>279.5 0</intersection>
<intersection>280.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>278.5,-226.5,279.5,-226.5</points>
<connection>
<GID>3142</GID>
<name>N_in1</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-226.5,247.5,-210</points>
<connection>
<GID>3141</GID>
<name>N_in1</name></connection>
<intersection>-210 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>249.5,-210,249.5,-194</points>
<connection>
<GID>2173</GID>
<name>N_in0</name></connection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-210,249.5,-210</points>
<intersection>247.5 0</intersection>
<intersection>249.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-399.5,250.5,-384.5</points>
<connection>
<GID>3381</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>247.5,-384.5,247.5,-370</points>
<connection>
<GID>3133</GID>
<name>N_in0</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-384.5,250.5,-384.5</points>
<intersection>247.5 1</intersection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-392.5,279.5,-385.5</points>
<connection>
<GID>3482</GID>
<name>N_in1</name></connection>
<intersection>-385.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>276.5,-385.5,276.5,-378.5</points>
<connection>
<GID>3243</GID>
<name>N_in0</name></connection>
<intersection>-385.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>276.5,-385.5,279.5,-385.5</points>
<intersection>276.5 1</intersection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-399.5,281.5,-385</points>
<connection>
<GID>3382</GID>
<name>N_in1</name></connection>
<intersection>-385 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>278.5,-385,278.5,-370.5</points>
<connection>
<GID>3134</GID>
<name>N_in0</name></connection>
<intersection>-385 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>278.5,-385,281.5,-385</points>
<intersection>278.5 1</intersection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-392.5,310.5,-383.5</points>
<connection>
<GID>3496</GID>
<name>N_in1</name></connection>
<intersection>-383.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>303.5,-383.5,303.5,-375</points>
<connection>
<GID>5779</GID>
<name>N_in0</name></connection>
<intersection>-383.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-383.5,310.5,-383.5</points>
<intersection>303.5 1</intersection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-399.5,313.5,-385</points>
<connection>
<GID>3383</GID>
<name>N_in1</name></connection>
<intersection>-385 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>313,-385,313,-370.5</points>
<intersection>-385 2</intersection>
<intersection>-370.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>313,-385,313.5,-385</points>
<intersection>313 1</intersection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>310.5,-370.5,313,-370.5</points>
<connection>
<GID>3135</GID>
<name>N_in0</name></connection>
<intersection>313 1</intersection></hsegment></shape></wire>
<wire>
<ID>4167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342.5,-392.5,342.5,-385</points>
<connection>
<GID>3495</GID>
<name>N_in1</name></connection>
<intersection>-385 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>339.5,-385,339.5,-377.5</points>
<connection>
<GID>3244</GID>
<name>N_in0</name></connection>
<intersection>-385 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-385,342.5,-385</points>
<intersection>339.5 1</intersection>
<intersection>342.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,-399.5,344.5,-384.5</points>
<connection>
<GID>3477</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>341.5,-384.5,341.5,-369.5</points>
<connection>
<GID>3136</GID>
<name>N_in0</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-384.5,344.5,-384.5</points>
<intersection>341.5 1</intersection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,-392.5,373,-384.5</points>
<connection>
<GID>3494</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>370,-384.5,370,-377</points>
<connection>
<GID>3245</GID>
<name>N_in0</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>370,-384.5,373,-384.5</points>
<intersection>370 1</intersection>
<intersection>373 0</intersection></hsegment></shape></wire>
<wire>
<ID>4170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-400,375.5,-384</points>
<connection>
<GID>3478</GID>
<name>N_in1</name></connection>
<intersection>-384 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>371.5,-384,371.5,-368.5</points>
<connection>
<GID>3137</GID>
<name>N_in0</name></connection>
<intersection>-384 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>371.5,-384,375.5,-384</points>
<intersection>371.5 1</intersection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,-392.5,403.5,-384.5</points>
<connection>
<GID>3493</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>400.5,-384.5,400.5,-377</points>
<connection>
<GID>3246</GID>
<name>N_in0</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>400.5,-384.5,403.5,-384.5</points>
<intersection>400.5 1</intersection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405.5,-399.5,405.5,-383.5</points>
<connection>
<GID>3479</GID>
<name>N_in1</name></connection>
<intersection>-383.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>402.5,-383.5,402.5,-368</points>
<connection>
<GID>3138</GID>
<name>N_in0</name></connection>
<intersection>-383.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>402.5,-383.5,405.5,-383.5</points>
<intersection>402.5 1</intersection>
<intersection>405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-392.5,434.5,-384.5</points>
<connection>
<GID>3492</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>431.5,-384.5,431.5,-377</points>
<connection>
<GID>3247</GID>
<name>N_in0</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-384.5,434.5,-384.5</points>
<intersection>431.5 1</intersection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,-399.5,436.5,-383</points>
<connection>
<GID>3480</GID>
<name>N_in1</name></connection>
<intersection>-383 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>433.5,-383,433.5,-367</points>
<connection>
<GID>3140</GID>
<name>N_in0</name></connection>
<intersection>-383 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-383,436.5,-383</points>
<intersection>433.5 1</intersection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465.5,-391.5,465.5,-384.5</points>
<connection>
<GID>3491</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>462.5,-384.5,462.5,-377.5</points>
<connection>
<GID>3248</GID>
<name>N_in0</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462.5,-384.5,465.5,-384.5</points>
<intersection>462.5 1</intersection>
<intersection>465.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467.5,-400,467.5,-384.5</points>
<connection>
<GID>3481</GID>
<name>N_in1</name></connection>
<intersection>-384.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>466,-384.5,466,-369</points>
<intersection>-384.5 2</intersection>
<intersection>-369 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>466,-384.5,467.5,-384.5</points>
<intersection>466 1</intersection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>464.5,-369,466,-369</points>
<connection>
<GID>3139</GID>
<name>N_in0</name></connection>
<intersection>466 1</intersection></hsegment></shape></wire>
<wire>
<ID>4177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496,-391,496,-384</points>
<connection>
<GID>3490</GID>
<name>N_in1</name></connection>
<intersection>-384 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>493,-384,493,-377</points>
<connection>
<GID>3249</GID>
<name>N_in0</name></connection>
<intersection>-384 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>493,-384,496,-384</points>
<intersection>493 1</intersection>
<intersection>496 0</intersection></hsegment></shape></wire>
<wire>
<ID>4178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-585.5,246.5,-564</points>
<connection>
<GID>3861</GID>
<name>N_in1</name></connection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>250.5,-564,250.5,-543</points>
<connection>
<GID>3373</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>246.5,-564,250.5,-564</points>
<intersection>246.5 0</intersection>
<intersection>250.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-578.5,275.5,-565</points>
<connection>
<GID>3962</GID>
<name>N_in1</name></connection>
<intersection>-565 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>279.5,-565,279.5,-551.5</points>
<connection>
<GID>3483</GID>
<name>N_in0</name></connection>
<intersection>-565 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>275.5,-565,279.5,-565</points>
<intersection>275.5 0</intersection>
<intersection>279.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-585.5,277.5,-564.5</points>
<connection>
<GID>3862</GID>
<name>N_in1</name></connection>
<intersection>-564.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>281.5,-564.5,281.5,-543.5</points>
<connection>
<GID>3374</GID>
<name>N_in0</name></connection>
<intersection>-564.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>277.5,-564.5,281.5,-564.5</points>
<intersection>277.5 0</intersection>
<intersection>281.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306.5,-578.5,306.5,-566.5</points>
<connection>
<GID>3976</GID>
<name>N_in1</name></connection>
<intersection>-566.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>306,-566.5,306,-555</points>
<connection>
<GID>5783</GID>
<name>N_in0</name></connection>
<intersection>-566.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>306,-566.5,306.5,-566.5</points>
<intersection>306 1</intersection>
<intersection>306.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-585.5,309.5,-564.5</points>
<connection>
<GID>3863</GID>
<name>N_in1</name></connection>
<intersection>-564.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>313.5,-564.5,313.5,-543.5</points>
<connection>
<GID>3375</GID>
<name>N_in0</name></connection>
<intersection>-564.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-564.5,313.5,-564.5</points>
<intersection>309.5 0</intersection>
<intersection>313.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,-578.5,338.5,-564.5</points>
<connection>
<GID>3975</GID>
<name>N_in1</name></connection>
<intersection>-564.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>342.5,-564.5,342.5,-550.5</points>
<connection>
<GID>3484</GID>
<name>N_in0</name></connection>
<intersection>-564.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>338.5,-564.5,342.5,-564.5</points>
<intersection>338.5 0</intersection>
<intersection>342.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>340.5,-585.5,340.5,-564</points>
<connection>
<GID>3957</GID>
<name>N_in1</name></connection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>344.5,-564,344.5,-542.5</points>
<connection>
<GID>3376</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>340.5,-564,344.5,-564</points>
<intersection>340.5 0</intersection>
<intersection>344.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-578.5,369,-564</points>
<connection>
<GID>3974</GID>
<name>N_in1</name></connection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>373,-564,373,-550</points>
<connection>
<GID>3485</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>369,-564,373,-564</points>
<intersection>369 0</intersection>
<intersection>373 1</intersection></hsegment></shape></wire>
<wire>
<ID>4186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>371.5,-586,371.5,-563.5</points>
<connection>
<GID>3958</GID>
<name>N_in1</name></connection>
<intersection>-563.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>374.5,-563.5,374.5,-541.5</points>
<connection>
<GID>3377</GID>
<name>N_in0</name></connection>
<intersection>-563.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>371.5,-563.5,374.5,-563.5</points>
<intersection>371.5 0</intersection>
<intersection>374.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,-578.5,399.5,-564</points>
<connection>
<GID>3973</GID>
<name>N_in1</name></connection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>403.5,-564,403.5,-550</points>
<connection>
<GID>3486</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>399.5,-564,403.5,-564</points>
<intersection>399.5 0</intersection>
<intersection>403.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>401.5,-585.5,401.5,-563</points>
<connection>
<GID>3959</GID>
<name>N_in1</name></connection>
<intersection>-563 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>405.5,-563,405.5,-541</points>
<connection>
<GID>3378</GID>
<name>N_in0</name></connection>
<intersection>-563 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>401.5,-563,405.5,-563</points>
<intersection>401.5 0</intersection>
<intersection>405.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,-578.5,430.5,-564</points>
<connection>
<GID>3972</GID>
<name>N_in1</name></connection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>434.5,-564,434.5,-550</points>
<connection>
<GID>3487</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>430.5,-564,434.5,-564</points>
<intersection>430.5 0</intersection>
<intersection>434.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,-585.5,432.5,-562.5</points>
<connection>
<GID>3960</GID>
<name>N_in1</name></connection>
<intersection>-562.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>436.5,-562.5,436.5,-540</points>
<connection>
<GID>3380</GID>
<name>N_in0</name></connection>
<intersection>-562.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>432.5,-562.5,436.5,-562.5</points>
<intersection>432.5 0</intersection>
<intersection>436.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461.5,-577.5,461.5,-564</points>
<connection>
<GID>3971</GID>
<name>N_in1</name></connection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>465.5,-564,465.5,-550.5</points>
<connection>
<GID>3488</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>461.5,-564,465.5,-564</points>
<intersection>461.5 0</intersection>
<intersection>465.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466.5,-586,466.5,-564</points>
<intersection>-586 3</intersection>
<intersection>-564 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>467.5,-564,467.5,-542</points>
<connection>
<GID>3379</GID>
<name>N_in0</name></connection>
<intersection>-564 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>466.5,-564,467.5,-564</points>
<intersection>466.5 0</intersection>
<intersection>467.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>463.5,-586,466.5,-586</points>
<connection>
<GID>3961</GID>
<name>N_in1</name></connection>
<intersection>466.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492,-577,492,-563.5</points>
<connection>
<GID>3970</GID>
<name>N_in1</name></connection>
<intersection>-563.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>496,-563.5,496,-550</points>
<connection>
<GID>3489</GID>
<name>N_in0</name></connection>
<intersection>-563.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>492,-563.5,496,-563.5</points>
<intersection>492 0</intersection>
<intersection>496 1</intersection></hsegment></shape></wire>
<wire>
<ID>4194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>487,-751,487,-743.5</points>
<connection>
<GID>5410</GID>
<name>N_in1</name></connection>
<intersection>-743.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>492,-743.5,492,-736</points>
<connection>
<GID>3969</GID>
<name>N_in0</name></connection>
<intersection>-743.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>487,-743.5,492,-743.5</points>
<intersection>487 0</intersection>
<intersection>492 1</intersection></hsegment></shape></wire>
<wire>
<ID>4195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-751.5,456.5,-744</points>
<connection>
<GID>5411</GID>
<name>N_in1</name></connection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>461.5,-744,461.5,-736.5</points>
<connection>
<GID>3968</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>456.5,-744,461.5,-744</points>
<intersection>456.5 0</intersection>
<intersection>461.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,-760,463,-744</points>
<intersection>-760 3</intersection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>463.5,-744,463.5,-728</points>
<connection>
<GID>3859</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>463,-744,463.5,-744</points>
<intersection>463 0</intersection>
<intersection>463.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>458.5,-760,463,-760</points>
<connection>
<GID>5401</GID>
<name>N_in1</name></connection>
<intersection>463 0</intersection></hsegment></shape></wire>
<wire>
<ID>4197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-752.5,425.5,-744</points>
<connection>
<GID>5412</GID>
<name>N_in1</name></connection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>430.5,-744,430.5,-736</points>
<connection>
<GID>3967</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>425.5,-744,430.5,-744</points>
<intersection>425.5 0</intersection>
<intersection>430.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-759.5,427.5,-742.5</points>
<connection>
<GID>5400</GID>
<name>N_in1</name></connection>
<intersection>-742.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>432.5,-742.5,432.5,-726</points>
<connection>
<GID>3860</GID>
<name>N_in0</name></connection>
<intersection>-742.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>427.5,-742.5,432.5,-742.5</points>
<intersection>427.5 0</intersection>
<intersection>432.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,-752.5,394.5,-744</points>
<connection>
<GID>5413</GID>
<name>N_in1</name></connection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>399.5,-744,399.5,-736</points>
<connection>
<GID>3966</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>394.5,-744,399.5,-744</points>
<intersection>394.5 0</intersection>
<intersection>399.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,-759.5,396.5,-743</points>
<connection>
<GID>5399</GID>
<name>N_in1</name></connection>
<intersection>-743 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>401.5,-743,401.5,-727</points>
<connection>
<GID>3858</GID>
<name>N_in0</name></connection>
<intersection>-743 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>396.5,-743,401.5,-743</points>
<intersection>396.5 0</intersection>
<intersection>401.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364,-752.5,364,-744</points>
<connection>
<GID>5414</GID>
<name>N_in1</name></connection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>369,-744,369,-736</points>
<connection>
<GID>3965</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>364,-744,369,-744</points>
<intersection>364 0</intersection>
<intersection>369 1</intersection></hsegment></shape></wire>
<wire>
<ID>4202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-760,366.5,-743.5</points>
<connection>
<GID>5398</GID>
<name>N_in1</name></connection>
<intersection>-743.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>370.5,-743.5,370.5,-727.5</points>
<connection>
<GID>3857</GID>
<name>N_in0</name></connection>
<intersection>-743.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>366.5,-743.5,370.5,-743.5</points>
<intersection>366.5 0</intersection>
<intersection>370.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,-752.5,333.5,-744.5</points>
<connection>
<GID>5415</GID>
<name>N_in1</name></connection>
<intersection>-744.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>338.5,-744.5,338.5,-736.5</points>
<connection>
<GID>3964</GID>
<name>N_in0</name></connection>
<intersection>-744.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>333.5,-744.5,338.5,-744.5</points>
<intersection>333.5 0</intersection>
<intersection>338.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-759.5,335.5,-744</points>
<connection>
<GID>5397</GID>
<name>N_in1</name></connection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>340.5,-744,340.5,-728.5</points>
<connection>
<GID>3856</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>335.5,-744,340.5,-744</points>
<intersection>335.5 0</intersection>
<intersection>340.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,-759.5,304.5,-730.5</points>
<connection>
<GID>5303</GID>
<name>N_in1</name></connection>
<intersection>-730.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>309.5,-730.5,309.5,-729.5</points>
<connection>
<GID>3855</GID>
<name>N_in0</name></connection>
<intersection>-730.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-730.5,309.5,-730.5</points>
<intersection>304.5 0</intersection>
<intersection>309.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-752.5,301.5,-731</points>
<connection>
<GID>5416</GID>
<name>N_in1</name></connection>
<connection>
<GID>5785</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-752.5,270.5,-745</points>
<connection>
<GID>5402</GID>
<name>N_in1</name></connection>
<intersection>-745 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>275.5,-745,275.5,-737.5</points>
<connection>
<GID>3963</GID>
<name>N_in0</name></connection>
<intersection>-745 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-745,275.5,-745</points>
<intersection>270.5 0</intersection>
<intersection>275.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-759.5,272.5,-744.5</points>
<connection>
<GID>5302</GID>
<name>N_in1</name></connection>
<intersection>-744.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>277.5,-744.5,277.5,-729.5</points>
<connection>
<GID>3854</GID>
<name>N_in0</name></connection>
<intersection>-744.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>272.5,-744.5,277.5,-744.5</points>
<intersection>272.5 0</intersection>
<intersection>277.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-759.5,241.5,-744</points>
<connection>
<GID>5301</GID>
<name>N_in1</name></connection>
<intersection>-744 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>246.5,-744,246.5,-729</points>
<connection>
<GID>3853</GID>
<name>N_in0</name></connection>
<intersection>-744 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>241.5,-744,246.5,-744</points>
<intersection>241.5 0</intersection>
<intersection>246.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2753</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>265.5,-717,267.5,-717</points>
<connection>
<GID>3850</GID>
<name>OUT</name></connection>
<connection>
<GID>3851</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-720.5,269.5,-720</points>
<connection>
<GID>3851</GID>
<name>IN_0</name></connection>
<intersection>-720.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-720.5,269.5,-720.5</points>
<intersection>255.5 2</intersection>
<intersection>269.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>255.5,-720.5,255.5,-707.5</points>
<intersection>-720.5 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>255.5,-716,259.5,-716</points>
<connection>
<GID>3850</GID>
<name>IN_0</name></connection>
<intersection>255.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>253.5,-707.5,255.5,-707.5</points>
<connection>
<GID>3852</GID>
<name>OUT_0</name></connection>
<intersection>255.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2755</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-620,478,-620</points>
<connection>
<GID>4042</GID>
<name>IN_1</name></connection>
<connection>
<GID>4045</GID>
<name>IN_1</name></connection>
<connection>
<GID>4048</GID>
<name>IN_1</name></connection>
<connection>
<GID>4051</GID>
<name>IN_1</name></connection>
<connection>
<GID>4054</GID>
<name>IN_1</name></connection>
<connection>
<GID>4057</GID>
<name>IN_1</name></connection>
<connection>
<GID>4060</GID>
<name>IN_1</name></connection>
<connection>
<GID>4063</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-620,242,-617.5</points>
<connection>
<GID>3991</GID>
<name>OUT_0</name></connection>
<intersection>-620 1</intersection></vsegment></shape></wire>
<wire>
<ID>2756</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-612.5,465.5,-612.5</points>
<connection>
<GID>3993</GID>
<name>OUT</name></connection>
<connection>
<GID>4044</GID>
<name>clock</name></connection>
<connection>
<GID>4047</GID>
<name>clock</name></connection>
<connection>
<GID>4050</GID>
<name>clock</name></connection>
<connection>
<GID>4053</GID>
<name>clock</name></connection>
<connection>
<GID>4056</GID>
<name>clock</name></connection>
<connection>
<GID>4059</GID>
<name>clock</name></connection>
<connection>
<GID>4062</GID>
<name>clock</name></connection>
<connection>
<GID>4065</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2757</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-636,477.5,-636</points>
<connection>
<GID>4018</GID>
<name>IN_1</name></connection>
<connection>
<GID>4021</GID>
<name>IN_1</name></connection>
<connection>
<GID>4024</GID>
<name>IN_1</name></connection>
<connection>
<GID>4027</GID>
<name>IN_1</name></connection>
<connection>
<GID>4030</GID>
<name>IN_1</name></connection>
<connection>
<GID>4033</GID>
<name>IN_1</name></connection>
<connection>
<GID>4036</GID>
<name>IN_1</name></connection>
<connection>
<GID>4039</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-636,242,-633.5</points>
<connection>
<GID>3995</GID>
<name>OUT_0</name></connection>
<intersection>-636 1</intersection></vsegment></shape></wire>
<wire>
<ID>2758</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-628.5,465,-628.5</points>
<connection>
<GID>3997</GID>
<name>OUT</name></connection>
<connection>
<GID>4020</GID>
<name>clock</name></connection>
<connection>
<GID>4023</GID>
<name>clock</name></connection>
<connection>
<GID>4026</GID>
<name>clock</name></connection>
<connection>
<GID>4029</GID>
<name>clock</name></connection>
<connection>
<GID>4032</GID>
<name>clock</name></connection>
<connection>
<GID>4035</GID>
<name>clock</name></connection>
<connection>
<GID>4038</GID>
<name>clock</name></connection>
<connection>
<GID>4041</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2759</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-645.5,464.5,-645.5</points>
<connection>
<GID>4017</GID>
<name>clock</name></connection>
<connection>
<GID>4014</GID>
<name>clock</name></connection>
<connection>
<GID>4011</GID>
<name>clock</name></connection>
<connection>
<GID>4008</GID>
<name>clock</name></connection>
<connection>
<GID>4005</GID>
<name>clock</name></connection>
<connection>
<GID>4002</GID>
<name>clock</name></connection>
<connection>
<GID>4001</GID>
<name>OUT</name></connection>
<connection>
<GID>3996</GID>
<name>clock</name></connection>
<connection>
<GID>3988</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2760</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-653,477,-653</points>
<connection>
<GID>3986</GID>
<name>IN_1</name></connection>
<connection>
<GID>3992</GID>
<name>IN_1</name></connection>
<connection>
<GID>3998</GID>
<name>IN_1</name></connection>
<connection>
<GID>4003</GID>
<name>IN_1</name></connection>
<connection>
<GID>4006</GID>
<name>IN_1</name></connection>
<connection>
<GID>4009</GID>
<name>IN_1</name></connection>
<connection>
<GID>4012</GID>
<name>IN_1</name></connection>
<connection>
<GID>4015</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-653,242,-650.5</points>
<connection>
<GID>3999</GID>
<name>OUT_0</name></connection>
<intersection>-653 1</intersection></vsegment></shape></wire>
<wire>
<ID>2761</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-662,465,-662</points>
<connection>
<GID>3979</GID>
<name>OUT</name></connection>
<connection>
<GID>3956</GID>
<name>clock</name></connection>
<connection>
<GID>3953</GID>
<name>clock</name></connection>
<connection>
<GID>3950</GID>
<name>clock</name></connection>
<connection>
<GID>3947</GID>
<name>clock</name></connection>
<connection>
<GID>3944</GID>
<name>clock</name></connection>
<connection>
<GID>3941</GID>
<name>clock</name></connection>
<connection>
<GID>3938</GID>
<name>clock</name></connection>
<connection>
<GID>3935</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2762</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,-669.5,477.5,-669.5</points>
<connection>
<GID>3933</GID>
<name>IN_1</name></connection>
<connection>
<GID>3936</GID>
<name>IN_1</name></connection>
<connection>
<GID>3939</GID>
<name>IN_1</name></connection>
<connection>
<GID>3942</GID>
<name>IN_1</name></connection>
<connection>
<GID>3945</GID>
<name>IN_1</name></connection>
<connection>
<GID>3948</GID>
<name>IN_1</name></connection>
<connection>
<GID>3951</GID>
<name>IN_1</name></connection>
<connection>
<GID>3954</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,-669.5,241,-666.5</points>
<connection>
<GID>3978</GID>
<name>OUT_0</name></connection>
<intersection>-669.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2763</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-677.5,464.5,-677.5</points>
<connection>
<GID>3981</GID>
<name>OUT</name></connection>
<connection>
<GID>3932</GID>
<name>clock</name></connection>
<connection>
<GID>3929</GID>
<name>clock</name></connection>
<connection>
<GID>3926</GID>
<name>clock</name></connection>
<connection>
<GID>3923</GID>
<name>clock</name></connection>
<connection>
<GID>3920</GID>
<name>clock</name></connection>
<connection>
<GID>3917</GID>
<name>clock</name></connection>
<connection>
<GID>3914</GID>
<name>clock</name></connection>
<connection>
<GID>3911</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2764</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,-685,477,-685</points>
<connection>
<GID>3909</GID>
<name>IN_1</name></connection>
<connection>
<GID>3912</GID>
<name>IN_1</name></connection>
<connection>
<GID>3915</GID>
<name>IN_1</name></connection>
<connection>
<GID>3918</GID>
<name>IN_1</name></connection>
<connection>
<GID>3921</GID>
<name>IN_1</name></connection>
<connection>
<GID>3924</GID>
<name>IN_1</name></connection>
<connection>
<GID>3927</GID>
<name>IN_1</name></connection>
<connection>
<GID>3930</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,-685,241,-682.5</points>
<connection>
<GID>3980</GID>
<name>OUT_0</name></connection>
<intersection>-685 1</intersection></vsegment></shape></wire>
<wire>
<ID>2765</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297,-717,299,-717</points>
<connection>
<GID>3864</GID>
<name>OUT</name></connection>
<connection>
<GID>3865</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287,-720,301,-720</points>
<connection>
<GID>3865</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287,-720,287,-707.5</points>
<intersection>-720 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287,-716,291,-716</points>
<connection>
<GID>3864</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>284.5,-707.5,287,-707.5</points>
<connection>
<GID>3866</GID>
<name>OUT_0</name></connection>
<intersection>287 2</intersection></hsegment></shape></wire>
<wire>
<ID>2767</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>327.5,-717,329.5,-717</points>
<connection>
<GID>3867</GID>
<name>OUT</name></connection>
<connection>
<GID>3868</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,-720.5,331.5,-720</points>
<connection>
<GID>3868</GID>
<name>IN_0</name></connection>
<intersection>-720.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-720.5,331.5,-720.5</points>
<intersection>317.5 2</intersection>
<intersection>331.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>317.5,-720.5,317.5,-707.5</points>
<intersection>-720.5 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>317.5,-716,321.5,-716</points>
<connection>
<GID>3867</GID>
<name>IN_0</name></connection>
<intersection>317.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>315.5,-707.5,317.5,-707.5</points>
<connection>
<GID>3869</GID>
<name>OUT_0</name></connection>
<intersection>317.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2769</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359,-717,361,-717</points>
<connection>
<GID>3870</GID>
<name>OUT</name></connection>
<connection>
<GID>3871</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,-720,363,-720</points>
<connection>
<GID>3871</GID>
<name>IN_0</name></connection>
<intersection>349 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349,-720,349,-707.5</points>
<intersection>-720 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349,-716,353,-716</points>
<connection>
<GID>3870</GID>
<name>IN_0</name></connection>
<intersection>349 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>346.5,-707.5,349,-707.5</points>
<connection>
<GID>3872</GID>
<name>OUT_0</name></connection>
<intersection>349 2</intersection></hsegment></shape></wire>
<wire>
<ID>2771</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>388.5,-717,390.5,-717</points>
<connection>
<GID>3873</GID>
<name>OUT</name></connection>
<connection>
<GID>3874</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392.5,-720.5,392.5,-720</points>
<connection>
<GID>3874</GID>
<name>IN_0</name></connection>
<intersection>-720.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378.5,-720.5,392.5,-720.5</points>
<intersection>378.5 2</intersection>
<intersection>392.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>378.5,-720.5,378.5,-707.5</points>
<intersection>-720.5 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>378.5,-716,382.5,-716</points>
<connection>
<GID>3873</GID>
<name>IN_0</name></connection>
<intersection>378.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>376.5,-707.5,378.5,-707.5</points>
<connection>
<GID>3875</GID>
<name>OUT_0</name></connection>
<intersection>378.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2773</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420,-717,422,-717</points>
<connection>
<GID>3876</GID>
<name>OUT</name></connection>
<connection>
<GID>3877</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2774</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410,-720,424,-720</points>
<connection>
<GID>3877</GID>
<name>IN_0</name></connection>
<intersection>410 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410,-720,410,-707.5</points>
<intersection>-720 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410,-716,414,-716</points>
<connection>
<GID>3876</GID>
<name>IN_0</name></connection>
<intersection>410 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>407.5,-707.5,410,-707.5</points>
<connection>
<GID>3878</GID>
<name>OUT_0</name></connection>
<intersection>410 2</intersection></hsegment></shape></wire>
<wire>
<ID>2775</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>450.5,-717,452.5,-717</points>
<connection>
<GID>3879</GID>
<name>OUT</name></connection>
<connection>
<GID>3880</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,-720.5,454.5,-720</points>
<connection>
<GID>3880</GID>
<name>IN_0</name></connection>
<intersection>-720.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>440.5,-720.5,454.5,-720.5</points>
<intersection>440.5 2</intersection>
<intersection>454.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>440.5,-720.5,440.5,-707.5</points>
<intersection>-720.5 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>440.5,-716,444.5,-716</points>
<connection>
<GID>3879</GID>
<name>IN_0</name></connection>
<intersection>440.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>438.5,-707.5,440.5,-707.5</points>
<connection>
<GID>3881</GID>
<name>OUT_0</name></connection>
<intersection>440.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2777</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482,-717,484,-717</points>
<connection>
<GID>3882</GID>
<name>OUT</name></connection>
<connection>
<GID>3883</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2778</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472,-720,486,-720</points>
<connection>
<GID>3883</GID>
<name>IN_0</name></connection>
<intersection>472 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472,-720,472,-707.5</points>
<intersection>-720 1</intersection>
<intersection>-716 4</intersection>
<intersection>-707.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472,-716,476,-716</points>
<connection>
<GID>3882</GID>
<name>IN_0</name></connection>
<intersection>472 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>469.5,-707.5,472,-707.5</points>
<connection>
<GID>3884</GID>
<name>OUT_0</name></connection>
<intersection>472 2</intersection></hsegment></shape></wire>
<wire>
<ID>2779</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266,-700,268,-700</points>
<connection>
<GID>3885</GID>
<name>OUT</name></connection>
<connection>
<GID>3886</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-703.5,270,-703</points>
<connection>
<GID>3886</GID>
<name>IN_0</name></connection>
<intersection>-703.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,-703.5,270,-703.5</points>
<intersection>256 2</intersection>
<intersection>270 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256,-703.5,256,-690.5</points>
<intersection>-703.5 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256,-699,260,-699</points>
<connection>
<GID>3885</GID>
<name>IN_0</name></connection>
<intersection>256 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254,-690.5,256,-690.5</points>
<connection>
<GID>3887</GID>
<name>OUT_0</name></connection>
<intersection>256 2</intersection></hsegment></shape></wire>
<wire>
<ID>2781</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>297.5,-700,299.5,-700</points>
<connection>
<GID>3888</GID>
<name>OUT</name></connection>
<connection>
<GID>3889</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2782</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287.5,-703,301.5,-703</points>
<connection>
<GID>3889</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287.5,-703,287.5,-690.5</points>
<intersection>-703 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,-699,291.5,-699</points>
<connection>
<GID>3888</GID>
<name>IN_0</name></connection>
<intersection>287.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285,-690.5,287.5,-690.5</points>
<connection>
<GID>3890</GID>
<name>OUT_0</name></connection>
<intersection>287.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2783</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328,-700,330,-700</points>
<connection>
<GID>3891</GID>
<name>OUT</name></connection>
<connection>
<GID>3892</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,-703.5,332,-703</points>
<connection>
<GID>3892</GID>
<name>IN_0</name></connection>
<intersection>-703.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,-703.5,332,-703.5</points>
<intersection>318 2</intersection>
<intersection>332 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318,-703.5,318,-690.5</points>
<intersection>-703.5 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318,-699,322,-699</points>
<connection>
<GID>3891</GID>
<name>IN_0</name></connection>
<intersection>318 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316,-690.5,318,-690.5</points>
<connection>
<GID>3893</GID>
<name>OUT_0</name></connection>
<intersection>318 2</intersection></hsegment></shape></wire>
<wire>
<ID>2785</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>359.5,-700,361.5,-700</points>
<connection>
<GID>3894</GID>
<name>OUT</name></connection>
<connection>
<GID>3895</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2786</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349.5,-703,363.5,-703</points>
<connection>
<GID>3895</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>349.5,-703,349.5,-690.5</points>
<intersection>-703 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>349.5,-699,353.5,-699</points>
<connection>
<GID>3894</GID>
<name>IN_0</name></connection>
<intersection>349.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347,-690.5,349.5,-690.5</points>
<connection>
<GID>3896</GID>
<name>OUT_0</name></connection>
<intersection>349.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2787</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389,-700,391,-700</points>
<connection>
<GID>3897</GID>
<name>OUT</name></connection>
<connection>
<GID>3898</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,-703.5,393,-703</points>
<connection>
<GID>3898</GID>
<name>IN_0</name></connection>
<intersection>-703.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,-703.5,393,-703.5</points>
<intersection>379 2</intersection>
<intersection>393 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379,-703.5,379,-690.5</points>
<intersection>-703.5 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379,-699,383,-699</points>
<connection>
<GID>3897</GID>
<name>IN_0</name></connection>
<intersection>379 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377,-690.5,379,-690.5</points>
<connection>
<GID>3899</GID>
<name>OUT_0</name></connection>
<intersection>379 2</intersection></hsegment></shape></wire>
<wire>
<ID>2789</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>420.5,-700,422.5,-700</points>
<connection>
<GID>3900</GID>
<name>OUT</name></connection>
<connection>
<GID>3901</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2790</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>410.5,-703,424.5,-703</points>
<connection>
<GID>3901</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>410.5,-703,410.5,-690.5</points>
<intersection>-703 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>410.5,-699,414.5,-699</points>
<connection>
<GID>3900</GID>
<name>IN_0</name></connection>
<intersection>410.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408,-690.5,410.5,-690.5</points>
<connection>
<GID>3902</GID>
<name>OUT_0</name></connection>
<intersection>410.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2791</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451,-700,453,-700</points>
<connection>
<GID>3903</GID>
<name>OUT</name></connection>
<connection>
<GID>3904</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,-703.5,455,-703</points>
<connection>
<GID>3904</GID>
<name>IN_0</name></connection>
<intersection>-703.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,-703.5,455,-703.5</points>
<intersection>441 2</intersection>
<intersection>455 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441,-703.5,441,-690.5</points>
<intersection>-703.5 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441,-699,445,-699</points>
<connection>
<GID>3903</GID>
<name>IN_0</name></connection>
<intersection>441 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439,-690.5,441,-690.5</points>
<connection>
<GID>3905</GID>
<name>OUT_0</name></connection>
<intersection>441 2</intersection></hsegment></shape></wire>
<wire>
<ID>2793</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>482.5,-700,484.5,-700</points>
<connection>
<GID>3906</GID>
<name>OUT</name></connection>
<connection>
<GID>3907</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2794</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>472.5,-703,486.5,-703</points>
<connection>
<GID>3907</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472.5,-703,472.5,-690.5</points>
<intersection>-703 1</intersection>
<intersection>-699 4</intersection>
<intersection>-690.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>472.5,-699,476.5,-699</points>
<connection>
<GID>3906</GID>
<name>IN_0</name></connection>
<intersection>472.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470,-690.5,472.5,-690.5</points>
<connection>
<GID>3908</GID>
<name>OUT_0</name></connection>
<intersection>472.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2795</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266.5,-684,268.5,-684</points>
<connection>
<GID>3909</GID>
<name>OUT</name></connection>
<connection>
<GID>3910</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-687.5,270.5,-687</points>
<connection>
<GID>3910</GID>
<name>IN_0</name></connection>
<intersection>-687.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,-687.5,270.5,-687.5</points>
<intersection>256.5 2</intersection>
<intersection>270.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256.5,-687.5,256.5,-674.5</points>
<intersection>-687.5 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256.5,-683,260.5,-683</points>
<connection>
<GID>3909</GID>
<name>IN_0</name></connection>
<intersection>256.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254.5,-674.5,256.5,-674.5</points>
<connection>
<GID>3911</GID>
<name>OUT_0</name></connection>
<intersection>256.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2797</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,-684,300,-684</points>
<connection>
<GID>3912</GID>
<name>OUT</name></connection>
<connection>
<GID>3913</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2798</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,-687,302,-687</points>
<connection>
<GID>3913</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288,-687,288,-674.5</points>
<intersection>-687 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,-683,292,-683</points>
<connection>
<GID>3912</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285.5,-674.5,288,-674.5</points>
<connection>
<GID>3914</GID>
<name>OUT_0</name></connection>
<intersection>288 2</intersection></hsegment></shape></wire>
<wire>
<ID>2799</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328.5,-684,330.5,-684</points>
<connection>
<GID>3915</GID>
<name>OUT</name></connection>
<connection>
<GID>3916</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-687.5,332.5,-687</points>
<connection>
<GID>3916</GID>
<name>IN_0</name></connection>
<intersection>-687.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-687.5,332.5,-687.5</points>
<intersection>318.5 2</intersection>
<intersection>332.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318.5,-687.5,318.5,-674.5</points>
<intersection>-687.5 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318.5,-683,322.5,-683</points>
<connection>
<GID>3915</GID>
<name>IN_0</name></connection>
<intersection>318.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316.5,-674.5,318.5,-674.5</points>
<connection>
<GID>3917</GID>
<name>OUT_0</name></connection>
<intersection>318.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2801</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360,-684,362,-684</points>
<connection>
<GID>3918</GID>
<name>OUT</name></connection>
<connection>
<GID>3919</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2802</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-687,364,-687</points>
<connection>
<GID>3919</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,-687,350,-674.5</points>
<intersection>-687 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350,-683,354,-683</points>
<connection>
<GID>3918</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347.5,-674.5,350,-674.5</points>
<connection>
<GID>3920</GID>
<name>OUT_0</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>2803</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389.5,-684,391.5,-684</points>
<connection>
<GID>3921</GID>
<name>OUT</name></connection>
<connection>
<GID>3922</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,-687.5,393.5,-687</points>
<connection>
<GID>3922</GID>
<name>IN_0</name></connection>
<intersection>-687.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-687.5,393.5,-687.5</points>
<intersection>379.5 2</intersection>
<intersection>393.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379.5,-687.5,379.5,-674.5</points>
<intersection>-687.5 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379.5,-683,383.5,-683</points>
<connection>
<GID>3921</GID>
<name>IN_0</name></connection>
<intersection>379.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377.5,-674.5,379.5,-674.5</points>
<connection>
<GID>3923</GID>
<name>OUT_0</name></connection>
<intersection>379.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2805</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421,-684,423,-684</points>
<connection>
<GID>3924</GID>
<name>OUT</name></connection>
<connection>
<GID>3925</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2806</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411,-687,425,-687</points>
<connection>
<GID>3925</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411,-687,411,-674.5</points>
<intersection>-687 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411,-683,415,-683</points>
<connection>
<GID>3924</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408.5,-674.5,411,-674.5</points>
<connection>
<GID>3926</GID>
<name>OUT_0</name></connection>
<intersection>411 2</intersection></hsegment></shape></wire>
<wire>
<ID>2807</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451.5,-684,453.5,-684</points>
<connection>
<GID>3927</GID>
<name>OUT</name></connection>
<connection>
<GID>3928</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-687.5,455.5,-687</points>
<connection>
<GID>3928</GID>
<name>IN_0</name></connection>
<intersection>-687.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,-687.5,455.5,-687.5</points>
<intersection>441.5 2</intersection>
<intersection>455.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441.5,-687.5,441.5,-674.5</points>
<intersection>-687.5 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441.5,-683,445.5,-683</points>
<connection>
<GID>3927</GID>
<name>IN_0</name></connection>
<intersection>441.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439.5,-674.5,441.5,-674.5</points>
<connection>
<GID>3929</GID>
<name>OUT_0</name></connection>
<intersection>441.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2809</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483,-684,485,-684</points>
<connection>
<GID>3930</GID>
<name>OUT</name></connection>
<connection>
<GID>3931</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2810</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473,-687,487,-687</points>
<connection>
<GID>3931</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473,-687,473,-674.5</points>
<intersection>-687 1</intersection>
<intersection>-683 4</intersection>
<intersection>-674.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473,-683,477,-683</points>
<connection>
<GID>3930</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470.5,-674.5,473,-674.5</points>
<connection>
<GID>3932</GID>
<name>OUT_0</name></connection>
<intersection>473 2</intersection></hsegment></shape></wire>
<wire>
<ID>2811</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267,-668.5,269,-668.5</points>
<connection>
<GID>3933</GID>
<name>OUT</name></connection>
<connection>
<GID>3934</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-672,271,-671.5</points>
<connection>
<GID>3934</GID>
<name>IN_0</name></connection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-672,271,-672</points>
<intersection>257 2</intersection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257,-672,257,-659</points>
<intersection>-672 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,-667.5,261,-667.5</points>
<connection>
<GID>3933</GID>
<name>IN_0</name></connection>
<intersection>257 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255,-659,257,-659</points>
<connection>
<GID>3935</GID>
<name>OUT_0</name></connection>
<intersection>257 2</intersection></hsegment></shape></wire>
<wire>
<ID>2813</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,-668.5,300.5,-668.5</points>
<connection>
<GID>3936</GID>
<name>OUT</name></connection>
<connection>
<GID>3937</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2814</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288.5,-671.5,302.5,-671.5</points>
<connection>
<GID>3937</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288.5,-671.5,288.5,-659</points>
<intersection>-671.5 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,-667.5,292.5,-667.5</points>
<connection>
<GID>3936</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,-659,288.5,-659</points>
<connection>
<GID>3938</GID>
<name>OUT_0</name></connection>
<intersection>288.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2815</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329,-668.5,331,-668.5</points>
<connection>
<GID>3939</GID>
<name>OUT</name></connection>
<connection>
<GID>3940</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2816</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,-672,333,-671.5</points>
<connection>
<GID>3940</GID>
<name>IN_0</name></connection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-672,333,-672</points>
<intersection>319 2</intersection>
<intersection>333 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319,-672,319,-659</points>
<intersection>-672 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,-667.5,323,-667.5</points>
<connection>
<GID>3939</GID>
<name>IN_0</name></connection>
<intersection>319 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317,-659,319,-659</points>
<connection>
<GID>3941</GID>
<name>OUT_0</name></connection>
<intersection>319 2</intersection></hsegment></shape></wire>
<wire>
<ID>2817</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360.5,-668.5,362.5,-668.5</points>
<connection>
<GID>3942</GID>
<name>OUT</name></connection>
<connection>
<GID>3943</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2818</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350.5,-671.5,364.5,-671.5</points>
<connection>
<GID>3943</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,-671.5,350.5,-659</points>
<intersection>-671.5 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350.5,-667.5,354.5,-667.5</points>
<connection>
<GID>3942</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348,-659,350.5,-659</points>
<connection>
<GID>3944</GID>
<name>OUT_0</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2819</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390,-668.5,392,-668.5</points>
<connection>
<GID>3945</GID>
<name>OUT</name></connection>
<connection>
<GID>3946</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,-672,394,-671.5</points>
<connection>
<GID>3946</GID>
<name>IN_0</name></connection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-672,394,-672</points>
<intersection>380 2</intersection>
<intersection>394 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380,-672,380,-659</points>
<intersection>-672 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,-667.5,384,-667.5</points>
<connection>
<GID>3945</GID>
<name>IN_0</name></connection>
<intersection>380 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378,-659,380,-659</points>
<connection>
<GID>3947</GID>
<name>OUT_0</name></connection>
<intersection>380 2</intersection></hsegment></shape></wire>
<wire>
<ID>2821</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421.5,-668.5,423.5,-668.5</points>
<connection>
<GID>3948</GID>
<name>OUT</name></connection>
<connection>
<GID>3949</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2822</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411.5,-671.5,425.5,-671.5</points>
<connection>
<GID>3949</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411.5,-671.5,411.5,-659</points>
<intersection>-671.5 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411.5,-667.5,415.5,-667.5</points>
<connection>
<GID>3948</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409,-659,411.5,-659</points>
<connection>
<GID>3950</GID>
<name>OUT_0</name></connection>
<intersection>411.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2823</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452,-668.5,454,-668.5</points>
<connection>
<GID>3951</GID>
<name>OUT</name></connection>
<connection>
<GID>3952</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-672,456,-671.5</points>
<connection>
<GID>3952</GID>
<name>IN_0</name></connection>
<intersection>-672 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,-672,456,-672</points>
<intersection>442 2</intersection>
<intersection>456 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442,-672,442,-659</points>
<intersection>-672 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442,-667.5,446,-667.5</points>
<connection>
<GID>3951</GID>
<name>IN_0</name></connection>
<intersection>442 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,-659,442,-659</points>
<connection>
<GID>3953</GID>
<name>OUT_0</name></connection>
<intersection>442 2</intersection></hsegment></shape></wire>
<wire>
<ID>2825</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483.5,-668.5,485.5,-668.5</points>
<connection>
<GID>3954</GID>
<name>OUT</name></connection>
<connection>
<GID>3955</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473.5,-671.5,487.5,-671.5</points>
<connection>
<GID>3955</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473.5,-671.5,473.5,-659</points>
<intersection>-671.5 1</intersection>
<intersection>-667.5 4</intersection>
<intersection>-659 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473.5,-667.5,477.5,-667.5</points>
<connection>
<GID>3954</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471,-659,473.5,-659</points>
<connection>
<GID>3956</GID>
<name>OUT_0</name></connection>
<intersection>473.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2827</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-693.5,464,-693.5</points>
<connection>
<GID>3983</GID>
<name>OUT</name></connection>
<connection>
<GID>3908</GID>
<name>clock</name></connection>
<connection>
<GID>3905</GID>
<name>clock</name></connection>
<connection>
<GID>3902</GID>
<name>clock</name></connection>
<connection>
<GID>3899</GID>
<name>clock</name></connection>
<connection>
<GID>3896</GID>
<name>clock</name></connection>
<connection>
<GID>3893</GID>
<name>clock</name></connection>
<connection>
<GID>3890</GID>
<name>clock</name></connection>
<connection>
<GID>3887</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2828</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,-701,476.5,-701</points>
<connection>
<GID>3885</GID>
<name>IN_1</name></connection>
<connection>
<GID>3888</GID>
<name>IN_1</name></connection>
<connection>
<GID>3891</GID>
<name>IN_1</name></connection>
<connection>
<GID>3894</GID>
<name>IN_1</name></connection>
<connection>
<GID>3897</GID>
<name>IN_1</name></connection>
<connection>
<GID>3900</GID>
<name>IN_1</name></connection>
<connection>
<GID>3903</GID>
<name>IN_1</name></connection>
<connection>
<GID>3906</GID>
<name>IN_1</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,-701,241,-698.5</points>
<connection>
<GID>3982</GID>
<name>OUT_0</name></connection>
<intersection>-701 1</intersection></vsegment></shape></wire>
<wire>
<ID>2829</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-710.5,463.5,-710.5</points>
<connection>
<GID>3985</GID>
<name>OUT</name></connection>
<connection>
<GID>3884</GID>
<name>clock</name></connection>
<connection>
<GID>3881</GID>
<name>clock</name></connection>
<connection>
<GID>3878</GID>
<name>clock</name></connection>
<connection>
<GID>3875</GID>
<name>clock</name></connection>
<connection>
<GID>3872</GID>
<name>clock</name></connection>
<connection>
<GID>3869</GID>
<name>clock</name></connection>
<connection>
<GID>3866</GID>
<name>clock</name></connection>
<connection>
<GID>3852</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-718,242,-715.5</points>
<intersection>-718 2</intersection>
<intersection>-715.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>242,-718,476,-718</points>
<connection>
<GID>3850</GID>
<name>IN_1</name></connection>
<connection>
<GID>3864</GID>
<name>IN_1</name></connection>
<connection>
<GID>3867</GID>
<name>IN_1</name></connection>
<connection>
<GID>3870</GID>
<name>IN_1</name></connection>
<connection>
<GID>3873</GID>
<name>IN_1</name></connection>
<connection>
<GID>3876</GID>
<name>IN_1</name></connection>
<connection>
<GID>3879</GID>
<name>IN_1</name></connection>
<connection>
<GID>3882</GID>
<name>IN_1</name></connection>
<intersection>242 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>241,-715.5,242,-715.5</points>
<connection>
<GID>3984</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>2831</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-727.5,277.5,-587.5</points>
<connection>
<GID>3862</GID>
<name>N_in0</name></connection>
<connection>
<GID>3854</GID>
<name>N_in1</name></connection>
<intersection>-707.5 1</intersection>
<intersection>-690.5 3</intersection>
<intersection>-674.5 4</intersection>
<intersection>-659 5</intersection>
<intersection>-642.5 6</intersection>
<intersection>-625.5 7</intersection>
<intersection>-609.5 8</intersection>
<intersection>-594 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,-707.5,278.5,-707.5</points>
<connection>
<GID>3866</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277.5,-594,281,-594</points>
<connection>
<GID>4071</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>277.5,-690.5,279,-690.5</points>
<connection>
<GID>3890</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>277.5,-674.5,279.5,-674.5</points>
<connection>
<GID>3914</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>277.5,-659,280,-659</points>
<connection>
<GID>3938</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>277.5,-642.5,279.5,-642.5</points>
<connection>
<GID>3996</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>277.5,-625.5,280,-625.5</points>
<connection>
<GID>4023</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>277.5,-609.5,280.5,-609.5</points>
<connection>
<GID>4047</GID>
<name>IN_0</name></connection>
<intersection>277.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-727.5,309.5,-587.5</points>
<connection>
<GID>3863</GID>
<name>N_in0</name></connection>
<connection>
<GID>3869</GID>
<name>IN_0</name></connection>
<connection>
<GID>3855</GID>
<name>N_in1</name></connection>
<intersection>-690.5 9</intersection>
<intersection>-674.5 10</intersection>
<intersection>-659 7</intersection>
<intersection>-642.5 11</intersection>
<intersection>-625.5 5</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309.5,-594,312,-594</points>
<connection>
<GID>4074</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-609.5,311.5,-609.5</points>
<connection>
<GID>4050</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>309.5,-625.5,311,-625.5</points>
<connection>
<GID>4026</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>309.5,-659,311,-659</points>
<connection>
<GID>3941</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>309.5,-690.5,310,-690.5</points>
<connection>
<GID>3893</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>309.5,-674.5,310.5,-674.5</points>
<connection>
<GID>3917</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>309.5,-642.5,310.5,-642.5</points>
<connection>
<GID>4002</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2833</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>340.5,-726.5,340.5,-587.5</points>
<connection>
<GID>3957</GID>
<name>N_in0</name></connection>
<connection>
<GID>3872</GID>
<name>IN_0</name></connection>
<connection>
<GID>3856</GID>
<name>N_in1</name></connection>
<intersection>-690.5 38</intersection>
<intersection>-674.5 21</intersection>
<intersection>-659 7</intersection>
<intersection>-642.5 20</intersection>
<intersection>-625.5 5</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>340.5,-594,343,-594</points>
<connection>
<GID>4077</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>340.5,-609.5,342.5,-609.5</points>
<connection>
<GID>4053</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>340.5,-625.5,342,-625.5</points>
<connection>
<GID>4029</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>340.5,-659,342,-659</points>
<connection>
<GID>3944</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>340.5,-642.5,341.5,-642.5</points>
<connection>
<GID>4005</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>340.5,-674.5,341.5,-674.5</points>
<connection>
<GID>3920</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>340.5,-690.5,341,-690.5</points>
<connection>
<GID>3896</GID>
<name>IN_0</name></connection>
<intersection>340.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2834</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>371.5,-690.5,371.5,-588</points>
<connection>
<GID>4008</GID>
<name>IN_0</name></connection>
<connection>
<GID>3923</GID>
<name>IN_0</name></connection>
<connection>
<GID>3958</GID>
<name>N_in0</name></connection>
<intersection>-690.5 9</intersection>
<intersection>-659 7</intersection>
<intersection>-625.5 5</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>371.5,-594,373,-594</points>
<connection>
<GID>4080</GID>
<name>IN_0</name></connection>
<intersection>371.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>371.5,-609.5,372.5,-609.5</points>
<connection>
<GID>4056</GID>
<name>IN_0</name></connection>
<intersection>371.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>371.5,-625.5,372,-625.5</points>
<connection>
<GID>4032</GID>
<name>IN_0</name></connection>
<intersection>371.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>371.5,-659,372,-659</points>
<connection>
<GID>3947</GID>
<name>IN_0</name></connection>
<intersection>371.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>370.5,-690.5,371.5,-690.5</points>
<connection>
<GID>3899</GID>
<name>IN_0</name></connection>
<intersection>370.5 10</intersection>
<intersection>371.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>370.5,-725.5,370.5,-690.5</points>
<connection>
<GID>3875</GID>
<name>IN_0</name></connection>
<connection>
<GID>3857</GID>
<name>N_in1</name></connection>
<intersection>-690.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>2835</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>401.5,-725,401.5,-587.5</points>
<connection>
<GID>3959</GID>
<name>N_in0</name></connection>
<connection>
<GID>3878</GID>
<name>IN_0</name></connection>
<connection>
<GID>3858</GID>
<name>N_in1</name></connection>
<intersection>-690.5 13</intersection>
<intersection>-674.5 11</intersection>
<intersection>-659 9</intersection>
<intersection>-642.5 7</intersection>
<intersection>-625.5 5</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>401.5,-594,404,-594</points>
<connection>
<GID>4083</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>401.5,-609.5,403.5,-609.5</points>
<connection>
<GID>4059</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>401.5,-625.5,403,-625.5</points>
<connection>
<GID>4035</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>401.5,-642.5,402.5,-642.5</points>
<connection>
<GID>4011</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>401.5,-659,403,-659</points>
<connection>
<GID>3950</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>401.5,-674.5,402.5,-674.5</points>
<connection>
<GID>3926</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>401.5,-690.5,402,-690.5</points>
<connection>
<GID>3902</GID>
<name>IN_0</name></connection>
<intersection>401.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2836</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432.5,-724,432.5,-587.5</points>
<connection>
<GID>3960</GID>
<name>N_in0</name></connection>
<connection>
<GID>3881</GID>
<name>IN_0</name></connection>
<connection>
<GID>3860</GID>
<name>N_in1</name></connection>
<intersection>-690.5 13</intersection>
<intersection>-674.5 11</intersection>
<intersection>-659 9</intersection>
<intersection>-642.5 7</intersection>
<intersection>-625.5 5</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,-594,435,-594</points>
<connection>
<GID>4086</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432.5,-609.5,434.5,-609.5</points>
<connection>
<GID>4062</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>432.5,-625.5,434,-625.5</points>
<connection>
<GID>4038</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>432.5,-642.5,433.5,-642.5</points>
<connection>
<GID>4014</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>432.5,-659,434,-659</points>
<connection>
<GID>3953</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>432.5,-674.5,433.5,-674.5</points>
<connection>
<GID>3929</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>432.5,-690.5,433,-690.5</points>
<connection>
<GID>3905</GID>
<name>IN_0</name></connection>
<intersection>432.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463.5,-726,463.5,-588</points>
<connection>
<GID>3961</GID>
<name>N_in0</name></connection>
<connection>
<GID>3884</GID>
<name>IN_0</name></connection>
<connection>
<GID>3859</GID>
<name>N_in1</name></connection>
<intersection>-690.5 13</intersection>
<intersection>-674.5 10</intersection>
<intersection>-659 8</intersection>
<intersection>-642.5 6</intersection>
<intersection>-625.5 4</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463.5,-594,466,-594</points>
<connection>
<GID>4089</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>463.5,-609.5,465.5,-609.5</points>
<connection>
<GID>4065</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>463.5,-625.5,465,-625.5</points>
<connection>
<GID>4041</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>463.5,-642.5,464.5,-642.5</points>
<connection>
<GID>4017</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>463.5,-659,465,-659</points>
<connection>
<GID>3956</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>463.5,-674.5,464.5,-674.5</points>
<connection>
<GID>3932</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>463.5,-690.5,464,-690.5</points>
<connection>
<GID>3908</GID>
<name>IN_0</name></connection>
<intersection>463.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-735.5,275.5,-580.5</points>
<connection>
<GID>3963</GID>
<name>N_in1</name></connection>
<connection>
<GID>3962</GID>
<name>N_in0</name></connection>
<intersection>-714.5 13</intersection>
<intersection>-697.5 12</intersection>
<intersection>-681.5 11</intersection>
<intersection>-666 10</intersection>
<intersection>-649.5 9</intersection>
<intersection>-632.5 8</intersection>
<intersection>-616.5 7</intersection>
<intersection>-601 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>272,-601,275.5,-601</points>
<connection>
<GID>4067</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>271.5,-616.5,275.5,-616.5</points>
<connection>
<GID>4043</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>271,-632.5,275.5,-632.5</points>
<connection>
<GID>4019</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>270.5,-649.5,275.5,-649.5</points>
<connection>
<GID>3987</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>271,-666,275.5,-666</points>
<connection>
<GID>3934</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>270.5,-681.5,275.5,-681.5</points>
<connection>
<GID>3910</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>270,-697.5,275.5,-697.5</points>
<connection>
<GID>3886</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>269.5,-714.5,275.5,-714.5</points>
<connection>
<GID>3851</GID>
<name>OUT_0</name></connection>
<intersection>275.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306.5,-714.5,306.5,-580.5</points>
<connection>
<GID>3976</GID>
<name>N_in0</name></connection>
<intersection>-714.5 13</intersection>
<intersection>-697.5 12</intersection>
<intersection>-681.5 11</intersection>
<intersection>-666 10</intersection>
<intersection>-649.5 9</intersection>
<intersection>-632.5 8</intersection>
<intersection>-616.5 7</intersection>
<intersection>-601 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>303.5,-601,306.5,-601</points>
<connection>
<GID>4070</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>303,-616.5,306.5,-616.5</points>
<connection>
<GID>4046</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>302.5,-632.5,306.5,-632.5</points>
<connection>
<GID>4022</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>302,-649.5,306.5,-649.5</points>
<connection>
<GID>3994</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>302.5,-666,306.5,-666</points>
<connection>
<GID>3937</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>302,-681.5,306.5,-681.5</points>
<connection>
<GID>3913</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>301.5,-697.5,306.5,-697.5</points>
<connection>
<GID>3889</GID>
<name>OUT_0</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>301,-714.5,306.5,-714.5</points>
<connection>
<GID>3865</GID>
<name>OUT_0</name></connection>
<intersection>304 22</intersection>
<intersection>306.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>304,-729,304,-714.5</points>
<intersection>-729 23</intersection>
<intersection>-714.5 13</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>301.5,-729,304,-729</points>
<connection>
<GID>5785</GID>
<name>N_in1</name></connection>
<intersection>304 22</intersection></hsegment></shape></wire>
<wire>
<ID>2840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,-734.5,338.5,-580.5</points>
<connection>
<GID>3975</GID>
<name>N_in0</name></connection>
<connection>
<GID>3964</GID>
<name>N_in1</name></connection>
<intersection>-714.5 13</intersection>
<intersection>-697.5 12</intersection>
<intersection>-681.5 11</intersection>
<intersection>-666 10</intersection>
<intersection>-649.5 9</intersection>
<intersection>-632.5 8</intersection>
<intersection>-616.5 7</intersection>
<intersection>-601 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>334,-601,338.5,-601</points>
<connection>
<GID>4073</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>333.5,-616.5,338.5,-616.5</points>
<connection>
<GID>4049</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>333,-632.5,338.5,-632.5</points>
<connection>
<GID>4025</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>332.5,-649.5,338.5,-649.5</points>
<connection>
<GID>4000</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>333,-666,338.5,-666</points>
<connection>
<GID>3940</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>332.5,-681.5,338.5,-681.5</points>
<connection>
<GID>3916</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>332,-697.5,338.5,-697.5</points>
<connection>
<GID>3892</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>331.5,-714.5,338.5,-714.5</points>
<connection>
<GID>3868</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369,-734,369,-580.5</points>
<connection>
<GID>3974</GID>
<name>N_in0</name></connection>
<connection>
<GID>3965</GID>
<name>N_in1</name></connection>
<intersection>-714.5 18</intersection>
<intersection>-697.5 17</intersection>
<intersection>-681.5 16</intersection>
<intersection>-666 15</intersection>
<intersection>-649.5 14</intersection>
<intersection>-632.5 13</intersection>
<intersection>-616.5 12</intersection>
<intersection>-601 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>365.5,-601,369,-601</points>
<connection>
<GID>4076</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>365,-616.5,369,-616.5</points>
<connection>
<GID>4052</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>364.5,-632.5,369,-632.5</points>
<connection>
<GID>4028</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>364,-649.5,369,-649.5</points>
<connection>
<GID>4004</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>364.5,-666,369,-666</points>
<connection>
<GID>3943</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>364,-681.5,369,-681.5</points>
<connection>
<GID>3919</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>363.5,-697.5,369,-697.5</points>
<connection>
<GID>3895</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>363,-714.5,369,-714.5</points>
<connection>
<GID>3871</GID>
<name>OUT_0</name></connection>
<intersection>369 0</intersection></hsegment></shape></wire>
<wire>
<ID>2842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,-734,399.5,-580.5</points>
<connection>
<GID>3973</GID>
<name>N_in0</name></connection>
<connection>
<GID>3966</GID>
<name>N_in1</name></connection>
<intersection>-714.5 9</intersection>
<intersection>-697.5 10</intersection>
<intersection>-681.5 11</intersection>
<intersection>-666 12</intersection>
<intersection>-649.5 13</intersection>
<intersection>-632.5 14</intersection>
<intersection>-616.5 15</intersection>
<intersection>-601 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>392.5,-714.5,399.5,-714.5</points>
<connection>
<GID>3874</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>393,-697.5,399.5,-697.5</points>
<connection>
<GID>3898</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>393.5,-681.5,399.5,-681.5</points>
<connection>
<GID>3922</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>394,-666,399.5,-666</points>
<connection>
<GID>3946</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>393.5,-649.5,399.5,-649.5</points>
<connection>
<GID>4007</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>394,-632.5,399.5,-632.5</points>
<connection>
<GID>4031</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>394.5,-616.5,399.5,-616.5</points>
<connection>
<GID>4055</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>395,-601,399.5,-601</points>
<connection>
<GID>4079</GID>
<name>OUT_0</name></connection>
<intersection>399.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2843</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,-734,430.5,-580.5</points>
<connection>
<GID>3972</GID>
<name>N_in0</name></connection>
<connection>
<GID>3967</GID>
<name>N_in1</name></connection>
<intersection>-714.5 6</intersection>
<intersection>-697.5 7</intersection>
<intersection>-681.5 8</intersection>
<intersection>-666 9</intersection>
<intersection>-649.5 10</intersection>
<intersection>-632.5 11</intersection>
<intersection>-616.5 12</intersection>
<intersection>-601 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>424,-714.5,430.5,-714.5</points>
<connection>
<GID>3877</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>424.5,-697.5,430.5,-697.5</points>
<connection>
<GID>3901</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>425,-681.5,430.5,-681.5</points>
<connection>
<GID>3925</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>425.5,-666,430.5,-666</points>
<connection>
<GID>3949</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>425,-649.5,430.5,-649.5</points>
<connection>
<GID>4010</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>425.5,-632.5,430.5,-632.5</points>
<connection>
<GID>4034</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>426,-616.5,430.5,-616.5</points>
<connection>
<GID>4058</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>426.5,-601,430.5,-601</points>
<connection>
<GID>4082</GID>
<name>OUT_0</name></connection>
<intersection>430.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461.5,-734.5,461.5,-579.5</points>
<connection>
<GID>3971</GID>
<name>N_in0</name></connection>
<connection>
<GID>3968</GID>
<name>N_in1</name></connection>
<intersection>-714.5 6</intersection>
<intersection>-697.5 7</intersection>
<intersection>-681.5 8</intersection>
<intersection>-666 9</intersection>
<intersection>-649.5 10</intersection>
<intersection>-632.5 11</intersection>
<intersection>-616.5 12</intersection>
<intersection>-601 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>454.5,-714.5,461.5,-714.5</points>
<connection>
<GID>3880</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>455,-697.5,461.5,-697.5</points>
<connection>
<GID>3904</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>455.5,-681.5,461.5,-681.5</points>
<connection>
<GID>3928</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>456,-666,461.5,-666</points>
<connection>
<GID>3952</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>455.5,-649.5,461.5,-649.5</points>
<connection>
<GID>4013</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>456,-632.5,461.5,-632.5</points>
<connection>
<GID>4037</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>456.5,-616.5,461.5,-616.5</points>
<connection>
<GID>4061</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>457,-601,461.5,-601</points>
<connection>
<GID>4085</GID>
<name>OUT_0</name></connection>
<intersection>461.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492,-734,492,-579</points>
<connection>
<GID>3970</GID>
<name>N_in0</name></connection>
<connection>
<GID>3969</GID>
<name>N_in1</name></connection>
<intersection>-714.5 3</intersection>
<intersection>-697.5 4</intersection>
<intersection>-681.5 5</intersection>
<intersection>-666 6</intersection>
<intersection>-649.5 7</intersection>
<intersection>-632.5 8</intersection>
<intersection>-616.5 9</intersection>
<intersection>-601 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>486,-714.5,492,-714.5</points>
<connection>
<GID>3883</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>486.5,-697.5,492,-697.5</points>
<connection>
<GID>3907</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>487,-681.5,492,-681.5</points>
<connection>
<GID>3931</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>487.5,-666,492,-666</points>
<connection>
<GID>3955</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>487,-649.5,492,-649.5</points>
<connection>
<GID>4016</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>487.5,-632.5,492,-632.5</points>
<connection>
<GID>4040</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>488,-616.5,492,-616.5</points>
<connection>
<GID>4064</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>488.5,-601,492,-601</points>
<connection>
<GID>4088</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment></shape></wire>
<wire>
<ID>2846</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,-648.5,200.5,-599.5</points>
<intersection>-648.5 2</intersection>
<intersection>-599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,-599.5,239.5,-599.5</points>
<connection>
<GID>3989</GID>
<name>ENABLE_0</name></connection>
<intersection>200.5 0</intersection>
<intersection>225.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-648.5,200.5,-648.5</points>
<connection>
<GID>3977</GID>
<name>OUT_7</name></connection>
<intersection>200.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-599.5,225.5,-596</points>
<intersection>-599.5 1</intersection>
<intersection>-596 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-596,230,-596</points>
<connection>
<GID>3990</GID>
<name>IN_0</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-649.5,202.5,-615</points>
<intersection>-649.5 2</intersection>
<intersection>-615 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-615,239.5,-615</points>
<intersection>202.5 0</intersection>
<intersection>225.5 4</intersection>
<intersection>239.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-649.5,202.5,-649.5</points>
<connection>
<GID>3977</GID>
<name>OUT_6</name></connection>
<intersection>202.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239.5,-615.5,239.5,-615</points>
<connection>
<GID>3991</GID>
<name>ENABLE_0</name></connection>
<intersection>-615 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-615,225.5,-611.5</points>
<intersection>-615 1</intersection>
<intersection>-611.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-611.5,229.5,-611.5</points>
<connection>
<GID>3993</GID>
<name>IN_0</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-650.5,204.5,-627.5</points>
<intersection>-650.5 2</intersection>
<intersection>-627.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-627.5,229.5,-627.5</points>
<connection>
<GID>3997</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection>
<intersection>225.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-650.5,204.5,-650.5</points>
<connection>
<GID>3977</GID>
<name>OUT_5</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>225.5,-631.5,225.5,-627.5</points>
<intersection>-631.5 4</intersection>
<intersection>-627.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>225.5,-631.5,239.5,-631.5</points>
<connection>
<GID>3995</GID>
<name>ENABLE_0</name></connection>
<intersection>225.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-651.5,206.5,-644.5</points>
<intersection>-651.5 2</intersection>
<intersection>-644.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,-644.5,229.5,-644.5</points>
<connection>
<GID>4001</GID>
<name>IN_0</name></connection>
<intersection>206.5 0</intersection>
<intersection>225.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-651.5,206.5,-651.5</points>
<connection>
<GID>3977</GID>
<name>OUT_4</name></connection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>225.5,-648.5,225.5,-644.5</points>
<intersection>-648.5 4</intersection>
<intersection>-644.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>225.5,-648.5,239.5,-648.5</points>
<connection>
<GID>3999</GID>
<name>ENABLE_0</name></connection>
<intersection>225.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2850</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-664.5,206.5,-652.5</points>
<intersection>-664.5 1</intersection>
<intersection>-652.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,-664.5,238.5,-664.5</points>
<connection>
<GID>3978</GID>
<name>ENABLE_0</name></connection>
<intersection>206.5 0</intersection>
<intersection>225.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-652.5,206.5,-652.5</points>
<connection>
<GID>3977</GID>
<name>OUT_3</name></connection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-664.5,225.5,-661</points>
<intersection>-664.5 1</intersection>
<intersection>-661 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-661,229.5,-661</points>
<connection>
<GID>3979</GID>
<name>IN_0</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2851</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-680.5,204.5,-653.5</points>
<intersection>-680.5 1</intersection>
<intersection>-653.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-680.5,238.5,-680.5</points>
<connection>
<GID>3980</GID>
<name>ENABLE_0</name></connection>
<intersection>204.5 0</intersection>
<intersection>225.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-653.5,204.5,-653.5</points>
<connection>
<GID>3977</GID>
<name>OUT_2</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-680.5,225.5,-676.5</points>
<intersection>-680.5 1</intersection>
<intersection>-676.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-676.5,229.5,-676.5</points>
<connection>
<GID>3981</GID>
<name>IN_0</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2852</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-696,202.5,-654.5</points>
<intersection>-696 1</intersection>
<intersection>-654.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-696,238.5,-696</points>
<intersection>202.5 0</intersection>
<intersection>225.5 4</intersection>
<intersection>238.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-654.5,202.5,-654.5</points>
<connection>
<GID>3977</GID>
<name>OUT_1</name></connection>
<intersection>202.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>238.5,-696.5,238.5,-696</points>
<connection>
<GID>3982</GID>
<name>ENABLE_0</name></connection>
<intersection>-696 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-696,225.5,-692.5</points>
<intersection>-696 1</intersection>
<intersection>-692.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-692.5,229.5,-692.5</points>
<connection>
<GID>3983</GID>
<name>IN_0</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2853</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,-713.5,200.5,-655.5</points>
<intersection>-713.5 1</intersection>
<intersection>-655.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,-713.5,238.5,-713.5</points>
<connection>
<GID>3984</GID>
<name>ENABLE_0</name></connection>
<intersection>200.5 0</intersection>
<intersection>225.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-655.5,200.5,-655.5</points>
<connection>
<GID>3977</GID>
<name>OUT_0</name></connection>
<intersection>200.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-713.5,225.5,-709.5</points>
<intersection>-713.5 1</intersection>
<intersection>-709.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-709.5,229.5,-709.5</points>
<connection>
<GID>3985</GID>
<name>IN_0</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2854</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>266.5,-652,268.5,-652</points>
<connection>
<GID>3986</GID>
<name>OUT</name></connection>
<connection>
<GID>3987</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2855</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-655.5,270.5,-655</points>
<connection>
<GID>3987</GID>
<name>IN_0</name></connection>
<intersection>-655.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,-655.5,270.5,-655.5</points>
<intersection>256.5 2</intersection>
<intersection>270.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>256.5,-655.5,256.5,-642.5</points>
<intersection>-655.5 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>256.5,-651,260.5,-651</points>
<connection>
<GID>3986</GID>
<name>IN_0</name></connection>
<intersection>256.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>254.5,-642.5,256.5,-642.5</points>
<connection>
<GID>3988</GID>
<name>OUT_0</name></connection>
<intersection>256.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2856</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,-652,300,-652</points>
<connection>
<GID>3992</GID>
<name>OUT</name></connection>
<connection>
<GID>3994</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2857</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,-655,302,-655</points>
<connection>
<GID>3994</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288,-655,288,-642.5</points>
<intersection>-655 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,-651,292,-651</points>
<connection>
<GID>3992</GID>
<name>IN_0</name></connection>
<intersection>288 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>285.5,-642.5,288,-642.5</points>
<connection>
<GID>3996</GID>
<name>OUT_0</name></connection>
<intersection>288 2</intersection></hsegment></shape></wire>
<wire>
<ID>2858</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>328.5,-652,330.5,-652</points>
<connection>
<GID>3998</GID>
<name>OUT</name></connection>
<connection>
<GID>4000</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2859</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-655.5,332.5,-655</points>
<connection>
<GID>4000</GID>
<name>IN_0</name></connection>
<intersection>-655.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-655.5,332.5,-655.5</points>
<intersection>318.5 2</intersection>
<intersection>332.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>318.5,-655.5,318.5,-642.5</points>
<intersection>-655.5 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>318.5,-651,322.5,-651</points>
<connection>
<GID>3998</GID>
<name>IN_0</name></connection>
<intersection>318.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>316.5,-642.5,318.5,-642.5</points>
<connection>
<GID>4002</GID>
<name>OUT_0</name></connection>
<intersection>318.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2860</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360,-652,362,-652</points>
<connection>
<GID>4003</GID>
<name>OUT</name></connection>
<connection>
<GID>4004</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2861</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350,-655,364,-655</points>
<connection>
<GID>4004</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,-655,350,-642.5</points>
<intersection>-655 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350,-651,354,-651</points>
<connection>
<GID>4003</GID>
<name>IN_0</name></connection>
<intersection>350 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>347.5,-642.5,350,-642.5</points>
<connection>
<GID>4005</GID>
<name>OUT_0</name></connection>
<intersection>350 2</intersection></hsegment></shape></wire>
<wire>
<ID>2862</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>389.5,-652,391.5,-652</points>
<connection>
<GID>4006</GID>
<name>OUT</name></connection>
<connection>
<GID>4007</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2863</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,-655.5,393.5,-655</points>
<connection>
<GID>4007</GID>
<name>IN_0</name></connection>
<intersection>-655.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-655.5,393.5,-655.5</points>
<intersection>379.5 2</intersection>
<intersection>393.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>379.5,-655.5,379.5,-642.5</points>
<intersection>-655.5 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>379.5,-651,383.5,-651</points>
<connection>
<GID>4006</GID>
<name>IN_0</name></connection>
<intersection>379.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>377.5,-642.5,379.5,-642.5</points>
<connection>
<GID>4008</GID>
<name>OUT_0</name></connection>
<intersection>379.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2864</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421,-652,423,-652</points>
<connection>
<GID>4009</GID>
<name>OUT</name></connection>
<connection>
<GID>4010</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2865</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411,-655,425,-655</points>
<connection>
<GID>4010</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411,-655,411,-642.5</points>
<intersection>-655 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411,-651,415,-651</points>
<connection>
<GID>4009</GID>
<name>IN_0</name></connection>
<intersection>411 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>408.5,-642.5,411,-642.5</points>
<connection>
<GID>4011</GID>
<name>OUT_0</name></connection>
<intersection>411 2</intersection></hsegment></shape></wire>
<wire>
<ID>2866</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>451.5,-652,453.5,-652</points>
<connection>
<GID>4012</GID>
<name>OUT</name></connection>
<connection>
<GID>4013</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-655.5,455.5,-655</points>
<connection>
<GID>4013</GID>
<name>IN_0</name></connection>
<intersection>-655.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,-655.5,455.5,-655.5</points>
<intersection>441.5 2</intersection>
<intersection>455.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>441.5,-655.5,441.5,-642.5</points>
<intersection>-655.5 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>441.5,-651,445.5,-651</points>
<connection>
<GID>4012</GID>
<name>IN_0</name></connection>
<intersection>441.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>439.5,-642.5,441.5,-642.5</points>
<connection>
<GID>4014</GID>
<name>OUT_0</name></connection>
<intersection>441.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2868</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483,-652,485,-652</points>
<connection>
<GID>4015</GID>
<name>OUT</name></connection>
<connection>
<GID>4016</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2869</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473,-655,487,-655</points>
<connection>
<GID>4016</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473,-655,473,-642.5</points>
<intersection>-655 1</intersection>
<intersection>-651 4</intersection>
<intersection>-642.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473,-651,477,-651</points>
<connection>
<GID>4015</GID>
<name>IN_0</name></connection>
<intersection>473 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>470.5,-642.5,473,-642.5</points>
<connection>
<GID>4017</GID>
<name>OUT_0</name></connection>
<intersection>473 2</intersection></hsegment></shape></wire>
<wire>
<ID>2870</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267,-635,269,-635</points>
<connection>
<GID>4018</GID>
<name>OUT</name></connection>
<connection>
<GID>4019</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2871</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-638.5,271,-638</points>
<connection>
<GID>4019</GID>
<name>IN_0</name></connection>
<intersection>-638.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-638.5,271,-638.5</points>
<intersection>257 2</intersection>
<intersection>271 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257,-638.5,257,-625.5</points>
<intersection>-638.5 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,-634,261,-634</points>
<connection>
<GID>4018</GID>
<name>IN_0</name></connection>
<intersection>257 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255,-625.5,257,-625.5</points>
<connection>
<GID>4020</GID>
<name>OUT_0</name></connection>
<intersection>257 2</intersection></hsegment></shape></wire>
<wire>
<ID>2872</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,-635,300.5,-635</points>
<connection>
<GID>4021</GID>
<name>OUT</name></connection>
<connection>
<GID>4022</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2873</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288.5,-638,302.5,-638</points>
<connection>
<GID>4022</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>288.5,-638,288.5,-625.5</points>
<intersection>-638 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,-634,292.5,-634</points>
<connection>
<GID>4021</GID>
<name>IN_0</name></connection>
<intersection>288.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,-625.5,288.5,-625.5</points>
<connection>
<GID>4023</GID>
<name>OUT_0</name></connection>
<intersection>288.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2874</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329,-635,331,-635</points>
<connection>
<GID>4024</GID>
<name>OUT</name></connection>
<connection>
<GID>4025</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,-638.5,333,-638</points>
<connection>
<GID>4025</GID>
<name>IN_0</name></connection>
<intersection>-638.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-638.5,333,-638.5</points>
<intersection>319 2</intersection>
<intersection>333 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319,-638.5,319,-625.5</points>
<intersection>-638.5 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,-634,323,-634</points>
<connection>
<GID>4024</GID>
<name>IN_0</name></connection>
<intersection>319 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317,-625.5,319,-625.5</points>
<connection>
<GID>4026</GID>
<name>OUT_0</name></connection>
<intersection>319 2</intersection></hsegment></shape></wire>
<wire>
<ID>2876</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>360.5,-635,362.5,-635</points>
<connection>
<GID>4027</GID>
<name>OUT</name></connection>
<connection>
<GID>4028</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2877</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>350.5,-638,364.5,-638</points>
<connection>
<GID>4028</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350.5,-638,350.5,-625.5</points>
<intersection>-638 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>350.5,-634,354.5,-634</points>
<connection>
<GID>4027</GID>
<name>IN_0</name></connection>
<intersection>350.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348,-625.5,350.5,-625.5</points>
<connection>
<GID>4029</GID>
<name>OUT_0</name></connection>
<intersection>350.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2878</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390,-635,392,-635</points>
<connection>
<GID>4030</GID>
<name>OUT</name></connection>
<connection>
<GID>4031</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,-638.5,394,-638</points>
<connection>
<GID>4031</GID>
<name>IN_0</name></connection>
<intersection>-638.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-638.5,394,-638.5</points>
<intersection>380 2</intersection>
<intersection>394 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380,-638.5,380,-625.5</points>
<intersection>-638.5 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,-634,384,-634</points>
<connection>
<GID>4030</GID>
<name>IN_0</name></connection>
<intersection>380 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378,-625.5,380,-625.5</points>
<connection>
<GID>4032</GID>
<name>OUT_0</name></connection>
<intersection>380 2</intersection></hsegment></shape></wire>
<wire>
<ID>2880</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>421.5,-635,423.5,-635</points>
<connection>
<GID>4033</GID>
<name>OUT</name></connection>
<connection>
<GID>4034</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2881</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>411.5,-638,425.5,-638</points>
<connection>
<GID>4034</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411.5,-638,411.5,-625.5</points>
<intersection>-638 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>411.5,-634,415.5,-634</points>
<connection>
<GID>4033</GID>
<name>IN_0</name></connection>
<intersection>411.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409,-625.5,411.5,-625.5</points>
<connection>
<GID>4035</GID>
<name>OUT_0</name></connection>
<intersection>411.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2882</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452,-635,454,-635</points>
<connection>
<GID>4036</GID>
<name>OUT</name></connection>
<connection>
<GID>4037</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2883</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-638.5,456,-638</points>
<connection>
<GID>4037</GID>
<name>IN_0</name></connection>
<intersection>-638.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,-638.5,456,-638.5</points>
<intersection>442 2</intersection>
<intersection>456 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442,-638.5,442,-625.5</points>
<intersection>-638.5 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442,-634,446,-634</points>
<connection>
<GID>4036</GID>
<name>IN_0</name></connection>
<intersection>442 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,-625.5,442,-625.5</points>
<connection>
<GID>4038</GID>
<name>OUT_0</name></connection>
<intersection>442 2</intersection></hsegment></shape></wire>
<wire>
<ID>2884</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>483.5,-635,485.5,-635</points>
<connection>
<GID>4039</GID>
<name>OUT</name></connection>
<connection>
<GID>4040</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2885</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>473.5,-638,487.5,-638</points>
<connection>
<GID>4040</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473.5,-638,473.5,-625.5</points>
<intersection>-638 1</intersection>
<intersection>-634 4</intersection>
<intersection>-625.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>473.5,-634,477.5,-634</points>
<connection>
<GID>4039</GID>
<name>IN_0</name></connection>
<intersection>473.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471,-625.5,473.5,-625.5</points>
<connection>
<GID>4041</GID>
<name>OUT_0</name></connection>
<intersection>473.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2886</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>267.5,-619,269.5,-619</points>
<connection>
<GID>4042</GID>
<name>OUT</name></connection>
<connection>
<GID>4043</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2887</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-622.5,271.5,-622</points>
<connection>
<GID>4043</GID>
<name>IN_0</name></connection>
<intersection>-622.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-622.5,271.5,-622.5</points>
<intersection>257.5 2</intersection>
<intersection>271.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>257.5,-622.5,257.5,-609.5</points>
<intersection>-622.5 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257.5,-618,261.5,-618</points>
<connection>
<GID>4042</GID>
<name>IN_0</name></connection>
<intersection>257.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>255.5,-609.5,257.5,-609.5</points>
<connection>
<GID>4044</GID>
<name>OUT_0</name></connection>
<intersection>257.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2888</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299,-619,301,-619</points>
<connection>
<GID>4045</GID>
<name>OUT</name></connection>
<connection>
<GID>4046</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2889</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-622,303,-622</points>
<connection>
<GID>4046</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289,-622,289,-609.5</points>
<intersection>-622 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289,-618,293,-618</points>
<connection>
<GID>4045</GID>
<name>IN_0</name></connection>
<intersection>289 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286.5,-609.5,289,-609.5</points>
<connection>
<GID>4047</GID>
<name>OUT_0</name></connection>
<intersection>289 2</intersection></hsegment></shape></wire>
<wire>
<ID>2890</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>329.5,-619,331.5,-619</points>
<connection>
<GID>4048</GID>
<name>OUT</name></connection>
<connection>
<GID>4049</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,-622.5,333.5,-622</points>
<connection>
<GID>4049</GID>
<name>IN_0</name></connection>
<intersection>-622.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-622.5,333.5,-622.5</points>
<intersection>319.5 2</intersection>
<intersection>333.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>319.5,-622.5,319.5,-609.5</points>
<intersection>-622.5 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319.5,-618,323.5,-618</points>
<connection>
<GID>4048</GID>
<name>IN_0</name></connection>
<intersection>319.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>317.5,-609.5,319.5,-609.5</points>
<connection>
<GID>4050</GID>
<name>OUT_0</name></connection>
<intersection>319.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2892</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361,-619,363,-619</points>
<connection>
<GID>4051</GID>
<name>OUT</name></connection>
<connection>
<GID>4052</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2893</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351,-622,365,-622</points>
<connection>
<GID>4052</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351,-622,351,-609.5</points>
<intersection>-622 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351,-618,355,-618</points>
<connection>
<GID>4051</GID>
<name>IN_0</name></connection>
<intersection>351 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348.5,-609.5,351,-609.5</points>
<connection>
<GID>4053</GID>
<name>OUT_0</name></connection>
<intersection>351 2</intersection></hsegment></shape></wire>
<wire>
<ID>2894</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>390.5,-619,392.5,-619</points>
<connection>
<GID>4054</GID>
<name>OUT</name></connection>
<connection>
<GID>4055</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2895</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394.5,-622.5,394.5,-622</points>
<connection>
<GID>4055</GID>
<name>IN_0</name></connection>
<intersection>-622.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,-622.5,394.5,-622.5</points>
<intersection>380.5 2</intersection>
<intersection>394.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>380.5,-622.5,380.5,-609.5</points>
<intersection>-622.5 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380.5,-618,384.5,-618</points>
<connection>
<GID>4054</GID>
<name>IN_0</name></connection>
<intersection>380.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>378.5,-609.5,380.5,-609.5</points>
<connection>
<GID>4056</GID>
<name>OUT_0</name></connection>
<intersection>380.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2896</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422,-619,424,-619</points>
<connection>
<GID>4057</GID>
<name>OUT</name></connection>
<connection>
<GID>4058</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2897</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,-622,426,-622</points>
<connection>
<GID>4058</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412,-622,412,-609.5</points>
<intersection>-622 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412,-618,416,-618</points>
<connection>
<GID>4057</GID>
<name>IN_0</name></connection>
<intersection>412 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>409.5,-609.5,412,-609.5</points>
<connection>
<GID>4059</GID>
<name>OUT_0</name></connection>
<intersection>412 2</intersection></hsegment></shape></wire>
<wire>
<ID>2898</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>452.5,-619,454.5,-619</points>
<connection>
<GID>4060</GID>
<name>OUT</name></connection>
<connection>
<GID>4061</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2899</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-622.5,456.5,-622</points>
<connection>
<GID>4061</GID>
<name>IN_0</name></connection>
<intersection>-622.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,-622.5,456.5,-622.5</points>
<intersection>442.5 2</intersection>
<intersection>456.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>442.5,-622.5,442.5,-609.5</points>
<intersection>-622.5 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>442.5,-618,446.5,-618</points>
<connection>
<GID>4060</GID>
<name>IN_0</name></connection>
<intersection>442.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,-609.5,442.5,-609.5</points>
<connection>
<GID>4062</GID>
<name>OUT_0</name></connection>
<intersection>442.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2900</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484,-619,486,-619</points>
<connection>
<GID>4063</GID>
<name>OUT</name></connection>
<connection>
<GID>4064</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2901</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474,-622,488,-622</points>
<connection>
<GID>4064</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474,-622,474,-609.5</points>
<intersection>-622 1</intersection>
<intersection>-618 4</intersection>
<intersection>-609.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474,-618,478,-618</points>
<connection>
<GID>4063</GID>
<name>IN_0</name></connection>
<intersection>474 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>471.5,-609.5,474,-609.5</points>
<connection>
<GID>4065</GID>
<name>OUT_0</name></connection>
<intersection>474 2</intersection></hsegment></shape></wire>
<wire>
<ID>2902</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>268,-603.5,270,-603.5</points>
<connection>
<GID>4066</GID>
<name>OUT</name></connection>
<connection>
<GID>4067</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2903</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-607,272,-606.5</points>
<connection>
<GID>4067</GID>
<name>IN_0</name></connection>
<intersection>-607 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-607,272,-607</points>
<intersection>258 2</intersection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,-607,258,-594</points>
<intersection>-607 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258,-602.5,262,-602.5</points>
<connection>
<GID>4066</GID>
<name>IN_0</name></connection>
<intersection>258 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>256,-594,258,-594</points>
<connection>
<GID>4068</GID>
<name>OUT_0</name></connection>
<intersection>258 2</intersection></hsegment></shape></wire>
<wire>
<ID>2904</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>299.5,-603.5,301.5,-603.5</points>
<connection>
<GID>4069</GID>
<name>OUT</name></connection>
<connection>
<GID>4070</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2905</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289.5,-606.5,303.5,-606.5</points>
<connection>
<GID>4070</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>289.5,-606.5,289.5,-594</points>
<intersection>-606.5 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>289.5,-602.5,293.5,-602.5</points>
<connection>
<GID>4069</GID>
<name>IN_0</name></connection>
<intersection>289.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287,-594,289.5,-594</points>
<connection>
<GID>4071</GID>
<name>OUT_0</name></connection>
<intersection>289.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2906</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>330,-603.5,332,-603.5</points>
<connection>
<GID>4072</GID>
<name>OUT</name></connection>
<connection>
<GID>4073</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2907</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-607,334,-606.5</points>
<connection>
<GID>4073</GID>
<name>IN_0</name></connection>
<intersection>-607 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-607,334,-607</points>
<intersection>320 2</intersection>
<intersection>334 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>320,-607,320,-594</points>
<intersection>-607 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>320,-602.5,324,-602.5</points>
<connection>
<GID>4072</GID>
<name>IN_0</name></connection>
<intersection>320 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>318,-594,320,-594</points>
<connection>
<GID>4074</GID>
<name>OUT_0</name></connection>
<intersection>320 2</intersection></hsegment></shape></wire>
<wire>
<ID>2908</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>361.5,-603.5,363.5,-603.5</points>
<connection>
<GID>4075</GID>
<name>OUT</name></connection>
<connection>
<GID>4076</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2909</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>351.5,-606.5,365.5,-606.5</points>
<connection>
<GID>4076</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>351.5,-606.5,351.5,-594</points>
<intersection>-606.5 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>351.5,-602.5,355.5,-602.5</points>
<connection>
<GID>4075</GID>
<name>IN_0</name></connection>
<intersection>351.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>349,-594,351.5,-594</points>
<connection>
<GID>4077</GID>
<name>OUT_0</name></connection>
<intersection>351.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2910</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>391,-603.5,393,-603.5</points>
<connection>
<GID>4078</GID>
<name>OUT</name></connection>
<connection>
<GID>4079</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395,-607,395,-606.5</points>
<connection>
<GID>4079</GID>
<name>IN_0</name></connection>
<intersection>-607 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-607,395,-607</points>
<intersection>381 2</intersection>
<intersection>395 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>381,-607,381,-594</points>
<intersection>-607 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>381,-602.5,385,-602.5</points>
<connection>
<GID>4078</GID>
<name>IN_0</name></connection>
<intersection>381 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>379,-594,381,-594</points>
<connection>
<GID>4080</GID>
<name>OUT_0</name></connection>
<intersection>381 2</intersection></hsegment></shape></wire>
<wire>
<ID>2912</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>422.5,-603.5,424.5,-603.5</points>
<connection>
<GID>4081</GID>
<name>OUT</name></connection>
<connection>
<GID>4082</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2913</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,-606.5,426.5,-606.5</points>
<connection>
<GID>4082</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412.5,-606.5,412.5,-594</points>
<intersection>-606.5 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412.5,-602.5,416.5,-602.5</points>
<connection>
<GID>4081</GID>
<name>IN_0</name></connection>
<intersection>412.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>410,-594,412.5,-594</points>
<connection>
<GID>4083</GID>
<name>OUT_0</name></connection>
<intersection>412.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2914</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>453,-603.5,455,-603.5</points>
<connection>
<GID>4084</GID>
<name>OUT</name></connection>
<connection>
<GID>4085</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-607,457,-606.5</points>
<connection>
<GID>4085</GID>
<name>IN_0</name></connection>
<intersection>-607 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443,-607,457,-607</points>
<intersection>443 2</intersection>
<intersection>457 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>443,-607,443,-594</points>
<intersection>-607 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>443,-602.5,447,-602.5</points>
<connection>
<GID>4084</GID>
<name>IN_0</name></connection>
<intersection>443 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>441,-594,443,-594</points>
<connection>
<GID>4086</GID>
<name>OUT_0</name></connection>
<intersection>443 2</intersection></hsegment></shape></wire>
<wire>
<ID>2916</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>484.5,-603.5,486.5,-603.5</points>
<connection>
<GID>4087</GID>
<name>OUT</name></connection>
<connection>
<GID>4088</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2917</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>474.5,-606.5,488.5,-606.5</points>
<connection>
<GID>4088</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>474.5,-606.5,474.5,-594</points>
<intersection>-606.5 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>474.5,-602.5,478.5,-602.5</points>
<connection>
<GID>4087</GID>
<name>IN_0</name></connection>
<intersection>474.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>472,-594,474.5,-594</points>
<connection>
<GID>4089</GID>
<name>OUT_0</name></connection>
<intersection>474.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-727,246.5,-587.5</points>
<connection>
<GID>3861</GID>
<name>N_in0</name></connection>
<connection>
<GID>3853</GID>
<name>N_in1</name></connection>
<intersection>-707.5 14</intersection>
<intersection>-690.5 12</intersection>
<intersection>-674.5 10</intersection>
<intersection>-659 8</intersection>
<intersection>-642.5 6</intersection>
<intersection>-625.5 4</intersection>
<intersection>-609.5 2</intersection>
<intersection>-594 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246.5,-594,250,-594</points>
<connection>
<GID>4068</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>246.5,-609.5,249.5,-609.5</points>
<connection>
<GID>4044</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>246.5,-625.5,249,-625.5</points>
<connection>
<GID>4020</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>246.5,-642.5,248.5,-642.5</points>
<connection>
<GID>3988</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>246.5,-659,249,-659</points>
<connection>
<GID>3935</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>246.5,-674.5,248.5,-674.5</points>
<connection>
<GID>3911</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>246.5,-690.5,248,-690.5</points>
<connection>
<GID>3887</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>246.5,-707.5,247.5,-707.5</points>
<connection>
<GID>3852</GID>
<name>IN_0</name></connection>
<intersection>246.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2919</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-604.5,478.5,-604.5</points>
<connection>
<GID>4066</GID>
<name>IN_1</name></connection>
<connection>
<GID>4069</GID>
<name>IN_1</name></connection>
<connection>
<GID>4072</GID>
<name>IN_1</name></connection>
<connection>
<GID>4075</GID>
<name>IN_1</name></connection>
<connection>
<GID>4078</GID>
<name>IN_1</name></connection>
<connection>
<GID>4081</GID>
<name>IN_1</name></connection>
<connection>
<GID>4084</GID>
<name>IN_1</name></connection>
<connection>
<GID>4087</GID>
<name>IN_1</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,-604.5,242,-601.5</points>
<connection>
<GID>3989</GID>
<name>OUT_0</name></connection>
<intersection>-604.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2920</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236,-597,466,-597</points>
<connection>
<GID>3990</GID>
<name>OUT</name></connection>
<connection>
<GID>4068</GID>
<name>clock</name></connection>
<connection>
<GID>4071</GID>
<name>clock</name></connection>
<connection>
<GID>4074</GID>
<name>clock</name></connection>
<connection>
<GID>4077</GID>
<name>clock</name></connection>
<connection>
<GID>4080</GID>
<name>clock</name></connection>
<connection>
<GID>4083</GID>
<name>clock</name></connection>
<connection>
<GID>4086</GID>
<name>clock</name></connection>
<connection>
<GID>4089</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2921</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>269.5,22,271.5,22</points>
<connection>
<GID>4090</GID>
<name>OUT</name></connection>
<connection>
<GID>4091</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,18.5,273.5,19</points>
<connection>
<GID>4091</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,18.5,273.5,18.5</points>
<intersection>259.5 2</intersection>
<intersection>273.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>259.5,18.5,259.5,31.5</points>
<intersection>18.5 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,23,263.5,23</points>
<connection>
<GID>4090</GID>
<name>IN_0</name></connection>
<intersection>259.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>257.5,31.5,259.5,31.5</points>
<connection>
<GID>4092</GID>
<name>OUT_0</name></connection>
<intersection>259.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2923</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,119,482,119</points>
<connection>
<GID>4282</GID>
<name>IN_1</name></connection>
<connection>
<GID>4285</GID>
<name>IN_1</name></connection>
<connection>
<GID>4288</GID>
<name>IN_1</name></connection>
<connection>
<GID>4291</GID>
<name>IN_1</name></connection>
<connection>
<GID>4294</GID>
<name>IN_1</name></connection>
<connection>
<GID>4297</GID>
<name>IN_1</name></connection>
<connection>
<GID>4300</GID>
<name>IN_1</name></connection>
<connection>
<GID>4303</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,119,246,121.5</points>
<connection>
<GID>4231</GID>
<name>OUT_0</name></connection>
<intersection>119 1</intersection></vsegment></shape></wire>
<wire>
<ID>2924</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,126.5,469.5,126.5</points>
<connection>
<GID>4233</GID>
<name>OUT</name></connection>
<connection>
<GID>4284</GID>
<name>clock</name></connection>
<connection>
<GID>4287</GID>
<name>clock</name></connection>
<connection>
<GID>4290</GID>
<name>clock</name></connection>
<connection>
<GID>4293</GID>
<name>clock</name></connection>
<connection>
<GID>4296</GID>
<name>clock</name></connection>
<connection>
<GID>4299</GID>
<name>clock</name></connection>
<connection>
<GID>4302</GID>
<name>clock</name></connection>
<connection>
<GID>4305</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2925</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,103,481.5,103</points>
<connection>
<GID>4258</GID>
<name>IN_1</name></connection>
<connection>
<GID>4261</GID>
<name>IN_1</name></connection>
<connection>
<GID>4264</GID>
<name>IN_1</name></connection>
<connection>
<GID>4267</GID>
<name>IN_1</name></connection>
<connection>
<GID>4270</GID>
<name>IN_1</name></connection>
<connection>
<GID>4273</GID>
<name>IN_1</name></connection>
<connection>
<GID>4276</GID>
<name>IN_1</name></connection>
<connection>
<GID>4279</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,103,246,105.5</points>
<connection>
<GID>4235</GID>
<name>OUT_0</name></connection>
<intersection>103 1</intersection></vsegment></shape></wire>
<wire>
<ID>2926</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,110.5,469,110.5</points>
<connection>
<GID>4237</GID>
<name>OUT</name></connection>
<connection>
<GID>4260</GID>
<name>clock</name></connection>
<connection>
<GID>4263</GID>
<name>clock</name></connection>
<connection>
<GID>4266</GID>
<name>clock</name></connection>
<connection>
<GID>4269</GID>
<name>clock</name></connection>
<connection>
<GID>4272</GID>
<name>clock</name></connection>
<connection>
<GID>4275</GID>
<name>clock</name></connection>
<connection>
<GID>4278</GID>
<name>clock</name></connection>
<connection>
<GID>4281</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2927</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,93.5,468.5,93.5</points>
<connection>
<GID>4257</GID>
<name>clock</name></connection>
<connection>
<GID>4254</GID>
<name>clock</name></connection>
<connection>
<GID>4251</GID>
<name>clock</name></connection>
<connection>
<GID>4248</GID>
<name>clock</name></connection>
<connection>
<GID>4245</GID>
<name>clock</name></connection>
<connection>
<GID>4242</GID>
<name>clock</name></connection>
<connection>
<GID>4241</GID>
<name>OUT</name></connection>
<connection>
<GID>4236</GID>
<name>clock</name></connection>
<connection>
<GID>4228</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246,86,481,86</points>
<connection>
<GID>4226</GID>
<name>IN_1</name></connection>
<connection>
<GID>4232</GID>
<name>IN_1</name></connection>
<connection>
<GID>4238</GID>
<name>IN_1</name></connection>
<connection>
<GID>4243</GID>
<name>IN_1</name></connection>
<connection>
<GID>4246</GID>
<name>IN_1</name></connection>
<connection>
<GID>4249</GID>
<name>IN_1</name></connection>
<connection>
<GID>4252</GID>
<name>IN_1</name></connection>
<connection>
<GID>4255</GID>
<name>IN_1</name></connection>
<intersection>246 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>246,86,246,88.5</points>
<connection>
<GID>4239</GID>
<name>OUT_0</name></connection>
<intersection>86 1</intersection></vsegment></shape></wire>
<wire>
<ID>2929</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,77,469,77</points>
<connection>
<GID>4219</GID>
<name>OUT</name></connection>
<connection>
<GID>4196</GID>
<name>clock</name></connection>
<connection>
<GID>4193</GID>
<name>clock</name></connection>
<connection>
<GID>4190</GID>
<name>clock</name></connection>
<connection>
<GID>4187</GID>
<name>clock</name></connection>
<connection>
<GID>4184</GID>
<name>clock</name></connection>
<connection>
<GID>4181</GID>
<name>clock</name></connection>
<connection>
<GID>4178</GID>
<name>clock</name></connection>
<connection>
<GID>4175</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2930</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,69.5,481.5,69.5</points>
<connection>
<GID>4173</GID>
<name>IN_1</name></connection>
<connection>
<GID>4176</GID>
<name>IN_1</name></connection>
<connection>
<GID>4179</GID>
<name>IN_1</name></connection>
<connection>
<GID>4182</GID>
<name>IN_1</name></connection>
<connection>
<GID>4185</GID>
<name>IN_1</name></connection>
<connection>
<GID>4188</GID>
<name>IN_1</name></connection>
<connection>
<GID>4191</GID>
<name>IN_1</name></connection>
<connection>
<GID>4194</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,69.5,245,72.5</points>
<connection>
<GID>4218</GID>
<name>OUT_0</name></connection>
<intersection>69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2931</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,61.5,468.5,61.5</points>
<connection>
<GID>4221</GID>
<name>OUT</name></connection>
<connection>
<GID>4172</GID>
<name>clock</name></connection>
<connection>
<GID>4169</GID>
<name>clock</name></connection>
<connection>
<GID>4166</GID>
<name>clock</name></connection>
<connection>
<GID>4163</GID>
<name>clock</name></connection>
<connection>
<GID>4160</GID>
<name>clock</name></connection>
<connection>
<GID>4157</GID>
<name>clock</name></connection>
<connection>
<GID>4154</GID>
<name>clock</name></connection>
<connection>
<GID>4151</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2932</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,54,481,54</points>
<connection>
<GID>4149</GID>
<name>IN_1</name></connection>
<connection>
<GID>4152</GID>
<name>IN_1</name></connection>
<connection>
<GID>4155</GID>
<name>IN_1</name></connection>
<connection>
<GID>4158</GID>
<name>IN_1</name></connection>
<connection>
<GID>4161</GID>
<name>IN_1</name></connection>
<connection>
<GID>4164</GID>
<name>IN_1</name></connection>
<connection>
<GID>4167</GID>
<name>IN_1</name></connection>
<connection>
<GID>4170</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,54,245,56.5</points>
<connection>
<GID>4220</GID>
<name>OUT_0</name></connection>
<intersection>54 1</intersection></vsegment></shape></wire>
<wire>
<ID>2933</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301,22,303,22</points>
<connection>
<GID>4104</GID>
<name>OUT</name></connection>
<connection>
<GID>4105</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2934</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291,19,305,19</points>
<connection>
<GID>4105</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291,19,291,31.5</points>
<intersection>19 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291,23,295,23</points>
<connection>
<GID>4104</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>288.5,31.5,291,31.5</points>
<connection>
<GID>4106</GID>
<name>OUT_0</name></connection>
<intersection>291 2</intersection></hsegment></shape></wire>
<wire>
<ID>2935</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>331.5,22,333.5,22</points>
<connection>
<GID>4107</GID>
<name>OUT</name></connection>
<connection>
<GID>4108</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,18.5,335.5,19</points>
<connection>
<GID>4108</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,18.5,335.5,18.5</points>
<intersection>321.5 2</intersection>
<intersection>335.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321.5,18.5,321.5,31.5</points>
<intersection>18.5 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321.5,23,325.5,23</points>
<connection>
<GID>4107</GID>
<name>IN_0</name></connection>
<intersection>321.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>319.5,31.5,321.5,31.5</points>
<connection>
<GID>4109</GID>
<name>OUT_0</name></connection>
<intersection>321.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2937</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363,22,365,22</points>
<connection>
<GID>4110</GID>
<name>OUT</name></connection>
<connection>
<GID>4111</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2938</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353,19,367,19</points>
<connection>
<GID>4111</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353,19,353,31.5</points>
<intersection>19 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353,23,357,23</points>
<connection>
<GID>4110</GID>
<name>IN_0</name></connection>
<intersection>353 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>350.5,31.5,353,31.5</points>
<connection>
<GID>4112</GID>
<name>OUT_0</name></connection>
<intersection>353 2</intersection></hsegment></shape></wire>
<wire>
<ID>2939</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>392.5,22,394.5,22</points>
<connection>
<GID>4113</GID>
<name>OUT</name></connection>
<connection>
<GID>4114</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,18.5,396.5,19</points>
<connection>
<GID>4114</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382.5,18.5,396.5,18.5</points>
<intersection>382.5 2</intersection>
<intersection>396.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>382.5,18.5,382.5,31.5</points>
<intersection>18.5 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>382.5,23,386.5,23</points>
<connection>
<GID>4113</GID>
<name>IN_0</name></connection>
<intersection>382.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>380.5,31.5,382.5,31.5</points>
<connection>
<GID>4115</GID>
<name>OUT_0</name></connection>
<intersection>382.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2941</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424,22,426,22</points>
<connection>
<GID>4116</GID>
<name>OUT</name></connection>
<connection>
<GID>4117</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414,19,428,19</points>
<connection>
<GID>4117</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414,19,414,31.5</points>
<intersection>19 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414,23,418,23</points>
<connection>
<GID>4116</GID>
<name>IN_0</name></connection>
<intersection>414 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>411.5,31.5,414,31.5</points>
<connection>
<GID>4118</GID>
<name>OUT_0</name></connection>
<intersection>414 2</intersection></hsegment></shape></wire>
<wire>
<ID>2943</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>454.5,22,456.5,22</points>
<connection>
<GID>4119</GID>
<name>OUT</name></connection>
<connection>
<GID>4120</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,18.5,458.5,19</points>
<connection>
<GID>4120</GID>
<name>IN_0</name></connection>
<intersection>18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,18.5,458.5,18.5</points>
<intersection>444.5 2</intersection>
<intersection>458.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>444.5,18.5,444.5,31.5</points>
<intersection>18.5 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>444.5,23,448.5,23</points>
<connection>
<GID>4119</GID>
<name>IN_0</name></connection>
<intersection>444.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>442.5,31.5,444.5,31.5</points>
<connection>
<GID>4121</GID>
<name>OUT_0</name></connection>
<intersection>444.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2945</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486,22,488,22</points>
<connection>
<GID>4122</GID>
<name>OUT</name></connection>
<connection>
<GID>4123</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2946</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476,19,490,19</points>
<connection>
<GID>4123</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476,19,476,31.5</points>
<intersection>19 1</intersection>
<intersection>23 4</intersection>
<intersection>31.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476,23,480,23</points>
<connection>
<GID>4122</GID>
<name>IN_0</name></connection>
<intersection>476 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>473.5,31.5,476,31.5</points>
<connection>
<GID>4124</GID>
<name>OUT_0</name></connection>
<intersection>476 2</intersection></hsegment></shape></wire>
<wire>
<ID>2947</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270,39,272,39</points>
<connection>
<GID>4125</GID>
<name>OUT</name></connection>
<connection>
<GID>4126</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,35.5,274,36</points>
<connection>
<GID>4126</GID>
<name>IN_0</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,35.5,274,35.5</points>
<intersection>260 2</intersection>
<intersection>274 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260,35.5,260,48.5</points>
<intersection>35.5 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260,40,264,40</points>
<connection>
<GID>4125</GID>
<name>IN_0</name></connection>
<intersection>260 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258,48.5,260,48.5</points>
<connection>
<GID>4127</GID>
<name>OUT_0</name></connection>
<intersection>260 2</intersection></hsegment></shape></wire>
<wire>
<ID>2949</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,39,303.5,39</points>
<connection>
<GID>4128</GID>
<name>OUT</name></connection>
<connection>
<GID>4129</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2950</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>291.5,36,305.5,36</points>
<connection>
<GID>4129</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>291.5,36,291.5,48.5</points>
<intersection>36 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>291.5,40,295.5,40</points>
<connection>
<GID>4128</GID>
<name>IN_0</name></connection>
<intersection>291.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289,48.5,291.5,48.5</points>
<connection>
<GID>4130</GID>
<name>OUT_0</name></connection>
<intersection>291.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2951</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332,39,334,39</points>
<connection>
<GID>4131</GID>
<name>OUT</name></connection>
<connection>
<GID>4132</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,35.5,336,36</points>
<connection>
<GID>4132</GID>
<name>IN_0</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,35.5,336,35.5</points>
<intersection>322 2</intersection>
<intersection>336 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322,35.5,322,48.5</points>
<intersection>35.5 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322,40,326,40</points>
<connection>
<GID>4131</GID>
<name>IN_0</name></connection>
<intersection>322 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320,48.5,322,48.5</points>
<connection>
<GID>4133</GID>
<name>OUT_0</name></connection>
<intersection>322 2</intersection></hsegment></shape></wire>
<wire>
<ID>2953</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>363.5,39,365.5,39</points>
<connection>
<GID>4134</GID>
<name>OUT</name></connection>
<connection>
<GID>4135</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2954</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353.5,36,367.5,36</points>
<connection>
<GID>4135</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>353.5,36,353.5,48.5</points>
<intersection>36 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>353.5,40,357.5,40</points>
<connection>
<GID>4134</GID>
<name>IN_0</name></connection>
<intersection>353.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351,48.5,353.5,48.5</points>
<connection>
<GID>4136</GID>
<name>OUT_0</name></connection>
<intersection>353.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2955</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393,39,395,39</points>
<connection>
<GID>4137</GID>
<name>OUT</name></connection>
<connection>
<GID>4138</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,35.5,397,36</points>
<connection>
<GID>4138</GID>
<name>IN_0</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383,35.5,397,35.5</points>
<intersection>383 2</intersection>
<intersection>397 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,35.5,383,48.5</points>
<intersection>35.5 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383,40,387,40</points>
<connection>
<GID>4137</GID>
<name>IN_0</name></connection>
<intersection>383 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381,48.5,383,48.5</points>
<connection>
<GID>4139</GID>
<name>OUT_0</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>2957</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>424.5,39,426.5,39</points>
<connection>
<GID>4140</GID>
<name>OUT</name></connection>
<connection>
<GID>4141</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2958</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414.5,36,428.5,36</points>
<connection>
<GID>4141</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>414.5,36,414.5,48.5</points>
<intersection>36 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>414.5,40,418.5,40</points>
<connection>
<GID>4140</GID>
<name>IN_0</name></connection>
<intersection>414.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412,48.5,414.5,48.5</points>
<connection>
<GID>4142</GID>
<name>OUT_0</name></connection>
<intersection>414.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2959</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455,39,457,39</points>
<connection>
<GID>4143</GID>
<name>OUT</name></connection>
<connection>
<GID>4144</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,35.5,459,36</points>
<connection>
<GID>4144</GID>
<name>IN_0</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,35.5,459,35.5</points>
<intersection>445 2</intersection>
<intersection>459 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445,35.5,445,48.5</points>
<intersection>35.5 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445,40,449,40</points>
<connection>
<GID>4143</GID>
<name>IN_0</name></connection>
<intersection>445 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443,48.5,445,48.5</points>
<connection>
<GID>4145</GID>
<name>OUT_0</name></connection>
<intersection>445 2</intersection></hsegment></shape></wire>
<wire>
<ID>2961</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>486.5,39,488.5,39</points>
<connection>
<GID>4146</GID>
<name>OUT</name></connection>
<connection>
<GID>4147</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2962</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476.5,36,490.5,36</points>
<connection>
<GID>4147</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>476.5,36,476.5,48.5</points>
<intersection>36 1</intersection>
<intersection>40 4</intersection>
<intersection>48.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>476.5,40,480.5,40</points>
<connection>
<GID>4146</GID>
<name>IN_0</name></connection>
<intersection>476.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474,48.5,476.5,48.5</points>
<connection>
<GID>4148</GID>
<name>OUT_0</name></connection>
<intersection>476.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2963</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270.5,55,272.5,55</points>
<connection>
<GID>4149</GID>
<name>OUT</name></connection>
<connection>
<GID>4150</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,51.5,274.5,52</points>
<connection>
<GID>4150</GID>
<name>IN_0</name></connection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,51.5,274.5,51.5</points>
<intersection>260.5 2</intersection>
<intersection>274.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260.5,51.5,260.5,64.5</points>
<intersection>51.5 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,56,264.5,56</points>
<connection>
<GID>4149</GID>
<name>IN_0</name></connection>
<intersection>260.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258.5,64.5,260.5,64.5</points>
<connection>
<GID>4151</GID>
<name>OUT_0</name></connection>
<intersection>260.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2965</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302,55,304,55</points>
<connection>
<GID>4152</GID>
<name>OUT</name></connection>
<connection>
<GID>4153</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,52,306,52</points>
<connection>
<GID>4153</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292,52,292,64.5</points>
<intersection>52 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292,56,296,56</points>
<connection>
<GID>4152</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289.5,64.5,292,64.5</points>
<connection>
<GID>4154</GID>
<name>OUT_0</name></connection>
<intersection>292 2</intersection></hsegment></shape></wire>
<wire>
<ID>2967</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332.5,55,334.5,55</points>
<connection>
<GID>4155</GID>
<name>OUT</name></connection>
<connection>
<GID>4156</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,51.5,336.5,52</points>
<connection>
<GID>4156</GID>
<name>IN_0</name></connection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,51.5,336.5,51.5</points>
<intersection>322.5 2</intersection>
<intersection>336.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322.5,51.5,322.5,64.5</points>
<intersection>51.5 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322.5,56,326.5,56</points>
<connection>
<GID>4155</GID>
<name>IN_0</name></connection>
<intersection>322.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320.5,64.5,322.5,64.5</points>
<connection>
<GID>4157</GID>
<name>OUT_0</name></connection>
<intersection>322.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2969</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364,55,366,55</points>
<connection>
<GID>4158</GID>
<name>OUT</name></connection>
<connection>
<GID>4159</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2970</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354,52,368,52</points>
<connection>
<GID>4159</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354,52,354,64.5</points>
<intersection>52 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354,56,358,56</points>
<connection>
<GID>4158</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351.5,64.5,354,64.5</points>
<connection>
<GID>4160</GID>
<name>OUT_0</name></connection>
<intersection>354 2</intersection></hsegment></shape></wire>
<wire>
<ID>2971</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393.5,55,395.5,55</points>
<connection>
<GID>4161</GID>
<name>OUT</name></connection>
<connection>
<GID>4162</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,51.5,397.5,52</points>
<connection>
<GID>4162</GID>
<name>IN_0</name></connection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,51.5,397.5,51.5</points>
<intersection>383.5 2</intersection>
<intersection>397.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,51.5,383.5,64.5</points>
<intersection>51.5 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383.5,56,387.5,56</points>
<connection>
<GID>4161</GID>
<name>IN_0</name></connection>
<intersection>383.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381.5,64.5,383.5,64.5</points>
<connection>
<GID>4163</GID>
<name>OUT_0</name></connection>
<intersection>383.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2973</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425,55,427,55</points>
<connection>
<GID>4164</GID>
<name>OUT</name></connection>
<connection>
<GID>4165</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415,52,429,52</points>
<connection>
<GID>4165</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415,52,415,64.5</points>
<intersection>52 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415,56,419,56</points>
<connection>
<GID>4164</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412.5,64.5,415,64.5</points>
<connection>
<GID>4166</GID>
<name>OUT_0</name></connection>
<intersection>415 2</intersection></hsegment></shape></wire>
<wire>
<ID>2975</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455.5,55,457.5,55</points>
<connection>
<GID>4167</GID>
<name>OUT</name></connection>
<connection>
<GID>4168</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,51.5,459.5,52</points>
<connection>
<GID>4168</GID>
<name>IN_0</name></connection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,51.5,459.5,51.5</points>
<intersection>445.5 2</intersection>
<intersection>459.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445.5,51.5,445.5,64.5</points>
<intersection>51.5 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445.5,56,449.5,56</points>
<connection>
<GID>4167</GID>
<name>IN_0</name></connection>
<intersection>445.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443.5,64.5,445.5,64.5</points>
<connection>
<GID>4169</GID>
<name>OUT_0</name></connection>
<intersection>445.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2977</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487,55,489,55</points>
<connection>
<GID>4170</GID>
<name>OUT</name></connection>
<connection>
<GID>4171</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2978</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,52,491,52</points>
<connection>
<GID>4171</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477,52,477,64.5</points>
<intersection>52 1</intersection>
<intersection>56 4</intersection>
<intersection>64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477,56,481,56</points>
<connection>
<GID>4170</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474.5,64.5,477,64.5</points>
<connection>
<GID>4172</GID>
<name>OUT_0</name></connection>
<intersection>477 2</intersection></hsegment></shape></wire>
<wire>
<ID>2979</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271,70.5,273,70.5</points>
<connection>
<GID>4173</GID>
<name>OUT</name></connection>
<connection>
<GID>4174</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,67,275,67.5</points>
<connection>
<GID>4174</GID>
<name>IN_0</name></connection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,67,275,67</points>
<intersection>261 2</intersection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261,67,261,80</points>
<intersection>67 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,71.5,265,71.5</points>
<connection>
<GID>4173</GID>
<name>IN_0</name></connection>
<intersection>261 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259,80,261,80</points>
<connection>
<GID>4175</GID>
<name>OUT_0</name></connection>
<intersection>261 2</intersection></hsegment></shape></wire>
<wire>
<ID>2981</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302.5,70.5,304.5,70.5</points>
<connection>
<GID>4176</GID>
<name>OUT</name></connection>
<connection>
<GID>4177</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2982</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,67.5,306.5,67.5</points>
<connection>
<GID>4177</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292.5,67.5,292.5,80</points>
<intersection>67.5 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292.5,71.5,296.5,71.5</points>
<connection>
<GID>4176</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290,80,292.5,80</points>
<connection>
<GID>4178</GID>
<name>OUT_0</name></connection>
<intersection>292.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2983</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333,70.5,335,70.5</points>
<connection>
<GID>4179</GID>
<name>OUT</name></connection>
<connection>
<GID>4180</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,67,337,67.5</points>
<connection>
<GID>4180</GID>
<name>IN_0</name></connection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,67,337,67</points>
<intersection>323 2</intersection>
<intersection>337 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323,67,323,80</points>
<intersection>67 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323,71.5,327,71.5</points>
<connection>
<GID>4179</GID>
<name>IN_0</name></connection>
<intersection>323 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321,80,323,80</points>
<connection>
<GID>4181</GID>
<name>OUT_0</name></connection>
<intersection>323 2</intersection></hsegment></shape></wire>
<wire>
<ID>2985</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364.5,70.5,366.5,70.5</points>
<connection>
<GID>4182</GID>
<name>OUT</name></connection>
<connection>
<GID>4183</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2986</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,67.5,368.5,67.5</points>
<connection>
<GID>4183</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354.5,67.5,354.5,80</points>
<intersection>67.5 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354.5,71.5,358.5,71.5</points>
<connection>
<GID>4182</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352,80,354.5,80</points>
<connection>
<GID>4184</GID>
<name>OUT_0</name></connection>
<intersection>354.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2987</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394,70.5,396,70.5</points>
<connection>
<GID>4185</GID>
<name>OUT</name></connection>
<connection>
<GID>4186</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,67,398,67.5</points>
<connection>
<GID>4186</GID>
<name>IN_0</name></connection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,67,398,67</points>
<intersection>384 2</intersection>
<intersection>398 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384,67,384,80</points>
<intersection>67 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384,71.5,388,71.5</points>
<connection>
<GID>4185</GID>
<name>IN_0</name></connection>
<intersection>384 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382,80,384,80</points>
<connection>
<GID>4187</GID>
<name>OUT_0</name></connection>
<intersection>384 2</intersection></hsegment></shape></wire>
<wire>
<ID>2989</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425.5,70.5,427.5,70.5</points>
<connection>
<GID>4188</GID>
<name>OUT</name></connection>
<connection>
<GID>4189</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2990</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415.5,67.5,429.5,67.5</points>
<connection>
<GID>4189</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415.5,67.5,415.5,80</points>
<intersection>67.5 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415.5,71.5,419.5,71.5</points>
<connection>
<GID>4188</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413,80,415.5,80</points>
<connection>
<GID>4190</GID>
<name>OUT_0</name></connection>
<intersection>415.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2991</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456,70.5,458,70.5</points>
<connection>
<GID>4191</GID>
<name>OUT</name></connection>
<connection>
<GID>4192</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460,67,460,67.5</points>
<connection>
<GID>4192</GID>
<name>IN_0</name></connection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446,67,460,67</points>
<intersection>446 2</intersection>
<intersection>460 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446,67,446,80</points>
<intersection>67 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446,71.5,450,71.5</points>
<connection>
<GID>4191</GID>
<name>IN_0</name></connection>
<intersection>446 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444,80,446,80</points>
<connection>
<GID>4193</GID>
<name>OUT_0</name></connection>
<intersection>446 2</intersection></hsegment></shape></wire>
<wire>
<ID>2993</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487.5,70.5,489.5,70.5</points>
<connection>
<GID>4194</GID>
<name>OUT</name></connection>
<connection>
<GID>4195</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2994</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,67.5,491.5,67.5</points>
<connection>
<GID>4195</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477.5,67.5,477.5,80</points>
<intersection>67.5 1</intersection>
<intersection>71.5 4</intersection>
<intersection>80 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477.5,71.5,481.5,71.5</points>
<connection>
<GID>4194</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475,80,477.5,80</points>
<connection>
<GID>4196</GID>
<name>OUT_0</name></connection>
<intersection>477.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2995</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,45.5,468,45.5</points>
<connection>
<GID>4223</GID>
<name>OUT</name></connection>
<connection>
<GID>4148</GID>
<name>clock</name></connection>
<connection>
<GID>4145</GID>
<name>clock</name></connection>
<connection>
<GID>4142</GID>
<name>clock</name></connection>
<connection>
<GID>4139</GID>
<name>clock</name></connection>
<connection>
<GID>4136</GID>
<name>clock</name></connection>
<connection>
<GID>4133</GID>
<name>clock</name></connection>
<connection>
<GID>4130</GID>
<name>clock</name></connection>
<connection>
<GID>4127</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2996</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,38,480.5,38</points>
<connection>
<GID>4125</GID>
<name>IN_1</name></connection>
<connection>
<GID>4128</GID>
<name>IN_1</name></connection>
<connection>
<GID>4131</GID>
<name>IN_1</name></connection>
<connection>
<GID>4134</GID>
<name>IN_1</name></connection>
<connection>
<GID>4137</GID>
<name>IN_1</name></connection>
<connection>
<GID>4140</GID>
<name>IN_1</name></connection>
<connection>
<GID>4143</GID>
<name>IN_1</name></connection>
<connection>
<GID>4146</GID>
<name>IN_1</name></connection>
<intersection>245 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245,38,245,40.5</points>
<connection>
<GID>4222</GID>
<name>OUT_0</name></connection>
<intersection>38 1</intersection></vsegment></shape></wire>
<wire>
<ID>2997</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,28.5,467.5,28.5</points>
<connection>
<GID>4225</GID>
<name>OUT</name></connection>
<connection>
<GID>4124</GID>
<name>clock</name></connection>
<connection>
<GID>4121</GID>
<name>clock</name></connection>
<connection>
<GID>4118</GID>
<name>clock</name></connection>
<connection>
<GID>4115</GID>
<name>clock</name></connection>
<connection>
<GID>4112</GID>
<name>clock</name></connection>
<connection>
<GID>4109</GID>
<name>clock</name></connection>
<connection>
<GID>4106</GID>
<name>clock</name></connection>
<connection>
<GID>4092</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>2998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,21,246,23.5</points>
<intersection>21 2</intersection>
<intersection>23.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>246,21,480,21</points>
<connection>
<GID>4090</GID>
<name>IN_1</name></connection>
<connection>
<GID>4104</GID>
<name>IN_1</name></connection>
<connection>
<GID>4107</GID>
<name>IN_1</name></connection>
<connection>
<GID>4110</GID>
<name>IN_1</name></connection>
<connection>
<GID>4113</GID>
<name>IN_1</name></connection>
<connection>
<GID>4116</GID>
<name>IN_1</name></connection>
<connection>
<GID>4119</GID>
<name>IN_1</name></connection>
<connection>
<GID>4122</GID>
<name>IN_1</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>245,23.5,246,23.5</points>
<connection>
<GID>4224</GID>
<name>OUT_0</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>2999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,11.5,281.5,151.5</points>
<connection>
<GID>4102</GID>
<name>N_in0</name></connection>
<connection>
<GID>4094</GID>
<name>N_in1</name></connection>
<intersection>31.5 1</intersection>
<intersection>48.5 3</intersection>
<intersection>64.5 4</intersection>
<intersection>80 5</intersection>
<intersection>96.5 6</intersection>
<intersection>113.5 7</intersection>
<intersection>129.5 8</intersection>
<intersection>145 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,31.5,282.5,31.5</points>
<connection>
<GID>4106</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,145,285,145</points>
<connection>
<GID>4311</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281.5,48.5,283,48.5</points>
<connection>
<GID>4130</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>281.5,64.5,283.5,64.5</points>
<connection>
<GID>4154</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>281.5,80,284,80</points>
<connection>
<GID>4178</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>281.5,96.5,283.5,96.5</points>
<connection>
<GID>4236</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>281.5,113.5,284,113.5</points>
<connection>
<GID>4263</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>281.5,129.5,284.5,129.5</points>
<connection>
<GID>4287</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,11.5,313.5,151.5</points>
<connection>
<GID>4103</GID>
<name>N_in0</name></connection>
<connection>
<GID>4109</GID>
<name>IN_0</name></connection>
<connection>
<GID>4095</GID>
<name>N_in1</name></connection>
<intersection>48.5 9</intersection>
<intersection>64.5 10</intersection>
<intersection>80 7</intersection>
<intersection>96.5 11</intersection>
<intersection>113.5 5</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,145,316,145</points>
<connection>
<GID>4314</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313.5,129.5,315.5,129.5</points>
<connection>
<GID>4290</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>313.5,113.5,315,113.5</points>
<connection>
<GID>4266</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>313.5,80,315,80</points>
<connection>
<GID>4181</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>313.5,48.5,314,48.5</points>
<connection>
<GID>4133</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>313.5,64.5,314.5,64.5</points>
<connection>
<GID>4157</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>313.5,96.5,314.5,96.5</points>
<connection>
<GID>4242</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3001</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,12.5,344.5,151.5</points>
<connection>
<GID>4197</GID>
<name>N_in0</name></connection>
<connection>
<GID>4112</GID>
<name>IN_0</name></connection>
<connection>
<GID>4096</GID>
<name>N_in1</name></connection>
<intersection>48.5 38</intersection>
<intersection>64.5 21</intersection>
<intersection>80 7</intersection>
<intersection>96.5 20</intersection>
<intersection>113.5 5</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,145,347,145</points>
<connection>
<GID>4317</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>344.5,129.5,346.5,129.5</points>
<connection>
<GID>4293</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>344.5,113.5,346,113.5</points>
<connection>
<GID>4269</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>344.5,80,346,80</points>
<connection>
<GID>4184</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>344.5,96.5,345.5,96.5</points>
<connection>
<GID>4245</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>344.5,64.5,345.5,64.5</points>
<connection>
<GID>4160</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>344.5,48.5,345,48.5</points>
<connection>
<GID>4136</GID>
<name>IN_0</name></connection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,48.5,375.5,151</points>
<connection>
<GID>4248</GID>
<name>IN_0</name></connection>
<connection>
<GID>4163</GID>
<name>IN_0</name></connection>
<connection>
<GID>4198</GID>
<name>N_in0</name></connection>
<intersection>48.5 9</intersection>
<intersection>80 7</intersection>
<intersection>113.5 5</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,145,377,145</points>
<connection>
<GID>4320</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,129.5,376.5,129.5</points>
<connection>
<GID>4296</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>375.5,113.5,376,113.5</points>
<connection>
<GID>4272</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>375.5,80,376,80</points>
<connection>
<GID>4187</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>374.5,48.5,375.5,48.5</points>
<connection>
<GID>4139</GID>
<name>IN_0</name></connection>
<intersection>374.5 10</intersection>
<intersection>375.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>374.5,13.5,374.5,48.5</points>
<connection>
<GID>4115</GID>
<name>IN_0</name></connection>
<connection>
<GID>4097</GID>
<name>N_in1</name></connection>
<intersection>48.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>3003</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405.5,14,405.5,151.5</points>
<connection>
<GID>4199</GID>
<name>N_in0</name></connection>
<connection>
<GID>4118</GID>
<name>IN_0</name></connection>
<connection>
<GID>4098</GID>
<name>N_in1</name></connection>
<intersection>48.5 13</intersection>
<intersection>64.5 11</intersection>
<intersection>80 9</intersection>
<intersection>96.5 7</intersection>
<intersection>113.5 5</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>405.5,145,408,145</points>
<connection>
<GID>4323</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>405.5,129.5,407.5,129.5</points>
<connection>
<GID>4299</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>405.5,113.5,407,113.5</points>
<connection>
<GID>4275</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>405.5,96.5,406.5,96.5</points>
<connection>
<GID>4251</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>405.5,80,407,80</points>
<connection>
<GID>4190</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>405.5,64.5,406.5,64.5</points>
<connection>
<GID>4166</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>405.5,48.5,406,48.5</points>
<connection>
<GID>4142</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436.5,15,436.5,151.5</points>
<connection>
<GID>4200</GID>
<name>N_in0</name></connection>
<connection>
<GID>4121</GID>
<name>IN_0</name></connection>
<connection>
<GID>4100</GID>
<name>N_in1</name></connection>
<intersection>48.5 13</intersection>
<intersection>64.5 11</intersection>
<intersection>80 9</intersection>
<intersection>96.5 7</intersection>
<intersection>113.5 5</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,145,439,145</points>
<connection>
<GID>4326</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436.5,129.5,438.5,129.5</points>
<connection>
<GID>4302</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>436.5,113.5,438,113.5</points>
<connection>
<GID>4278</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>436.5,96.5,437.5,96.5</points>
<connection>
<GID>4254</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>436.5,80,438,80</points>
<connection>
<GID>4193</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>436.5,64.5,437.5,64.5</points>
<connection>
<GID>4169</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>436.5,48.5,437,48.5</points>
<connection>
<GID>4145</GID>
<name>IN_0</name></connection>
<intersection>436.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467.5,13,467.5,151</points>
<connection>
<GID>4201</GID>
<name>N_in0</name></connection>
<connection>
<GID>4124</GID>
<name>IN_0</name></connection>
<connection>
<GID>4099</GID>
<name>N_in1</name></connection>
<intersection>48.5 13</intersection>
<intersection>64.5 10</intersection>
<intersection>80 8</intersection>
<intersection>96.5 6</intersection>
<intersection>113.5 4</intersection>
<intersection>129.5 2</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467.5,145,470,145</points>
<connection>
<GID>4329</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>467.5,129.5,469.5,129.5</points>
<connection>
<GID>4305</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>467.5,113.5,469,113.5</points>
<connection>
<GID>4281</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>467.5,96.5,468.5,96.5</points>
<connection>
<GID>4257</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>467.5,80,469,80</points>
<connection>
<GID>4196</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>467.5,64.5,468.5,64.5</points>
<connection>
<GID>4172</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>467.5,48.5,468,48.5</points>
<connection>
<GID>4148</GID>
<name>IN_0</name></connection>
<intersection>467.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,3.5,279.5,158.5</points>
<connection>
<GID>4203</GID>
<name>N_in1</name></connection>
<connection>
<GID>4202</GID>
<name>N_in0</name></connection>
<intersection>24.5 13</intersection>
<intersection>41.5 12</intersection>
<intersection>57.5 11</intersection>
<intersection>73 10</intersection>
<intersection>89.5 9</intersection>
<intersection>106.5 8</intersection>
<intersection>122.5 7</intersection>
<intersection>138 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>276,138,279.5,138</points>
<connection>
<GID>4307</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>275.5,122.5,279.5,122.5</points>
<connection>
<GID>4283</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>275,106.5,279.5,106.5</points>
<connection>
<GID>4259</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>274.5,89.5,279.5,89.5</points>
<connection>
<GID>4227</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>275,73,279.5,73</points>
<connection>
<GID>4174</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>274.5,57.5,279.5,57.5</points>
<connection>
<GID>4150</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>274,41.5,279.5,41.5</points>
<connection>
<GID>4126</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>273.5,24.5,279.5,24.5</points>
<connection>
<GID>4091</GID>
<name>OUT_0</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3007</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,24.5,310.5,158.5</points>
<connection>
<GID>4216</GID>
<name>N_in0</name></connection>
<intersection>24.5 13</intersection>
<intersection>41.5 12</intersection>
<intersection>57.5 11</intersection>
<intersection>73 10</intersection>
<intersection>89.5 9</intersection>
<intersection>106.5 8</intersection>
<intersection>122.5 7</intersection>
<intersection>138 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>307.5,138,310.5,138</points>
<connection>
<GID>4310</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>307,122.5,310.5,122.5</points>
<connection>
<GID>4286</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>306.5,106.5,310.5,106.5</points>
<connection>
<GID>4262</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>306,89.5,310.5,89.5</points>
<connection>
<GID>4234</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>306.5,73,310.5,73</points>
<connection>
<GID>4177</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>306,57.5,310.5,57.5</points>
<connection>
<GID>4153</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>305.5,41.5,310.5,41.5</points>
<connection>
<GID>4129</GID>
<name>OUT_0</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>305,24.5,310.5,24.5</points>
<connection>
<GID>4105</GID>
<name>OUT_0</name></connection>
<intersection>309 22</intersection>
<intersection>310.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>309,5,309,24.5</points>
<connection>
<GID>5775</GID>
<name>N_in1</name></connection>
<intersection>24.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>3008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342.5,4.5,342.5,158.5</points>
<connection>
<GID>4215</GID>
<name>N_in0</name></connection>
<connection>
<GID>4204</GID>
<name>N_in1</name></connection>
<intersection>24.5 13</intersection>
<intersection>41.5 12</intersection>
<intersection>57.5 11</intersection>
<intersection>73 10</intersection>
<intersection>89.5 9</intersection>
<intersection>106.5 8</intersection>
<intersection>122.5 7</intersection>
<intersection>138 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>338,138,342.5,138</points>
<connection>
<GID>4313</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>337.5,122.5,342.5,122.5</points>
<connection>
<GID>4289</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>337,106.5,342.5,106.5</points>
<connection>
<GID>4265</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>336.5,89.5,342.5,89.5</points>
<connection>
<GID>4240</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>337,73,342.5,73</points>
<connection>
<GID>4180</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>336.5,57.5,342.5,57.5</points>
<connection>
<GID>4156</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>336,41.5,342.5,41.5</points>
<connection>
<GID>4132</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>335.5,24.5,342.5,24.5</points>
<connection>
<GID>4108</GID>
<name>OUT_0</name></connection>
<intersection>342.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3009</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,5,373,158.5</points>
<connection>
<GID>4214</GID>
<name>N_in0</name></connection>
<connection>
<GID>4205</GID>
<name>N_in1</name></connection>
<intersection>24.5 18</intersection>
<intersection>41.5 17</intersection>
<intersection>57.5 16</intersection>
<intersection>73 15</intersection>
<intersection>89.5 14</intersection>
<intersection>106.5 13</intersection>
<intersection>122.5 12</intersection>
<intersection>138 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>369.5,138,373,138</points>
<connection>
<GID>4316</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>369,122.5,373,122.5</points>
<connection>
<GID>4292</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>368.5,106.5,373,106.5</points>
<connection>
<GID>4268</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>368,89.5,373,89.5</points>
<connection>
<GID>4244</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>368.5,73,373,73</points>
<connection>
<GID>4183</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>368,57.5,373,57.5</points>
<connection>
<GID>4159</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>367.5,41.5,373,41.5</points>
<connection>
<GID>4135</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>367,24.5,373,24.5</points>
<connection>
<GID>4111</GID>
<name>OUT_0</name></connection>
<intersection>373 0</intersection></hsegment></shape></wire>
<wire>
<ID>3010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403.5,5,403.5,158.5</points>
<connection>
<GID>4213</GID>
<name>N_in0</name></connection>
<connection>
<GID>4206</GID>
<name>N_in1</name></connection>
<intersection>24.5 9</intersection>
<intersection>41.5 10</intersection>
<intersection>57.5 11</intersection>
<intersection>73 12</intersection>
<intersection>89.5 13</intersection>
<intersection>106.5 14</intersection>
<intersection>122.5 15</intersection>
<intersection>138 16</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>396.5,24.5,403.5,24.5</points>
<connection>
<GID>4114</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>397,41.5,403.5,41.5</points>
<connection>
<GID>4138</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>397.5,57.5,403.5,57.5</points>
<connection>
<GID>4162</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>398,73,403.5,73</points>
<connection>
<GID>4186</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>397.5,89.5,403.5,89.5</points>
<connection>
<GID>4247</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>398,106.5,403.5,106.5</points>
<connection>
<GID>4271</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>398.5,122.5,403.5,122.5</points>
<connection>
<GID>4295</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>399,138,403.5,138</points>
<connection>
<GID>4319</GID>
<name>OUT_0</name></connection>
<intersection>403.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,5,434.5,158.5</points>
<connection>
<GID>4212</GID>
<name>N_in0</name></connection>
<connection>
<GID>4207</GID>
<name>N_in1</name></connection>
<intersection>24.5 6</intersection>
<intersection>41.5 7</intersection>
<intersection>57.5 8</intersection>
<intersection>73 9</intersection>
<intersection>89.5 10</intersection>
<intersection>106.5 11</intersection>
<intersection>122.5 12</intersection>
<intersection>138 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>428,24.5,434.5,24.5</points>
<connection>
<GID>4117</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>428.5,41.5,434.5,41.5</points>
<connection>
<GID>4141</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>429,57.5,434.5,57.5</points>
<connection>
<GID>4165</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>429.5,73,434.5,73</points>
<connection>
<GID>4189</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>429,89.5,434.5,89.5</points>
<connection>
<GID>4250</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>429.5,106.5,434.5,106.5</points>
<connection>
<GID>4274</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>430,122.5,434.5,122.5</points>
<connection>
<GID>4298</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>430.5,138,434.5,138</points>
<connection>
<GID>4322</GID>
<name>OUT_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465.5,4.5,465.5,159.5</points>
<connection>
<GID>4211</GID>
<name>N_in0</name></connection>
<connection>
<GID>4208</GID>
<name>N_in1</name></connection>
<intersection>24.5 6</intersection>
<intersection>41.5 7</intersection>
<intersection>57.5 8</intersection>
<intersection>73 9</intersection>
<intersection>89.5 10</intersection>
<intersection>106.5 11</intersection>
<intersection>122.5 12</intersection>
<intersection>138 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>458.5,24.5,465.5,24.5</points>
<connection>
<GID>4120</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>459,41.5,465.5,41.5</points>
<connection>
<GID>4144</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>459.5,57.5,465.5,57.5</points>
<connection>
<GID>4168</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>460,73,465.5,73</points>
<connection>
<GID>4192</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>459.5,89.5,465.5,89.5</points>
<connection>
<GID>4253</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>460,106.5,465.5,106.5</points>
<connection>
<GID>4277</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>460.5,122.5,465.5,122.5</points>
<connection>
<GID>4301</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>461,138,465.5,138</points>
<connection>
<GID>4325</GID>
<name>OUT_0</name></connection>
<intersection>465.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496,5,496,160</points>
<connection>
<GID>4210</GID>
<name>N_in0</name></connection>
<connection>
<GID>4209</GID>
<name>N_in1</name></connection>
<intersection>24.5 3</intersection>
<intersection>41.5 4</intersection>
<intersection>57.5 5</intersection>
<intersection>73 6</intersection>
<intersection>89.5 7</intersection>
<intersection>106.5 8</intersection>
<intersection>122.5 9</intersection>
<intersection>138 10</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>490,24.5,496,24.5</points>
<connection>
<GID>4123</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>490.5,41.5,496,41.5</points>
<connection>
<GID>4147</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>491,57.5,496,57.5</points>
<connection>
<GID>4171</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>491.5,73,496,73</points>
<connection>
<GID>4195</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>491,89.5,496,89.5</points>
<connection>
<GID>4256</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>491.5,106.5,496,106.5</points>
<connection>
<GID>4280</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>492,122.5,496,122.5</points>
<connection>
<GID>4304</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>492.5,138,496,138</points>
<connection>
<GID>4328</GID>
<name>OUT_0</name></connection>
<intersection>496 0</intersection></hsegment></shape></wire>
<wire>
<ID>3014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,90.5,204.5,139.5</points>
<intersection>90.5 2</intersection>
<intersection>139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,139.5,243.5,139.5</points>
<connection>
<GID>4229</GID>
<name>ENABLE_0</name></connection>
<intersection>204.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,90.5,204.5,90.5</points>
<connection>
<GID>4217</GID>
<name>OUT_7</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,139.5,229.5,143</points>
<intersection>139.5 1</intersection>
<intersection>143 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,143,234,143</points>
<connection>
<GID>4230</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,89.5,206.5,124</points>
<intersection>89.5 2</intersection>
<intersection>124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,124,243.5,124</points>
<intersection>206.5 0</intersection>
<intersection>229.5 4</intersection>
<intersection>243.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,89.5,206.5,89.5</points>
<connection>
<GID>4217</GID>
<name>OUT_6</name></connection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243.5,123.5,243.5,124</points>
<connection>
<GID>4231</GID>
<name>ENABLE_0</name></connection>
<intersection>124 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>229.5,124,229.5,127.5</points>
<intersection>124 1</intersection>
<intersection>127.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,127.5,233.5,127.5</points>
<connection>
<GID>4233</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,88.5,208.5,111.5</points>
<intersection>88.5 2</intersection>
<intersection>111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,111.5,233.5,111.5</points>
<connection>
<GID>4237</GID>
<name>IN_0</name></connection>
<intersection>208.5 0</intersection>
<intersection>229.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,88.5,208.5,88.5</points>
<connection>
<GID>4217</GID>
<name>OUT_5</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229.5,107.5,229.5,111.5</points>
<intersection>107.5 4</intersection>
<intersection>111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229.5,107.5,243.5,107.5</points>
<connection>
<GID>4235</GID>
<name>ENABLE_0</name></connection>
<intersection>229.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,87.5,210.5,94.5</points>
<intersection>87.5 2</intersection>
<intersection>94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,94.5,233.5,94.5</points>
<connection>
<GID>4241</GID>
<name>IN_0</name></connection>
<intersection>210.5 0</intersection>
<intersection>229.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,87.5,210.5,87.5</points>
<connection>
<GID>4217</GID>
<name>OUT_4</name></connection>
<intersection>210.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>229.5,90.5,229.5,94.5</points>
<intersection>90.5 4</intersection>
<intersection>94.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>229.5,90.5,243.5,90.5</points>
<connection>
<GID>4239</GID>
<name>ENABLE_0</name></connection>
<intersection>229.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,74.5,210.5,86.5</points>
<intersection>74.5 1</intersection>
<intersection>86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,74.5,242.5,74.5</points>
<connection>
<GID>4218</GID>
<name>ENABLE_0</name></connection>
<intersection>210.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,86.5,210.5,86.5</points>
<connection>
<GID>4217</GID>
<name>OUT_3</name></connection>
<intersection>210.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,74.5,229.5,78</points>
<intersection>74.5 1</intersection>
<intersection>78 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,78,233.5,78</points>
<connection>
<GID>4219</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,58.5,208.5,85.5</points>
<intersection>58.5 1</intersection>
<intersection>85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,58.5,242.5,58.5</points>
<connection>
<GID>4220</GID>
<name>ENABLE_0</name></connection>
<intersection>208.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,85.5,208.5,85.5</points>
<connection>
<GID>4217</GID>
<name>OUT_2</name></connection>
<intersection>208.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,58.5,229.5,62.5</points>
<intersection>58.5 1</intersection>
<intersection>62.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,62.5,233.5,62.5</points>
<connection>
<GID>4221</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,43,206.5,84.5</points>
<intersection>43 1</intersection>
<intersection>84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206.5,43,242.5,43</points>
<intersection>206.5 0</intersection>
<intersection>229.5 4</intersection>
<intersection>242.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,84.5,206.5,84.5</points>
<connection>
<GID>4217</GID>
<name>OUT_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242.5,42.5,242.5,43</points>
<connection>
<GID>4222</GID>
<name>ENABLE_0</name></connection>
<intersection>43 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>229.5,43,229.5,46.5</points>
<intersection>43 1</intersection>
<intersection>46.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,46.5,233.5,46.5</points>
<connection>
<GID>4223</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,25.5,204.5,83.5</points>
<intersection>25.5 1</intersection>
<intersection>83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,25.5,242.5,25.5</points>
<connection>
<GID>4224</GID>
<name>ENABLE_0</name></connection>
<intersection>204.5 0</intersection>
<intersection>229.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,83.5,204.5,83.5</points>
<connection>
<GID>4217</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>229.5,25.5,229.5,29.5</points>
<intersection>25.5 1</intersection>
<intersection>29.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>229.5,29.5,233.5,29.5</points>
<connection>
<GID>4225</GID>
<name>IN_0</name></connection>
<intersection>229.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3022</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>270.5,87,272.5,87</points>
<connection>
<GID>4226</GID>
<name>OUT</name></connection>
<connection>
<GID>4227</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,83.5,274.5,84</points>
<connection>
<GID>4227</GID>
<name>IN_0</name></connection>
<intersection>83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260.5,83.5,274.5,83.5</points>
<intersection>260.5 2</intersection>
<intersection>274.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>260.5,83.5,260.5,96.5</points>
<intersection>83.5 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260.5,88,264.5,88</points>
<connection>
<GID>4226</GID>
<name>IN_0</name></connection>
<intersection>260.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>258.5,96.5,260.5,96.5</points>
<connection>
<GID>4228</GID>
<name>OUT_0</name></connection>
<intersection>260.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3024</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302,87,304,87</points>
<connection>
<GID>4232</GID>
<name>OUT</name></connection>
<connection>
<GID>4234</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3025</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292,84,306,84</points>
<connection>
<GID>4234</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292,84,292,96.5</points>
<intersection>84 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292,88,296,88</points>
<connection>
<GID>4232</GID>
<name>IN_0</name></connection>
<intersection>292 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289.5,96.5,292,96.5</points>
<connection>
<GID>4236</GID>
<name>OUT_0</name></connection>
<intersection>292 2</intersection></hsegment></shape></wire>
<wire>
<ID>3026</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>332.5,87,334.5,87</points>
<connection>
<GID>4238</GID>
<name>OUT</name></connection>
<connection>
<GID>4240</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3027</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,83.5,336.5,84</points>
<connection>
<GID>4240</GID>
<name>IN_0</name></connection>
<intersection>83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,83.5,336.5,83.5</points>
<intersection>322.5 2</intersection>
<intersection>336.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322.5,83.5,322.5,96.5</points>
<intersection>83.5 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>322.5,88,326.5,88</points>
<connection>
<GID>4238</GID>
<name>IN_0</name></connection>
<intersection>322.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320.5,96.5,322.5,96.5</points>
<connection>
<GID>4242</GID>
<name>OUT_0</name></connection>
<intersection>322.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3028</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364,87,366,87</points>
<connection>
<GID>4243</GID>
<name>OUT</name></connection>
<connection>
<GID>4244</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3029</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354,84,368,84</points>
<connection>
<GID>4244</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354,84,354,96.5</points>
<intersection>84 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354,88,358,88</points>
<connection>
<GID>4243</GID>
<name>IN_0</name></connection>
<intersection>354 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>351.5,96.5,354,96.5</points>
<connection>
<GID>4245</GID>
<name>OUT_0</name></connection>
<intersection>354 2</intersection></hsegment></shape></wire>
<wire>
<ID>3030</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>393.5,87,395.5,87</points>
<connection>
<GID>4246</GID>
<name>OUT</name></connection>
<connection>
<GID>4247</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,83.5,397.5,84</points>
<connection>
<GID>4247</GID>
<name>IN_0</name></connection>
<intersection>83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,83.5,397.5,83.5</points>
<intersection>383.5 2</intersection>
<intersection>397.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383.5,83.5,383.5,96.5</points>
<intersection>83.5 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>383.5,88,387.5,88</points>
<connection>
<GID>4246</GID>
<name>IN_0</name></connection>
<intersection>383.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>381.5,96.5,383.5,96.5</points>
<connection>
<GID>4248</GID>
<name>OUT_0</name></connection>
<intersection>383.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3032</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425,87,427,87</points>
<connection>
<GID>4249</GID>
<name>OUT</name></connection>
<connection>
<GID>4250</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415,84,429,84</points>
<connection>
<GID>4250</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415,84,415,96.5</points>
<intersection>84 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415,88,419,88</points>
<connection>
<GID>4249</GID>
<name>IN_0</name></connection>
<intersection>415 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>412.5,96.5,415,96.5</points>
<connection>
<GID>4251</GID>
<name>OUT_0</name></connection>
<intersection>415 2</intersection></hsegment></shape></wire>
<wire>
<ID>3034</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>455.5,87,457.5,87</points>
<connection>
<GID>4252</GID>
<name>OUT</name></connection>
<connection>
<GID>4253</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,83.5,459.5,84</points>
<connection>
<GID>4253</GID>
<name>IN_0</name></connection>
<intersection>83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,83.5,459.5,83.5</points>
<intersection>445.5 2</intersection>
<intersection>459.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>445.5,83.5,445.5,96.5</points>
<intersection>83.5 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>445.5,88,449.5,88</points>
<connection>
<GID>4252</GID>
<name>IN_0</name></connection>
<intersection>445.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443.5,96.5,445.5,96.5</points>
<connection>
<GID>4254</GID>
<name>OUT_0</name></connection>
<intersection>445.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3036</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487,87,489,87</points>
<connection>
<GID>4255</GID>
<name>OUT</name></connection>
<connection>
<GID>4256</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,84,491,84</points>
<connection>
<GID>4256</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477,84,477,96.5</points>
<intersection>84 1</intersection>
<intersection>88 4</intersection>
<intersection>96.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477,88,481,88</points>
<connection>
<GID>4255</GID>
<name>IN_0</name></connection>
<intersection>477 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>474.5,96.5,477,96.5</points>
<connection>
<GID>4257</GID>
<name>OUT_0</name></connection>
<intersection>477 2</intersection></hsegment></shape></wire>
<wire>
<ID>3038</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271,104,273,104</points>
<connection>
<GID>4258</GID>
<name>OUT</name></connection>
<connection>
<GID>4259</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,100.5,275,101</points>
<connection>
<GID>4259</GID>
<name>IN_0</name></connection>
<intersection>100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,100.5,275,100.5</points>
<intersection>261 2</intersection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261,100.5,261,113.5</points>
<intersection>100.5 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,105,265,105</points>
<connection>
<GID>4258</GID>
<name>IN_0</name></connection>
<intersection>261 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259,113.5,261,113.5</points>
<connection>
<GID>4260</GID>
<name>OUT_0</name></connection>
<intersection>261 2</intersection></hsegment></shape></wire>
<wire>
<ID>3040</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>302.5,104,304.5,104</points>
<connection>
<GID>4261</GID>
<name>OUT</name></connection>
<connection>
<GID>4262</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,101,306.5,101</points>
<connection>
<GID>4262</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>292.5,101,292.5,113.5</points>
<intersection>101 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>292.5,105,296.5,105</points>
<connection>
<GID>4261</GID>
<name>IN_0</name></connection>
<intersection>292.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290,113.5,292.5,113.5</points>
<connection>
<GID>4263</GID>
<name>OUT_0</name></connection>
<intersection>292.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3042</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333,104,335,104</points>
<connection>
<GID>4264</GID>
<name>OUT</name></connection>
<connection>
<GID>4265</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,100.5,337,101</points>
<connection>
<GID>4265</GID>
<name>IN_0</name></connection>
<intersection>100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,100.5,337,100.5</points>
<intersection>323 2</intersection>
<intersection>337 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323,100.5,323,113.5</points>
<intersection>100.5 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323,105,327,105</points>
<connection>
<GID>4264</GID>
<name>IN_0</name></connection>
<intersection>323 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321,113.5,323,113.5</points>
<connection>
<GID>4266</GID>
<name>OUT_0</name></connection>
<intersection>323 2</intersection></hsegment></shape></wire>
<wire>
<ID>3044</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>364.5,104,366.5,104</points>
<connection>
<GID>4267</GID>
<name>OUT</name></connection>
<connection>
<GID>4268</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,101,368.5,101</points>
<connection>
<GID>4268</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>354.5,101,354.5,113.5</points>
<intersection>101 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354.5,105,358.5,105</points>
<connection>
<GID>4267</GID>
<name>IN_0</name></connection>
<intersection>354.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352,113.5,354.5,113.5</points>
<connection>
<GID>4269</GID>
<name>OUT_0</name></connection>
<intersection>354.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3046</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394,104,396,104</points>
<connection>
<GID>4270</GID>
<name>OUT</name></connection>
<connection>
<GID>4271</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,100.5,398,101</points>
<connection>
<GID>4271</GID>
<name>IN_0</name></connection>
<intersection>100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,100.5,398,100.5</points>
<intersection>384 2</intersection>
<intersection>398 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384,100.5,384,113.5</points>
<intersection>100.5 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384,105,388,105</points>
<connection>
<GID>4270</GID>
<name>IN_0</name></connection>
<intersection>384 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382,113.5,384,113.5</points>
<connection>
<GID>4272</GID>
<name>OUT_0</name></connection>
<intersection>384 2</intersection></hsegment></shape></wire>
<wire>
<ID>3048</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425.5,104,427.5,104</points>
<connection>
<GID>4273</GID>
<name>OUT</name></connection>
<connection>
<GID>4274</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>415.5,101,429.5,101</points>
<connection>
<GID>4274</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>415.5,101,415.5,113.5</points>
<intersection>101 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415.5,105,419.5,105</points>
<connection>
<GID>4273</GID>
<name>IN_0</name></connection>
<intersection>415.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413,113.5,415.5,113.5</points>
<connection>
<GID>4275</GID>
<name>OUT_0</name></connection>
<intersection>415.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3050</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456,104,458,104</points>
<connection>
<GID>4276</GID>
<name>OUT</name></connection>
<connection>
<GID>4277</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460,100.5,460,101</points>
<connection>
<GID>4277</GID>
<name>IN_0</name></connection>
<intersection>100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446,100.5,460,100.5</points>
<intersection>446 2</intersection>
<intersection>460 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446,100.5,446,113.5</points>
<intersection>100.5 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446,105,450,105</points>
<connection>
<GID>4276</GID>
<name>IN_0</name></connection>
<intersection>446 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444,113.5,446,113.5</points>
<connection>
<GID>4278</GID>
<name>OUT_0</name></connection>
<intersection>446 2</intersection></hsegment></shape></wire>
<wire>
<ID>3052</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>487.5,104,489.5,104</points>
<connection>
<GID>4279</GID>
<name>OUT</name></connection>
<connection>
<GID>4280</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,101,491.5,101</points>
<connection>
<GID>4280</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477.5,101,477.5,113.5</points>
<intersection>101 1</intersection>
<intersection>105 4</intersection>
<intersection>113.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477.5,105,481.5,105</points>
<connection>
<GID>4279</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475,113.5,477.5,113.5</points>
<connection>
<GID>4281</GID>
<name>OUT_0</name></connection>
<intersection>477.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3054</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>271.5,120,273.5,120</points>
<connection>
<GID>4282</GID>
<name>OUT</name></connection>
<connection>
<GID>4283</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,116.5,275.5,117</points>
<connection>
<GID>4283</GID>
<name>IN_0</name></connection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,116.5,275.5,116.5</points>
<intersection>261.5 2</intersection>
<intersection>275.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>261.5,116.5,261.5,129.5</points>
<intersection>116.5 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261.5,121,265.5,121</points>
<connection>
<GID>4282</GID>
<name>IN_0</name></connection>
<intersection>261.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>259.5,129.5,261.5,129.5</points>
<connection>
<GID>4284</GID>
<name>OUT_0</name></connection>
<intersection>261.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3056</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>303,120,305,120</points>
<connection>
<GID>4285</GID>
<name>OUT</name></connection>
<connection>
<GID>4286</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293,117,307,117</points>
<connection>
<GID>4286</GID>
<name>IN_0</name></connection>
<intersection>293 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>293,117,293,129.5</points>
<intersection>117 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>293,121,297,121</points>
<connection>
<GID>4285</GID>
<name>IN_0</name></connection>
<intersection>293 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>290.5,129.5,293,129.5</points>
<connection>
<GID>4287</GID>
<name>OUT_0</name></connection>
<intersection>293 2</intersection></hsegment></shape></wire>
<wire>
<ID>3058</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>333.5,120,335.5,120</points>
<connection>
<GID>4288</GID>
<name>OUT</name></connection>
<connection>
<GID>4289</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,116.5,337.5,117</points>
<connection>
<GID>4289</GID>
<name>IN_0</name></connection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,116.5,337.5,116.5</points>
<intersection>323.5 2</intersection>
<intersection>337.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323.5,116.5,323.5,129.5</points>
<intersection>116.5 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>323.5,121,327.5,121</points>
<connection>
<GID>4288</GID>
<name>IN_0</name></connection>
<intersection>323.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>321.5,129.5,323.5,129.5</points>
<connection>
<GID>4290</GID>
<name>OUT_0</name></connection>
<intersection>323.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3060</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>365,120,367,120</points>
<connection>
<GID>4291</GID>
<name>OUT</name></connection>
<connection>
<GID>4292</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,117,369,117</points>
<connection>
<GID>4292</GID>
<name>IN_0</name></connection>
<intersection>355 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>355,117,355,129.5</points>
<intersection>117 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>355,121,359,121</points>
<connection>
<GID>4291</GID>
<name>IN_0</name></connection>
<intersection>355 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352.5,129.5,355,129.5</points>
<connection>
<GID>4293</GID>
<name>OUT_0</name></connection>
<intersection>355 2</intersection></hsegment></shape></wire>
<wire>
<ID>3062</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>394.5,120,396.5,120</points>
<connection>
<GID>4294</GID>
<name>OUT</name></connection>
<connection>
<GID>4295</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3063</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398.5,116.5,398.5,117</points>
<connection>
<GID>4295</GID>
<name>IN_0</name></connection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,116.5,398.5,116.5</points>
<intersection>384.5 2</intersection>
<intersection>398.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>384.5,116.5,384.5,129.5</points>
<intersection>116.5 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>384.5,121,388.5,121</points>
<connection>
<GID>4294</GID>
<name>IN_0</name></connection>
<intersection>384.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>382.5,129.5,384.5,129.5</points>
<connection>
<GID>4296</GID>
<name>OUT_0</name></connection>
<intersection>384.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3064</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>426,120,428,120</points>
<connection>
<GID>4297</GID>
<name>OUT</name></connection>
<connection>
<GID>4298</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>416,117,430,117</points>
<connection>
<GID>4298</GID>
<name>IN_0</name></connection>
<intersection>416 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>416,117,416,129.5</points>
<intersection>117 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>416,121,420,121</points>
<connection>
<GID>4297</GID>
<name>IN_0</name></connection>
<intersection>416 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>413.5,129.5,416,129.5</points>
<connection>
<GID>4299</GID>
<name>OUT_0</name></connection>
<intersection>416 2</intersection></hsegment></shape></wire>
<wire>
<ID>3066</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>456.5,120,458.5,120</points>
<connection>
<GID>4300</GID>
<name>OUT</name></connection>
<connection>
<GID>4301</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3067</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>460.5,116.5,460.5,117</points>
<connection>
<GID>4301</GID>
<name>IN_0</name></connection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446.5,116.5,460.5,116.5</points>
<intersection>446.5 2</intersection>
<intersection>460.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>446.5,116.5,446.5,129.5</points>
<intersection>116.5 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>446.5,121,450.5,121</points>
<connection>
<GID>4300</GID>
<name>IN_0</name></connection>
<intersection>446.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444.5,129.5,446.5,129.5</points>
<connection>
<GID>4302</GID>
<name>OUT_0</name></connection>
<intersection>446.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3068</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>488,120,490,120</points>
<connection>
<GID>4303</GID>
<name>OUT</name></connection>
<connection>
<GID>4304</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>478,117,492,117</points>
<connection>
<GID>4304</GID>
<name>IN_0</name></connection>
<intersection>478 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>478,117,478,129.5</points>
<intersection>117 1</intersection>
<intersection>121 4</intersection>
<intersection>129.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>478,121,482,121</points>
<connection>
<GID>4303</GID>
<name>IN_0</name></connection>
<intersection>478 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>475.5,129.5,478,129.5</points>
<connection>
<GID>4305</GID>
<name>OUT_0</name></connection>
<intersection>478 2</intersection></hsegment></shape></wire>
<wire>
<ID>3070</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>272,135.5,274,135.5</points>
<connection>
<GID>4306</GID>
<name>OUT</name></connection>
<connection>
<GID>4307</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,132,276,132.5</points>
<connection>
<GID>4307</GID>
<name>IN_0</name></connection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,132,276,132</points>
<intersection>262 2</intersection>
<intersection>276 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>262,132,262,145</points>
<intersection>132 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>262,136.5,266,136.5</points>
<connection>
<GID>4306</GID>
<name>IN_0</name></connection>
<intersection>262 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>260,145,262,145</points>
<connection>
<GID>4308</GID>
<name>OUT_0</name></connection>
<intersection>262 2</intersection></hsegment></shape></wire>
<wire>
<ID>3072</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>303.5,135.5,305.5,135.5</points>
<connection>
<GID>4309</GID>
<name>OUT</name></connection>
<connection>
<GID>4310</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>293.5,132.5,307.5,132.5</points>
<connection>
<GID>4310</GID>
<name>IN_0</name></connection>
<intersection>293.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>293.5,132.5,293.5,145</points>
<intersection>132.5 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>293.5,136.5,297.5,136.5</points>
<connection>
<GID>4309</GID>
<name>IN_0</name></connection>
<intersection>293.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>291,145,293.5,145</points>
<connection>
<GID>4311</GID>
<name>OUT_0</name></connection>
<intersection>293.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3074</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>334,135.5,336,135.5</points>
<connection>
<GID>4312</GID>
<name>OUT</name></connection>
<connection>
<GID>4313</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338,132,338,132.5</points>
<connection>
<GID>4313</GID>
<name>IN_0</name></connection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324,132,338,132</points>
<intersection>324 2</intersection>
<intersection>338 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>324,132,324,145</points>
<intersection>132 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>324,136.5,328,136.5</points>
<connection>
<GID>4312</GID>
<name>IN_0</name></connection>
<intersection>324 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>322,145,324,145</points>
<connection>
<GID>4314</GID>
<name>OUT_0</name></connection>
<intersection>324 2</intersection></hsegment></shape></wire>
<wire>
<ID>3076</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>365.5,135.5,367.5,135.5</points>
<connection>
<GID>4315</GID>
<name>OUT</name></connection>
<connection>
<GID>4316</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355.5,132.5,369.5,132.5</points>
<connection>
<GID>4316</GID>
<name>IN_0</name></connection>
<intersection>355.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>355.5,132.5,355.5,145</points>
<intersection>132.5 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>355.5,136.5,359.5,136.5</points>
<connection>
<GID>4315</GID>
<name>IN_0</name></connection>
<intersection>355.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>353,145,355.5,145</points>
<connection>
<GID>4317</GID>
<name>OUT_0</name></connection>
<intersection>355.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3078</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>395,135.5,397,135.5</points>
<connection>
<GID>4318</GID>
<name>OUT</name></connection>
<connection>
<GID>4319</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,132,399,132.5</points>
<connection>
<GID>4319</GID>
<name>IN_0</name></connection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>385,132,399,132</points>
<intersection>385 2</intersection>
<intersection>399 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>385,132,385,145</points>
<intersection>132 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>385,136.5,389,136.5</points>
<connection>
<GID>4318</GID>
<name>IN_0</name></connection>
<intersection>385 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>383,145,385,145</points>
<connection>
<GID>4320</GID>
<name>OUT_0</name></connection>
<intersection>385 2</intersection></hsegment></shape></wire>
<wire>
<ID>3080</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>426.5,135.5,428.5,135.5</points>
<connection>
<GID>4321</GID>
<name>OUT</name></connection>
<connection>
<GID>4322</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3081</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>416.5,132.5,430.5,132.5</points>
<connection>
<GID>4322</GID>
<name>IN_0</name></connection>
<intersection>416.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>416.5,132.5,416.5,145</points>
<intersection>132.5 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>416.5,136.5,420.5,136.5</points>
<connection>
<GID>4321</GID>
<name>IN_0</name></connection>
<intersection>416.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>414,145,416.5,145</points>
<connection>
<GID>4323</GID>
<name>OUT_0</name></connection>
<intersection>416.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>3082</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>457,135.5,459,135.5</points>
<connection>
<GID>4324</GID>
<name>OUT</name></connection>
<connection>
<GID>4325</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461,132,461,132.5</points>
<connection>
<GID>4325</GID>
<name>IN_0</name></connection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>447,132,461,132</points>
<intersection>447 2</intersection>
<intersection>461 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>447,132,447,145</points>
<intersection>132 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>447,136.5,451,136.5</points>
<connection>
<GID>4324</GID>
<name>IN_0</name></connection>
<intersection>447 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>445,145,447,145</points>
<connection>
<GID>4326</GID>
<name>OUT_0</name></connection>
<intersection>447 2</intersection></hsegment></shape></wire>
<wire>
<ID>3084</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>488.5,135.5,490.5,135.5</points>
<connection>
<GID>4327</GID>
<name>OUT</name></connection>
<connection>
<GID>4328</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3085</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>478.5,132.5,492.5,132.5</points>
<connection>
<GID>4328</GID>
<name>IN_0</name></connection>
<intersection>478.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>478.5,132.5,478.5,145</points>
<intersection>132.5 1</intersection>
<intersection>136.5 4</intersection>
<intersection>145 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>478.5,136.5,482.5,136.5</points>
<connection>
<GID>4327</GID>
<name>IN_0</name></connection>
<intersection>478.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>476,145,478.5,145</points>
<connection>
<GID>4329</GID>
<name>OUT_0</name></connection>
<intersection>478.5 2</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 1>
<page 2>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 2>
<page 3>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 3>
<page 4>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 4>
<page 5>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>-0.000378015,33.5808,338.954,-133.958</PageViewport></page 9></circuit>